magic
tech sky130A
timestamp 1634045183
<< pwell >>
rect -717 5029 -209 5050
rect -717 -574 3227 5029
rect -510 -585 3227 -574
<< mvpsubdiff >>
rect -683 3447 -313 3532
rect -683 3300 -640 3447
rect -683 988 -644 3300
rect -372 1135 -313 3447
rect -376 988 -313 1135
rect -683 960 -313 988
<< mvpsubdiffcont >>
rect -640 3300 -372 3447
rect -644 1135 -372 3300
rect -644 988 -376 1135
<< poly >>
rect 72 4796 2770 4827
rect 47 3747 548 3781
rect 1061 3746 1562 3780
rect 2191 3747 2692 3781
rect 38 2700 539 2734
rect 1075 2700 1576 2734
rect 2104 2701 2605 2735
rect 77 1649 578 1683
rect 1121 1651 1622 1685
rect 2125 1650 2626 1684
rect 71 602 572 636
rect 1146 603 1647 637
rect 2226 604 2727 638
<< locali >>
rect -187 4649 -155 4674
rect 1874 4649 1906 4667
rect -189 4610 1906 4649
rect -187 4394 -155 4610
rect 1874 4387 1906 4610
rect -683 3447 -313 3532
rect -683 3300 -640 3447
rect -683 988 -644 3300
rect -372 1135 -313 3447
rect -376 988 -313 1135
rect -683 960 -313 988
rect -181 132 -154 4295
rect 839 119 866 4282
rect 1873 134 1900 4297
rect 2906 164 2933 4327
rect 845 -240 877 -1
rect 2901 -240 2934 2
rect 845 -281 2936 -240
rect 2901 -288 2934 -281
<< viali >>
rect -584 1358 -435 3204
<< metal1 >>
rect -683 3204 -313 3532
rect -683 1358 -584 3204
rect -435 1358 -313 3204
rect -683 960 -313 1358
use sky130_fd_pr__nfet_g5v0d10v5_C8TC2Y  sky130_fd_pr__nfet_g5v0d10v5_C8TC2Y_0 ~/layout test
timestamp 1634044821
transform 1 0 1373 0 1 2192
box -1558 -2607 1558 2607
<< end >>
