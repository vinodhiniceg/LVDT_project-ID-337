magic
tech sky130A
magscale 1 2
timestamp 1634365921
<< error_p >>
rect -70 -2600 -10 2600
rect 10 -2600 70 2600
<< metal3 >>
rect -4282 2572 -10 2600
rect -4282 -2572 -94 2572
rect -30 -2572 -10 2572
rect -4282 -2600 -10 -2572
rect 10 2572 4282 2600
rect 10 -2572 4198 2572
rect 4262 -2572 4282 2572
rect 10 -2600 4282 -2572
<< via3 >>
rect -94 -2572 -30 2572
rect 4198 -2572 4262 2572
<< mimcap >>
rect -4182 2460 -182 2500
rect -4182 -2460 -2770 2460
rect -1594 -2460 -182 2460
rect -4182 -2500 -182 -2460
rect 110 2460 4110 2500
rect 110 -2460 1522 2460
rect 2698 -2460 4110 2460
rect 110 -2500 4110 -2460
<< mimcapcontact >>
rect -2770 -2460 -1594 2460
rect 1522 -2460 2698 2460
<< metal4 >>
rect -110 2572 -14 2588
rect -2771 2460 -1593 2461
rect -2771 -2460 -2770 2460
rect -1594 -2460 -1593 2460
rect -2771 -2461 -1593 -2460
rect -110 -2572 -94 2572
rect -30 -2572 -14 2572
rect 4182 2572 4278 2588
rect 1521 2460 2699 2461
rect 1521 -2460 1522 2460
rect 2698 -2460 2699 2460
rect 1521 -2461 2699 -2460
rect -110 -2588 -14 -2572
rect 4182 -2572 4198 2572
rect 4262 -2572 4278 2572
rect 4182 -2588 4278 -2572
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX 10 -2600 4210 2600
string parameters w 20.00 l 25.00 val 1.017k carea 2.00 cperi 0.19 nx 2 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 30
string library sky130
<< end >>
