magic
tech sky130A
timestamp 1634044821
<< error_p >>
rect -1558 1594 -1529 2594
rect -529 1594 -500 2594
rect 500 1594 529 2594
rect 1529 1594 1558 2594
rect -1558 547 -1529 1547
rect -529 547 -500 1547
rect 500 547 529 1547
rect 1529 547 1558 1547
rect -1558 -500 -1529 500
rect -529 -500 -500 500
rect 500 -500 529 500
rect 1529 -500 1558 500
rect -1558 -1547 -1529 -547
rect -529 -1547 -500 -547
rect 500 -1547 529 -547
rect 1529 -1547 1558 -547
rect -1558 -2594 -1529 -1594
rect -529 -2594 -500 -1594
rect 500 -2594 529 -1594
rect 1529 -2594 1558 -1594
<< mvnmos >>
rect -1529 1594 -529 2594
rect -500 1594 500 2594
rect 529 1594 1529 2594
rect -1529 547 -529 1547
rect -500 547 500 1547
rect 529 547 1529 1547
rect -1529 -500 -529 500
rect -500 -500 500 500
rect 529 -500 1529 500
rect -1529 -1547 -529 -547
rect -500 -1547 500 -547
rect 529 -1547 1529 -547
rect -1529 -2594 -529 -1594
rect -500 -2594 500 -1594
rect 529 -2594 1529 -1594
<< mvndiff >>
rect -1558 2242 -1529 2594
rect -1558 1946 -1552 2242
rect -1535 1946 -1529 2242
rect -1558 1594 -1529 1946
rect -529 2242 -500 2594
rect -529 1946 -523 2242
rect -506 1946 -500 2242
rect -529 1594 -500 1946
rect 500 2242 529 2594
rect 500 1946 506 2242
rect 523 1946 529 2242
rect 500 1594 529 1946
rect 1529 2242 1558 2594
rect 1529 1946 1535 2242
rect 1552 1946 1558 2242
rect 1529 1594 1558 1946
rect -1558 1195 -1529 1547
rect -1558 899 -1552 1195
rect -1535 899 -1529 1195
rect -1558 547 -1529 899
rect -529 1195 -500 1547
rect -529 899 -523 1195
rect -506 899 -500 1195
rect -529 547 -500 899
rect 500 1195 529 1547
rect 500 899 506 1195
rect 523 899 529 1195
rect 500 547 529 899
rect 1529 1195 1558 1547
rect 1529 899 1535 1195
rect 1552 899 1558 1195
rect 1529 547 1558 899
rect -1558 148 -1529 500
rect -1558 -148 -1552 148
rect -1535 -148 -1529 148
rect -1558 -500 -1529 -148
rect -529 148 -500 500
rect -529 -148 -523 148
rect -506 -148 -500 148
rect -529 -500 -500 -148
rect 500 148 529 500
rect 500 -148 506 148
rect 523 -148 529 148
rect 500 -500 529 -148
rect 1529 148 1558 500
rect 1529 -148 1535 148
rect 1552 -148 1558 148
rect 1529 -500 1558 -148
rect -1558 -899 -1529 -547
rect -1558 -1195 -1552 -899
rect -1535 -1195 -1529 -899
rect -1558 -1547 -1529 -1195
rect -529 -899 -500 -547
rect -529 -1195 -523 -899
rect -506 -1195 -500 -899
rect -529 -1547 -500 -1195
rect 500 -899 529 -547
rect 500 -1195 506 -899
rect 523 -1195 529 -899
rect 500 -1547 529 -1195
rect 1529 -899 1558 -547
rect 1529 -1195 1535 -899
rect 1552 -1195 1558 -899
rect 1529 -1547 1558 -1195
rect -1558 -1946 -1529 -1594
rect -1558 -2242 -1552 -1946
rect -1535 -2242 -1529 -1946
rect -1558 -2594 -1529 -2242
rect -529 -1946 -500 -1594
rect -529 -2242 -523 -1946
rect -506 -2242 -500 -1946
rect -529 -2594 -500 -2242
rect 500 -1946 529 -1594
rect 500 -2242 506 -1946
rect 523 -2242 529 -1946
rect 500 -2594 529 -2242
rect 1529 -1946 1558 -1594
rect 1529 -2242 1535 -1946
rect 1552 -2242 1558 -1946
rect 1529 -2594 1558 -2242
<< mvndiffc >>
rect -1552 1946 -1535 2242
rect -523 1946 -506 2242
rect 506 1946 523 2242
rect 1535 1946 1552 2242
rect -1552 899 -1535 1195
rect -523 899 -506 1195
rect 506 899 523 1195
rect 1535 899 1552 1195
rect -1552 -148 -1535 148
rect -523 -148 -506 148
rect 506 -148 523 148
rect 1535 -148 1552 148
rect -1552 -1195 -1535 -899
rect -523 -1195 -506 -899
rect 506 -1195 523 -899
rect 1535 -1195 1552 -899
rect -1552 -2242 -1535 -1946
rect -523 -2242 -506 -1946
rect 506 -2242 523 -1946
rect 1535 -2242 1552 -1946
<< poly >>
rect -1529 2594 -529 2607
rect -500 2594 500 2607
rect 529 2594 1529 2607
rect -1529 1581 -529 1594
rect -500 1581 500 1594
rect 529 1581 1529 1594
rect -1529 1547 -529 1560
rect -500 1547 500 1560
rect 529 1547 1529 1560
rect -1529 534 -529 547
rect -500 534 500 547
rect 529 534 1529 547
rect -1529 500 -529 513
rect -500 500 500 513
rect 529 500 1529 513
rect -1529 -513 -529 -500
rect -500 -513 500 -500
rect 529 -513 1529 -500
rect -1529 -547 -529 -534
rect -500 -547 500 -534
rect 529 -547 1529 -534
rect -1529 -1560 -529 -1547
rect -500 -1560 500 -1547
rect 529 -1560 1529 -1547
rect -1529 -1594 -529 -1581
rect -500 -1594 500 -1581
rect 529 -1594 1529 -1581
rect -1529 -2607 -529 -2594
rect -500 -2607 500 -2594
rect 529 -2607 1529 -2594
<< locali >>
rect -1552 2242 -1535 2250
rect -1552 1938 -1535 1946
rect -523 2242 -506 2250
rect -523 1938 -506 1946
rect 506 2242 523 2250
rect 506 1938 523 1946
rect 1535 2242 1552 2250
rect 1535 1938 1552 1946
rect -1552 1195 -1535 1203
rect -1552 891 -1535 899
rect -523 1195 -506 1203
rect -523 891 -506 899
rect 506 1195 523 1203
rect 506 891 523 899
rect 1535 1195 1552 1203
rect 1535 891 1552 899
rect -1552 148 -1535 156
rect -1552 -156 -1535 -148
rect -523 148 -506 156
rect -523 -156 -506 -148
rect 506 148 523 156
rect 506 -156 523 -148
rect 1535 148 1552 156
rect 1535 -156 1552 -148
rect -1552 -899 -1535 -891
rect -1552 -1203 -1535 -1195
rect -523 -899 -506 -891
rect -523 -1203 -506 -1195
rect 506 -899 523 -891
rect 506 -1203 523 -1195
rect 1535 -899 1552 -891
rect 1535 -1203 1552 -1195
rect -1552 -1946 -1535 -1938
rect -1552 -2250 -1535 -2242
rect -523 -1946 -506 -1938
rect -523 -2250 -506 -2242
rect 506 -1946 523 -1938
rect 506 -2250 523 -2242
rect 1535 -1946 1552 -1938
rect 1535 -2250 1552 -2242
<< viali >>
rect -1552 1946 -1535 2242
rect -523 1946 -506 2242
rect 506 1946 523 2242
rect 1535 1946 1552 2242
rect -1552 899 -1535 1195
rect -523 899 -506 1195
rect 506 899 523 1195
rect 1535 899 1552 1195
rect -1552 -148 -1535 148
rect -523 -148 -506 148
rect 506 -148 523 148
rect 1535 -148 1552 148
rect -1552 -1195 -1535 -899
rect -523 -1195 -506 -899
rect 506 -1195 523 -899
rect 1535 -1195 1552 -899
rect -1552 -2242 -1535 -1946
rect -523 -2242 -506 -1946
rect 506 -2242 523 -1946
rect 1535 -2242 1552 -1946
<< metal1 >>
rect -1555 2242 -1532 2248
rect -1555 1946 -1552 2242
rect -1535 1946 -1532 2242
rect -1555 1940 -1532 1946
rect -526 2242 -503 2248
rect -526 1946 -523 2242
rect -506 1946 -503 2242
rect -526 1940 -503 1946
rect 503 2242 526 2248
rect 503 1946 506 2242
rect 523 1946 526 2242
rect 503 1940 526 1946
rect 1532 2242 1555 2248
rect 1532 1946 1535 2242
rect 1552 1946 1555 2242
rect 1532 1940 1555 1946
rect -1555 1195 -1532 1201
rect -1555 899 -1552 1195
rect -1535 899 -1532 1195
rect -1555 893 -1532 899
rect -526 1195 -503 1201
rect -526 899 -523 1195
rect -506 899 -503 1195
rect -526 893 -503 899
rect 503 1195 526 1201
rect 503 899 506 1195
rect 523 899 526 1195
rect 503 893 526 899
rect 1532 1195 1555 1201
rect 1532 899 1535 1195
rect 1552 899 1555 1195
rect 1532 893 1555 899
rect -1555 148 -1532 154
rect -1555 -148 -1552 148
rect -1535 -148 -1532 148
rect -1555 -154 -1532 -148
rect -526 148 -503 154
rect -526 -148 -523 148
rect -506 -148 -503 148
rect -526 -154 -503 -148
rect 503 148 526 154
rect 503 -148 506 148
rect 523 -148 526 148
rect 503 -154 526 -148
rect 1532 148 1555 154
rect 1532 -148 1535 148
rect 1552 -148 1555 148
rect 1532 -154 1555 -148
rect -1555 -899 -1532 -893
rect -1555 -1195 -1552 -899
rect -1535 -1195 -1532 -899
rect -1555 -1201 -1532 -1195
rect -526 -899 -503 -893
rect -526 -1195 -523 -899
rect -506 -1195 -503 -899
rect -526 -1201 -503 -1195
rect 503 -899 526 -893
rect 503 -1195 506 -899
rect 523 -1195 526 -899
rect 503 -1201 526 -1195
rect 1532 -899 1555 -893
rect 1532 -1195 1535 -899
rect 1552 -1195 1555 -899
rect 1532 -1201 1555 -1195
rect -1555 -1946 -1532 -1940
rect -1555 -2242 -1552 -1946
rect -1535 -2242 -1532 -1946
rect -1555 -2248 -1532 -2242
rect -526 -1946 -503 -1940
rect -526 -2242 -523 -1946
rect -506 -2242 -503 -1946
rect -526 -2248 -503 -2242
rect 503 -1946 526 -1940
rect 503 -2242 506 -1946
rect 523 -2242 526 -1946
rect 503 -2248 526 -2242
rect 1532 -1946 1555 -1940
rect 1532 -2242 1535 -1946
rect 1552 -2242 1555 -1946
rect 1532 -2248 1555 -2242
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string parameters w 10 l 10 m 5 nf 3 diffcov 30 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 30 viadrn 30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
