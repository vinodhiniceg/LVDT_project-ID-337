magic
tech sky130A
magscale 1 2
timestamp 1634119395
<< error_p >>
rect -2727 709 2727 713
rect -2727 -709 -2697 709
rect -2661 643 2661 647
rect -2661 47 -2631 643
rect 2631 47 2661 643
rect -2661 -643 -2631 -47
rect 2631 -643 2661 -47
rect -2661 -647 2661 -643
rect 2697 -709 2727 709
rect -2727 -713 2727 -709
<< nwell >>
rect -2697 -709 2697 709
<< mvpmos >>
rect -2603 47 -2003 647
rect -1945 47 -1345 647
rect -1287 47 -687 647
rect -629 47 -29 647
rect 29 47 629 647
rect 687 47 1287 647
rect 1345 47 1945 647
rect 2003 47 2603 647
rect -2603 -647 -2003 -47
rect -1945 -647 -1345 -47
rect -1287 -647 -687 -47
rect -629 -647 -29 -47
rect 29 -647 629 -47
rect 687 -647 1287 -47
rect 1345 -647 1945 -47
rect 2003 -647 2603 -47
<< mvpdiff >>
rect -2661 433 -2603 647
rect -2661 261 -2649 433
rect -2615 261 -2603 433
rect -2661 47 -2603 261
rect -2003 433 -1945 647
rect -2003 261 -1991 433
rect -1957 261 -1945 433
rect -2003 47 -1945 261
rect -1345 433 -1287 647
rect -1345 261 -1333 433
rect -1299 261 -1287 433
rect -1345 47 -1287 261
rect -687 433 -629 647
rect -687 261 -675 433
rect -641 261 -629 433
rect -687 47 -629 261
rect -29 433 29 647
rect -29 261 -17 433
rect 17 261 29 433
rect -29 47 29 261
rect 629 433 687 647
rect 629 261 641 433
rect 675 261 687 433
rect 629 47 687 261
rect 1287 433 1345 647
rect 1287 261 1299 433
rect 1333 261 1345 433
rect 1287 47 1345 261
rect 1945 433 2003 647
rect 1945 261 1957 433
rect 1991 261 2003 433
rect 1945 47 2003 261
rect 2603 433 2661 647
rect 2603 261 2615 433
rect 2649 261 2661 433
rect 2603 47 2661 261
rect -2661 -261 -2603 -47
rect -2661 -433 -2649 -261
rect -2615 -433 -2603 -261
rect -2661 -647 -2603 -433
rect -2003 -261 -1945 -47
rect -2003 -433 -1991 -261
rect -1957 -433 -1945 -261
rect -2003 -647 -1945 -433
rect -1345 -261 -1287 -47
rect -1345 -433 -1333 -261
rect -1299 -433 -1287 -261
rect -1345 -647 -1287 -433
rect -687 -261 -629 -47
rect -687 -433 -675 -261
rect -641 -433 -629 -261
rect -687 -647 -629 -433
rect -29 -261 29 -47
rect -29 -433 -17 -261
rect 17 -433 29 -261
rect -29 -647 29 -433
rect 629 -261 687 -47
rect 629 -433 641 -261
rect 675 -433 687 -261
rect 629 -647 687 -433
rect 1287 -261 1345 -47
rect 1287 -433 1299 -261
rect 1333 -433 1345 -261
rect 1287 -647 1345 -433
rect 1945 -261 2003 -47
rect 1945 -433 1957 -261
rect 1991 -433 2003 -261
rect 1945 -647 2003 -433
rect 2603 -261 2661 -47
rect 2603 -433 2615 -261
rect 2649 -433 2661 -261
rect 2603 -647 2661 -433
<< mvpdiffc >>
rect -2649 261 -2615 433
rect -1991 261 -1957 433
rect -1333 261 -1299 433
rect -675 261 -641 433
rect -17 261 17 433
rect 641 261 675 433
rect 1299 261 1333 433
rect 1957 261 1991 433
rect 2615 261 2649 433
rect -2649 -433 -2615 -261
rect -1991 -433 -1957 -261
rect -1333 -433 -1299 -261
rect -675 -433 -641 -261
rect -17 -433 17 -261
rect 641 -433 675 -261
rect 1299 -433 1333 -261
rect 1957 -433 1991 -261
rect 2615 -433 2649 -261
<< poly >>
rect -2603 647 -2003 673
rect -1945 647 -1345 673
rect -1287 647 -687 673
rect -629 647 -29 673
rect 29 647 629 673
rect 687 647 1287 673
rect 1345 647 1945 673
rect 2003 647 2603 673
rect -2603 21 -2003 47
rect -1945 21 -1345 47
rect -1287 21 -687 47
rect -629 21 -29 47
rect 29 21 629 47
rect 687 21 1287 47
rect 1345 21 1945 47
rect 2003 21 2603 47
rect -2603 -47 -2003 -21
rect -1945 -47 -1345 -21
rect -1287 -47 -687 -21
rect -629 -47 -29 -21
rect 29 -47 629 -21
rect 687 -47 1287 -21
rect 1345 -47 1945 -21
rect 2003 -47 2603 -21
rect -2603 -673 -2003 -647
rect -1945 -673 -1345 -647
rect -1287 -673 -687 -647
rect -629 -673 -29 -647
rect 29 -673 629 -647
rect 687 -673 1287 -647
rect 1345 -673 1945 -647
rect 2003 -673 2603 -647
<< locali >>
rect -2649 433 -2615 449
rect -2649 245 -2615 261
rect -1991 433 -1957 449
rect -1991 245 -1957 261
rect -1333 433 -1299 449
rect -1333 245 -1299 261
rect -675 433 -641 449
rect -675 245 -641 261
rect -17 433 17 449
rect -17 245 17 261
rect 641 433 675 449
rect 641 245 675 261
rect 1299 433 1333 449
rect 1299 245 1333 261
rect 1957 433 1991 449
rect 1957 245 1991 261
rect 2615 433 2649 449
rect 2615 245 2649 261
rect -2649 -261 -2615 -245
rect -2649 -449 -2615 -433
rect -1991 -261 -1957 -245
rect -1991 -449 -1957 -433
rect -1333 -261 -1299 -245
rect -1333 -449 -1299 -433
rect -675 -261 -641 -245
rect -675 -449 -641 -433
rect -17 -261 17 -245
rect -17 -449 17 -433
rect 641 -261 675 -245
rect 641 -449 675 -433
rect 1299 -261 1333 -245
rect 1299 -449 1333 -433
rect 1957 -261 1991 -245
rect 1957 -449 1991 -433
rect 2615 -261 2649 -245
rect 2615 -449 2649 -433
<< viali >>
rect -2649 261 -2615 433
rect -1991 261 -1957 433
rect -1333 261 -1299 433
rect -675 261 -641 433
rect -17 261 17 433
rect 641 261 675 433
rect 1299 261 1333 433
rect 1957 261 1991 433
rect 2615 261 2649 433
rect -2649 -433 -2615 -261
rect -1991 -433 -1957 -261
rect -1333 -433 -1299 -261
rect -675 -433 -641 -261
rect -17 -433 17 -261
rect 641 -433 675 -261
rect 1299 -433 1333 -261
rect 1957 -433 1991 -261
rect 2615 -433 2649 -261
<< metal1 >>
rect -2655 433 -2609 445
rect -2655 261 -2649 433
rect -2615 261 -2609 433
rect -2655 249 -2609 261
rect -1997 433 -1951 445
rect -1997 261 -1991 433
rect -1957 261 -1951 433
rect -1997 249 -1951 261
rect -1339 433 -1293 445
rect -1339 261 -1333 433
rect -1299 261 -1293 433
rect -1339 249 -1293 261
rect -681 433 -635 445
rect -681 261 -675 433
rect -641 261 -635 433
rect -681 249 -635 261
rect -23 433 23 445
rect -23 261 -17 433
rect 17 261 23 433
rect -23 249 23 261
rect 635 433 681 445
rect 635 261 641 433
rect 675 261 681 433
rect 635 249 681 261
rect 1293 433 1339 445
rect 1293 261 1299 433
rect 1333 261 1339 433
rect 1293 249 1339 261
rect 1951 433 1997 445
rect 1951 261 1957 433
rect 1991 261 1997 433
rect 1951 249 1997 261
rect 2609 433 2655 445
rect 2609 261 2615 433
rect 2649 261 2655 433
rect 2609 249 2655 261
rect -2655 -261 -2609 -249
rect -2655 -433 -2649 -261
rect -2615 -433 -2609 -261
rect -2655 -445 -2609 -433
rect -1997 -261 -1951 -249
rect -1997 -433 -1991 -261
rect -1957 -433 -1951 -261
rect -1997 -445 -1951 -433
rect -1339 -261 -1293 -249
rect -1339 -433 -1333 -261
rect -1299 -433 -1293 -261
rect -1339 -445 -1293 -433
rect -681 -261 -635 -249
rect -681 -433 -675 -261
rect -641 -433 -635 -261
rect -681 -445 -635 -433
rect -23 -261 23 -249
rect -23 -433 -17 -261
rect 17 -433 23 -261
rect -23 -445 23 -433
rect 635 -261 681 -249
rect 635 -433 641 -261
rect 675 -433 681 -261
rect 635 -445 681 -433
rect 1293 -261 1339 -249
rect 1293 -433 1299 -261
rect 1333 -433 1339 -261
rect 1293 -445 1339 -433
rect 1951 -261 1997 -249
rect 1951 -433 1957 -261
rect 1991 -433 1997 -261
rect 1951 -445 1997 -433
rect 2609 -261 2655 -249
rect 2609 -433 2615 -261
rect 2649 -433 2655 -261
rect 2609 -445 2655 -433
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string parameters w 3 l 3 m 2 nf 8 diffcov 30 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 30 viadrn 30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
