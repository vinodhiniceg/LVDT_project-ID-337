magic
tech sky130A
timestamp 1634629898
<< error_p >>
rect -54 -50 -25 50
rect 25 -50 54 50
<< mvnmos >>
rect -25 -50 25 50
<< mvndiff >>
rect -54 13 -25 50
rect -54 -13 -48 13
rect -31 -13 -25 13
rect -54 -50 -25 -13
rect 25 13 54 50
rect 25 -13 31 13
rect 48 -13 54 13
rect 25 -50 54 -13
<< mvndiffc >>
rect -48 -13 -31 13
rect 31 -13 48 13
<< poly >>
rect -25 50 25 63
rect -25 -63 25 -50
<< locali >>
rect -48 13 -31 21
rect -48 -21 -31 -13
rect 31 13 48 21
rect 31 -21 48 -13
<< viali >>
rect -48 -13 -31 13
rect 31 -13 48 13
<< metal1 >>
rect -51 13 -28 19
rect -51 -13 -48 13
rect -31 -13 -28 13
rect -51 -19 -28 -13
rect 28 13 51 19
rect 28 -13 31 13
rect 48 -13 51 13
rect 28 -19 51 -13
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string parameters w 1 l 0.5 m 1 nf 1 diffcov 30 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 30 viadrn 30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
