magic
tech sky130A
magscale 1 2
timestamp 1634229043
<< error_s >>
rect -46 3204 -10 3210
rect -12 3170 -10 3176
<< mvpsubdiff >>
rect -450 3050 -266 3090
rect -450 520 -432 3050
rect -302 520 -266 3050
rect -450 486 -266 520
<< mvpsubdiffcont >>
rect -432 520 -302 3050
<< poly >>
rect 476 3422 852 3478
rect 110 2718 574 2790
rect 850 2716 1314 2788
rect 152 2026 616 2098
rect 862 2022 1284 2094
rect 146 1332 610 1404
rect 742 1328 1234 1410
rect 168 640 632 712
rect 786 638 1122 706
<< locali >>
rect -100 3358 26 3432
rect -100 3356 68 3358
rect -100 3354 1382 3356
rect -100 3310 1386 3354
rect -100 3290 68 3310
rect -100 3204 62 3290
rect -10 3176 62 3204
rect -12 3114 66 3176
rect -450 3050 -266 3090
rect -450 520 -432 3050
rect -302 520 -266 3050
rect -450 486 -266 520
rect -2 316 64 3114
rect 650 376 716 3160
rect 1314 3142 1386 3310
rect 1314 2098 1380 3142
rect 1320 2016 1374 2098
rect 1314 1438 1380 2016
rect 1314 1314 1382 1438
rect 640 306 754 376
rect 1314 352 1380 1314
rect 604 110 784 306
<< viali >>
rect -420 602 -338 3004
<< metal1 >>
rect -450 3004 -266 3090
rect -450 602 -420 3004
rect -338 602 -266 3004
rect -450 486 -266 602
use sky130_fd_pr__nfet_g5v0d10v5_QWZYNS  sky130_fd_pr__nfet_g5v0d10v5_QWZYNS_0
timestamp 1634228860
transform 1 0 687 0 1 1714
box -687 -1714 687 1714
<< labels >>
flabel poly 650 3452 650 3452 0 FreeSans 1600 0 0 0 g
flabel locali -64 3306 -64 3306 0 FreeSans 1600 0 0 0 s
flabel locali 696 176 696 176 0 FreeSans 1600 0 0 0 d
<< end >>
