magic
tech sky130A
magscale 1 2
timestamp 1634929801
<< nwell >>
rect -1632 3426 738 3622
rect -1642 3382 738 3426
rect -1642 1848 734 3382
rect -1642 -88 1654 1848
<< pwell >>
rect -2456 5006 -1748 5010
rect -2684 4986 -1692 5006
rect -2684 -134 -1674 4986
rect 1022 3556 2004 3562
rect 850 3548 2004 3556
rect 2256 3548 2882 3572
rect 850 1908 2882 3548
rect 1684 -102 2882 1908
rect 2256 -124 2882 -102
rect -2456 -144 -1674 -134
<< mvnmos >>
rect -2316 4638 -2116 4838
rect -2058 4638 -1858 4838
rect -2316 4344 -2116 4544
rect -2058 4344 -1858 4544
rect -2316 4050 -2116 4250
rect -2058 4050 -1858 4250
rect -2316 3756 -2116 3956
rect -2058 3756 -1858 3956
rect -2316 3462 -2116 3662
rect -2058 3462 -1858 3662
rect -2316 3168 -2116 3368
rect -2058 3168 -1858 3368
rect -2316 2874 -2116 3074
rect -2058 2874 -1858 3074
rect 1146 3134 1346 3334
rect 1404 3134 1604 3334
rect -2316 2580 -2116 2780
rect -2058 2580 -1858 2780
rect 1146 2840 1346 3040
rect 1404 2840 1604 3040
rect -2316 2286 -2116 2486
rect -2058 2286 -1858 2486
rect 1146 2546 1346 2746
rect 1404 2546 1604 2746
rect -2316 1992 -2116 2192
rect -2058 1992 -1858 2192
rect 1146 2252 1346 2452
rect 1404 2252 1604 2452
rect -2316 1698 -2116 1898
rect -2058 1698 -1858 1898
rect 1146 1958 1346 2158
rect 1404 1958 1604 2158
rect -2316 1404 -2116 1604
rect -2058 1404 -1858 1604
rect -2316 1110 -2116 1310
rect -2058 1110 -1858 1310
rect 1804 1210 2004 1410
rect 2062 1210 2262 1410
rect -2316 816 -2116 1016
rect -2058 816 -1858 1016
rect -2316 522 -2116 722
rect -2058 522 -1858 722
rect -2316 228 -2116 428
rect -2058 228 -1858 428
rect -2316 -66 -2116 134
rect -2058 -66 -1858 134
rect 1804 916 2004 1116
rect 2062 916 2262 1116
rect 1804 622 2004 822
rect 2062 622 2262 822
rect 1804 328 2004 528
rect 2062 328 2262 528
rect 1804 34 2004 234
rect 2062 34 2262 234
<< mvpmos >>
rect 108 3024 308 3224
rect 366 3024 566 3224
rect -1404 2696 -1204 2896
rect -1146 2696 -946 2896
rect -888 2696 -688 2896
rect -630 2696 -430 2896
rect 108 2730 308 2930
rect 366 2730 566 2930
rect -1404 2402 -1204 2602
rect -1146 2402 -946 2602
rect -888 2402 -688 2602
rect -630 2402 -430 2602
rect 108 2436 308 2636
rect 366 2436 566 2636
rect -1404 2108 -1204 2308
rect -1146 2108 -946 2308
rect -888 2108 -688 2308
rect -630 2108 -430 2308
rect 108 2142 308 2342
rect 366 2142 566 2342
rect -1404 1814 -1204 2014
rect -1146 1814 -946 2014
rect -888 1814 -688 2014
rect -630 1814 -430 2014
rect 108 1848 308 2048
rect 366 1848 566 2048
rect -1404 1520 -1204 1720
rect -1146 1520 -946 1720
rect -888 1520 -688 1720
rect -630 1520 -430 1720
rect -1404 1226 -1204 1426
rect -1146 1226 -946 1426
rect -888 1226 -688 1426
rect -630 1226 -430 1426
rect 108 1224 308 1424
rect 366 1224 566 1424
rect 896 1222 1096 1422
rect 1154 1222 1354 1422
rect -1404 932 -1204 1132
rect -1146 932 -946 1132
rect -888 932 -688 1132
rect -630 932 -430 1132
rect 108 930 308 1130
rect 366 930 566 1130
rect 896 928 1096 1128
rect 1154 928 1354 1128
rect -1404 638 -1204 838
rect -1146 638 -946 838
rect -888 638 -688 838
rect -630 638 -430 838
rect 108 636 308 836
rect 366 636 566 836
rect 896 634 1096 834
rect 1154 634 1354 834
rect -1404 344 -1204 544
rect -1146 344 -946 544
rect -888 344 -688 544
rect -630 344 -430 544
rect 108 342 308 542
rect 366 342 566 542
rect 896 340 1096 540
rect 1154 340 1354 540
rect -1404 50 -1204 250
rect -1146 50 -946 250
rect -888 50 -688 250
rect -630 50 -430 250
rect 108 48 308 248
rect 366 48 566 248
rect 896 46 1096 246
rect 1154 46 1354 246
<< mvndiff >>
rect -2374 4764 -2316 4838
rect -2374 4712 -2362 4764
rect -2328 4712 -2316 4764
rect -2374 4638 -2316 4712
rect -2116 4764 -2058 4838
rect -2116 4712 -2104 4764
rect -2070 4712 -2058 4764
rect -2116 4638 -2058 4712
rect -1858 4764 -1800 4838
rect -1858 4712 -1846 4764
rect -1812 4712 -1800 4764
rect -1858 4638 -1800 4712
rect -2374 4470 -2316 4544
rect -2374 4418 -2362 4470
rect -2328 4418 -2316 4470
rect -2374 4344 -2316 4418
rect -2116 4470 -2058 4544
rect -2116 4418 -2104 4470
rect -2070 4418 -2058 4470
rect -2116 4344 -2058 4418
rect -1858 4470 -1800 4544
rect -1858 4418 -1846 4470
rect -1812 4418 -1800 4470
rect -1858 4344 -1800 4418
rect -2374 4176 -2316 4250
rect -2374 4124 -2362 4176
rect -2328 4124 -2316 4176
rect -2374 4050 -2316 4124
rect -2116 4176 -2058 4250
rect -2116 4124 -2104 4176
rect -2070 4124 -2058 4176
rect -2116 4050 -2058 4124
rect -1858 4176 -1800 4250
rect -1858 4124 -1846 4176
rect -1812 4124 -1800 4176
rect -1858 4050 -1800 4124
rect -2374 3882 -2316 3956
rect -2374 3830 -2362 3882
rect -2328 3830 -2316 3882
rect -2374 3756 -2316 3830
rect -2116 3882 -2058 3956
rect -2116 3830 -2104 3882
rect -2070 3830 -2058 3882
rect -2116 3756 -2058 3830
rect -1858 3882 -1800 3956
rect -1858 3830 -1846 3882
rect -1812 3830 -1800 3882
rect -1858 3756 -1800 3830
rect -2374 3588 -2316 3662
rect -2374 3536 -2362 3588
rect -2328 3536 -2316 3588
rect -2374 3462 -2316 3536
rect -2116 3588 -2058 3662
rect -2116 3536 -2104 3588
rect -2070 3536 -2058 3588
rect -2116 3462 -2058 3536
rect -1858 3588 -1800 3662
rect -1858 3536 -1846 3588
rect -1812 3536 -1800 3588
rect -1858 3462 -1800 3536
rect -2374 3294 -2316 3368
rect -2374 3242 -2362 3294
rect -2328 3242 -2316 3294
rect -2374 3168 -2316 3242
rect -2116 3294 -2058 3368
rect -2116 3242 -2104 3294
rect -2070 3242 -2058 3294
rect -2116 3168 -2058 3242
rect -1858 3294 -1800 3368
rect -1858 3242 -1846 3294
rect -1812 3242 -1800 3294
rect -1858 3168 -1800 3242
rect -2374 3000 -2316 3074
rect -2374 2948 -2362 3000
rect -2328 2948 -2316 3000
rect -2374 2874 -2316 2948
rect -2116 3000 -2058 3074
rect -2116 2948 -2104 3000
rect -2070 2948 -2058 3000
rect -2116 2874 -2058 2948
rect -1858 3000 -1800 3074
rect 1088 3260 1146 3334
rect 1088 3208 1100 3260
rect 1134 3208 1146 3260
rect 1088 3134 1146 3208
rect 1346 3260 1404 3334
rect 1346 3208 1358 3260
rect 1392 3208 1404 3260
rect 1346 3134 1404 3208
rect 1604 3260 1662 3334
rect 1604 3208 1616 3260
rect 1650 3208 1662 3260
rect 1604 3134 1662 3208
rect -1858 2948 -1846 3000
rect -1812 2948 -1800 3000
rect 1088 2966 1146 3040
rect -1858 2874 -1800 2948
rect -2374 2706 -2316 2780
rect -2374 2654 -2362 2706
rect -2328 2654 -2316 2706
rect -2374 2580 -2316 2654
rect -2116 2706 -2058 2780
rect -2116 2654 -2104 2706
rect -2070 2654 -2058 2706
rect -2116 2580 -2058 2654
rect -1858 2706 -1800 2780
rect -1858 2654 -1846 2706
rect -1812 2654 -1800 2706
rect 1088 2914 1100 2966
rect 1134 2914 1146 2966
rect 1088 2840 1146 2914
rect 1346 2966 1404 3040
rect 1346 2914 1358 2966
rect 1392 2914 1404 2966
rect 1346 2840 1404 2914
rect 1604 2966 1662 3040
rect 1604 2914 1616 2966
rect 1650 2914 1662 2966
rect 1604 2840 1662 2914
rect -1858 2580 -1800 2654
rect 1088 2672 1146 2746
rect -2374 2412 -2316 2486
rect -2374 2360 -2362 2412
rect -2328 2360 -2316 2412
rect -2374 2286 -2316 2360
rect -2116 2412 -2058 2486
rect -2116 2360 -2104 2412
rect -2070 2360 -2058 2412
rect -2116 2286 -2058 2360
rect -1858 2412 -1800 2486
rect -1858 2360 -1846 2412
rect -1812 2360 -1800 2412
rect 1088 2620 1100 2672
rect 1134 2620 1146 2672
rect 1088 2546 1146 2620
rect 1346 2672 1404 2746
rect 1346 2620 1358 2672
rect 1392 2620 1404 2672
rect 1346 2546 1404 2620
rect 1604 2672 1662 2746
rect 1604 2620 1616 2672
rect 1650 2620 1662 2672
rect 1604 2546 1662 2620
rect -1858 2286 -1800 2360
rect 1088 2378 1146 2452
rect -2374 2118 -2316 2192
rect -2374 2066 -2362 2118
rect -2328 2066 -2316 2118
rect -2374 1992 -2316 2066
rect -2116 2118 -2058 2192
rect -2116 2066 -2104 2118
rect -2070 2066 -2058 2118
rect -2116 1992 -2058 2066
rect -1858 2118 -1800 2192
rect -1858 2066 -1846 2118
rect -1812 2066 -1800 2118
rect 1088 2326 1100 2378
rect 1134 2326 1146 2378
rect 1088 2252 1146 2326
rect 1346 2378 1404 2452
rect 1346 2326 1358 2378
rect 1392 2326 1404 2378
rect 1346 2252 1404 2326
rect 1604 2378 1662 2452
rect 1604 2326 1616 2378
rect 1650 2326 1662 2378
rect 1604 2252 1662 2326
rect -1858 1992 -1800 2066
rect 1088 2084 1146 2158
rect -2374 1824 -2316 1898
rect -2374 1772 -2362 1824
rect -2328 1772 -2316 1824
rect -2374 1698 -2316 1772
rect -2116 1824 -2058 1898
rect -2116 1772 -2104 1824
rect -2070 1772 -2058 1824
rect -2116 1698 -2058 1772
rect -1858 1824 -1800 1898
rect -1858 1772 -1846 1824
rect -1812 1772 -1800 1824
rect 1088 2032 1100 2084
rect 1134 2032 1146 2084
rect 1088 1958 1146 2032
rect 1346 2084 1404 2158
rect 1346 2032 1358 2084
rect 1392 2032 1404 2084
rect 1346 1958 1404 2032
rect 1604 2084 1662 2158
rect 1604 2032 1616 2084
rect 1650 2032 1662 2084
rect 1604 1958 1662 2032
rect -1858 1698 -1800 1772
rect -2374 1530 -2316 1604
rect -2374 1478 -2362 1530
rect -2328 1478 -2316 1530
rect -2374 1404 -2316 1478
rect -2116 1530 -2058 1604
rect -2116 1478 -2104 1530
rect -2070 1478 -2058 1530
rect -2116 1404 -2058 1478
rect -1858 1530 -1800 1604
rect -1858 1478 -1846 1530
rect -1812 1478 -1800 1530
rect -1858 1404 -1800 1478
rect -2374 1236 -2316 1310
rect -2374 1184 -2362 1236
rect -2328 1184 -2316 1236
rect -2374 1110 -2316 1184
rect -2116 1236 -2058 1310
rect -2116 1184 -2104 1236
rect -2070 1184 -2058 1236
rect -2116 1110 -2058 1184
rect -1858 1236 -1800 1310
rect -1858 1184 -1846 1236
rect -1812 1184 -1800 1236
rect -1858 1110 -1800 1184
rect 1746 1336 1804 1410
rect 1746 1284 1758 1336
rect 1792 1284 1804 1336
rect 1746 1210 1804 1284
rect 2004 1336 2062 1410
rect 2004 1284 2016 1336
rect 2050 1284 2062 1336
rect 2004 1210 2062 1284
rect 2262 1336 2320 1410
rect 2262 1284 2274 1336
rect 2308 1284 2320 1336
rect 2262 1210 2320 1284
rect -2374 942 -2316 1016
rect -2374 890 -2362 942
rect -2328 890 -2316 942
rect -2374 816 -2316 890
rect -2116 942 -2058 1016
rect -2116 890 -2104 942
rect -2070 890 -2058 942
rect -2116 816 -2058 890
rect -1858 942 -1800 1016
rect -1858 890 -1846 942
rect -1812 890 -1800 942
rect -1858 816 -1800 890
rect 1746 1042 1804 1116
rect -2374 648 -2316 722
rect -2374 596 -2362 648
rect -2328 596 -2316 648
rect -2374 522 -2316 596
rect -2116 648 -2058 722
rect -2116 596 -2104 648
rect -2070 596 -2058 648
rect -2116 522 -2058 596
rect -1858 648 -1800 722
rect -1858 596 -1846 648
rect -1812 596 -1800 648
rect -1858 522 -1800 596
rect -2374 354 -2316 428
rect -2374 302 -2362 354
rect -2328 302 -2316 354
rect -2374 228 -2316 302
rect -2116 354 -2058 428
rect -2116 302 -2104 354
rect -2070 302 -2058 354
rect -2116 228 -2058 302
rect -1858 354 -1800 428
rect -1858 302 -1846 354
rect -1812 302 -1800 354
rect -1858 228 -1800 302
rect -2374 60 -2316 134
rect -2374 8 -2362 60
rect -2328 8 -2316 60
rect -2374 -66 -2316 8
rect -2116 60 -2058 134
rect -2116 8 -2104 60
rect -2070 8 -2058 60
rect -2116 -66 -2058 8
rect -1858 60 -1800 134
rect -1858 8 -1846 60
rect -1812 8 -1800 60
rect 1746 990 1758 1042
rect 1792 990 1804 1042
rect 1746 916 1804 990
rect 2004 1042 2062 1116
rect 2004 990 2016 1042
rect 2050 990 2062 1042
rect 2004 916 2062 990
rect 2262 1042 2320 1116
rect 2262 990 2274 1042
rect 2308 990 2320 1042
rect 2262 916 2320 990
rect 1746 748 1804 822
rect 1746 696 1758 748
rect 1792 696 1804 748
rect 1746 622 1804 696
rect 2004 748 2062 822
rect 2004 696 2016 748
rect 2050 696 2062 748
rect 2004 622 2062 696
rect 2262 748 2320 822
rect 2262 696 2274 748
rect 2308 696 2320 748
rect 2262 622 2320 696
rect 1746 454 1804 528
rect 1746 402 1758 454
rect 1792 402 1804 454
rect 1746 328 1804 402
rect 2004 454 2062 528
rect 2004 402 2016 454
rect 2050 402 2062 454
rect 2004 328 2062 402
rect 2262 454 2320 528
rect 2262 402 2274 454
rect 2308 402 2320 454
rect 2262 328 2320 402
rect 1746 160 1804 234
rect 1746 108 1758 160
rect 1792 108 1804 160
rect -1858 -66 -1800 8
rect 1746 34 1804 108
rect 2004 160 2062 234
rect 2004 108 2016 160
rect 2050 108 2062 160
rect 2004 34 2062 108
rect 2262 160 2320 234
rect 2262 108 2274 160
rect 2308 108 2320 160
rect 2262 34 2320 108
<< mvpdiff >>
rect 50 3150 108 3224
rect 50 3098 62 3150
rect 96 3098 108 3150
rect 50 3024 108 3098
rect 308 3150 366 3224
rect 308 3098 320 3150
rect 354 3098 366 3150
rect 308 3024 366 3098
rect 566 3150 624 3224
rect 566 3098 578 3150
rect 612 3098 624 3150
rect 566 3024 624 3098
rect -1462 2822 -1404 2896
rect -1462 2770 -1450 2822
rect -1416 2770 -1404 2822
rect -1462 2696 -1404 2770
rect -1204 2822 -1146 2896
rect -1204 2770 -1192 2822
rect -1158 2770 -1146 2822
rect -1204 2696 -1146 2770
rect -946 2822 -888 2896
rect -946 2770 -934 2822
rect -900 2770 -888 2822
rect -946 2696 -888 2770
rect -688 2822 -630 2896
rect -688 2770 -676 2822
rect -642 2770 -630 2822
rect -688 2696 -630 2770
rect -430 2822 -372 2896
rect -430 2770 -418 2822
rect -384 2770 -372 2822
rect -430 2696 -372 2770
rect 50 2856 108 2930
rect 50 2804 62 2856
rect 96 2804 108 2856
rect 50 2730 108 2804
rect 308 2856 366 2930
rect 308 2804 320 2856
rect 354 2804 366 2856
rect 308 2730 366 2804
rect 566 2856 624 2930
rect 566 2804 578 2856
rect 612 2804 624 2856
rect 566 2730 624 2804
rect -1462 2528 -1404 2602
rect -1462 2476 -1450 2528
rect -1416 2476 -1404 2528
rect -1462 2402 -1404 2476
rect -1204 2528 -1146 2602
rect -1204 2476 -1192 2528
rect -1158 2476 -1146 2528
rect -1204 2402 -1146 2476
rect -946 2528 -888 2602
rect -946 2476 -934 2528
rect -900 2476 -888 2528
rect -946 2402 -888 2476
rect -688 2528 -630 2602
rect -688 2476 -676 2528
rect -642 2476 -630 2528
rect -688 2402 -630 2476
rect -430 2528 -372 2602
rect -430 2476 -418 2528
rect -384 2476 -372 2528
rect -430 2402 -372 2476
rect 50 2562 108 2636
rect 50 2510 62 2562
rect 96 2510 108 2562
rect 50 2436 108 2510
rect 308 2562 366 2636
rect 308 2510 320 2562
rect 354 2510 366 2562
rect 308 2436 366 2510
rect 566 2562 624 2636
rect 566 2510 578 2562
rect 612 2510 624 2562
rect 566 2436 624 2510
rect -1462 2234 -1404 2308
rect -1462 2182 -1450 2234
rect -1416 2182 -1404 2234
rect -1462 2108 -1404 2182
rect -1204 2234 -1146 2308
rect -1204 2182 -1192 2234
rect -1158 2182 -1146 2234
rect -1204 2108 -1146 2182
rect -946 2234 -888 2308
rect -946 2182 -934 2234
rect -900 2182 -888 2234
rect -946 2108 -888 2182
rect -688 2234 -630 2308
rect -688 2182 -676 2234
rect -642 2182 -630 2234
rect -688 2108 -630 2182
rect -430 2234 -372 2308
rect -430 2182 -418 2234
rect -384 2182 -372 2234
rect -430 2108 -372 2182
rect 50 2268 108 2342
rect 50 2216 62 2268
rect 96 2216 108 2268
rect 50 2142 108 2216
rect 308 2268 366 2342
rect 308 2216 320 2268
rect 354 2216 366 2268
rect 308 2142 366 2216
rect 566 2268 624 2342
rect 566 2216 578 2268
rect 612 2216 624 2268
rect 566 2142 624 2216
rect -1462 1940 -1404 2014
rect -1462 1888 -1450 1940
rect -1416 1888 -1404 1940
rect -1462 1814 -1404 1888
rect -1204 1940 -1146 2014
rect -1204 1888 -1192 1940
rect -1158 1888 -1146 1940
rect -1204 1814 -1146 1888
rect -946 1940 -888 2014
rect -946 1888 -934 1940
rect -900 1888 -888 1940
rect -946 1814 -888 1888
rect -688 1940 -630 2014
rect -688 1888 -676 1940
rect -642 1888 -630 1940
rect -688 1814 -630 1888
rect -430 1940 -372 2014
rect -430 1888 -418 1940
rect -384 1888 -372 1940
rect -430 1814 -372 1888
rect 50 1974 108 2048
rect 50 1922 62 1974
rect 96 1922 108 1974
rect 50 1848 108 1922
rect 308 1974 366 2048
rect 308 1922 320 1974
rect 354 1922 366 1974
rect 308 1848 366 1922
rect 566 1974 624 2048
rect 566 1922 578 1974
rect 612 1922 624 1974
rect 566 1848 624 1922
rect -1462 1646 -1404 1720
rect -1462 1594 -1450 1646
rect -1416 1594 -1404 1646
rect -1462 1520 -1404 1594
rect -1204 1646 -1146 1720
rect -1204 1594 -1192 1646
rect -1158 1594 -1146 1646
rect -1204 1520 -1146 1594
rect -946 1646 -888 1720
rect -946 1594 -934 1646
rect -900 1594 -888 1646
rect -946 1520 -888 1594
rect -688 1646 -630 1720
rect -688 1594 -676 1646
rect -642 1594 -630 1646
rect -688 1520 -630 1594
rect -430 1646 -372 1720
rect -430 1594 -418 1646
rect -384 1594 -372 1646
rect -430 1520 -372 1594
rect -1462 1352 -1404 1426
rect -1462 1300 -1450 1352
rect -1416 1300 -1404 1352
rect -1462 1226 -1404 1300
rect -1204 1352 -1146 1426
rect -1204 1300 -1192 1352
rect -1158 1300 -1146 1352
rect -1204 1226 -1146 1300
rect -946 1352 -888 1426
rect -946 1300 -934 1352
rect -900 1300 -888 1352
rect -946 1226 -888 1300
rect -688 1352 -630 1426
rect -688 1300 -676 1352
rect -642 1300 -630 1352
rect -688 1226 -630 1300
rect -430 1352 -372 1426
rect -430 1300 -418 1352
rect -384 1300 -372 1352
rect -430 1226 -372 1300
rect 50 1350 108 1424
rect 50 1298 62 1350
rect 96 1298 108 1350
rect 50 1224 108 1298
rect 308 1350 366 1424
rect 308 1298 320 1350
rect 354 1298 366 1350
rect 308 1224 366 1298
rect 566 1350 624 1424
rect 566 1298 578 1350
rect 612 1298 624 1350
rect 566 1224 624 1298
rect 838 1348 896 1422
rect 838 1296 850 1348
rect 884 1296 896 1348
rect 838 1222 896 1296
rect 1096 1348 1154 1422
rect 1096 1296 1108 1348
rect 1142 1296 1154 1348
rect 1096 1222 1154 1296
rect 1354 1348 1412 1422
rect 1354 1296 1366 1348
rect 1400 1296 1412 1348
rect 1354 1222 1412 1296
rect -1462 1058 -1404 1132
rect -1462 1006 -1450 1058
rect -1416 1006 -1404 1058
rect -1462 932 -1404 1006
rect -1204 1058 -1146 1132
rect -1204 1006 -1192 1058
rect -1158 1006 -1146 1058
rect -1204 932 -1146 1006
rect -946 1058 -888 1132
rect -946 1006 -934 1058
rect -900 1006 -888 1058
rect -946 932 -888 1006
rect -688 1058 -630 1132
rect -688 1006 -676 1058
rect -642 1006 -630 1058
rect -688 932 -630 1006
rect -430 1058 -372 1132
rect -430 1006 -418 1058
rect -384 1006 -372 1058
rect -430 932 -372 1006
rect 50 1056 108 1130
rect 50 1004 62 1056
rect 96 1004 108 1056
rect 50 930 108 1004
rect 308 1056 366 1130
rect 308 1004 320 1056
rect 354 1004 366 1056
rect 308 930 366 1004
rect 566 1056 624 1130
rect 566 1004 578 1056
rect 612 1004 624 1056
rect 566 930 624 1004
rect 838 1054 896 1128
rect 838 1002 850 1054
rect 884 1002 896 1054
rect 838 928 896 1002
rect 1096 1054 1154 1128
rect 1096 1002 1108 1054
rect 1142 1002 1154 1054
rect 1096 928 1154 1002
rect 1354 1054 1412 1128
rect 1354 1002 1366 1054
rect 1400 1002 1412 1054
rect 1354 928 1412 1002
rect -1462 764 -1404 838
rect -1462 712 -1450 764
rect -1416 712 -1404 764
rect -1462 638 -1404 712
rect -1204 764 -1146 838
rect -1204 712 -1192 764
rect -1158 712 -1146 764
rect -1204 638 -1146 712
rect -946 764 -888 838
rect -946 712 -934 764
rect -900 712 -888 764
rect -946 638 -888 712
rect -688 764 -630 838
rect -688 712 -676 764
rect -642 712 -630 764
rect -688 638 -630 712
rect -430 764 -372 838
rect -430 712 -418 764
rect -384 712 -372 764
rect -430 638 -372 712
rect 50 762 108 836
rect 50 710 62 762
rect 96 710 108 762
rect 50 636 108 710
rect 308 762 366 836
rect 308 710 320 762
rect 354 710 366 762
rect 308 636 366 710
rect 566 762 624 836
rect 566 710 578 762
rect 612 710 624 762
rect 566 636 624 710
rect 838 760 896 834
rect 838 708 850 760
rect 884 708 896 760
rect 838 634 896 708
rect 1096 760 1154 834
rect 1096 708 1108 760
rect 1142 708 1154 760
rect 1096 634 1154 708
rect 1354 760 1412 834
rect 1354 708 1366 760
rect 1400 708 1412 760
rect 1354 634 1412 708
rect -1462 470 -1404 544
rect -1462 418 -1450 470
rect -1416 418 -1404 470
rect -1462 344 -1404 418
rect -1204 470 -1146 544
rect -1204 418 -1192 470
rect -1158 418 -1146 470
rect -1204 344 -1146 418
rect -946 470 -888 544
rect -946 418 -934 470
rect -900 418 -888 470
rect -946 344 -888 418
rect -688 470 -630 544
rect -688 418 -676 470
rect -642 418 -630 470
rect -688 344 -630 418
rect -430 470 -372 544
rect -430 418 -418 470
rect -384 418 -372 470
rect -430 344 -372 418
rect 50 468 108 542
rect 50 416 62 468
rect 96 416 108 468
rect 50 342 108 416
rect 308 468 366 542
rect 308 416 320 468
rect 354 416 366 468
rect 308 342 366 416
rect 566 468 624 542
rect 566 416 578 468
rect 612 416 624 468
rect 566 342 624 416
rect 838 466 896 540
rect 838 414 850 466
rect 884 414 896 466
rect 838 340 896 414
rect 1096 466 1154 540
rect 1096 414 1108 466
rect 1142 414 1154 466
rect 1096 340 1154 414
rect 1354 466 1412 540
rect 1354 414 1366 466
rect 1400 414 1412 466
rect 1354 340 1412 414
rect -1462 176 -1404 250
rect -1462 124 -1450 176
rect -1416 124 -1404 176
rect -1462 50 -1404 124
rect -1204 176 -1146 250
rect -1204 124 -1192 176
rect -1158 124 -1146 176
rect -1204 50 -1146 124
rect -946 176 -888 250
rect -946 124 -934 176
rect -900 124 -888 176
rect -946 50 -888 124
rect -688 176 -630 250
rect -688 124 -676 176
rect -642 124 -630 176
rect -688 50 -630 124
rect -430 176 -372 250
rect -430 124 -418 176
rect -384 124 -372 176
rect -430 50 -372 124
rect 50 174 108 248
rect 50 122 62 174
rect 96 122 108 174
rect 50 48 108 122
rect 308 174 366 248
rect 308 122 320 174
rect 354 122 366 174
rect 308 48 366 122
rect 566 174 624 248
rect 566 122 578 174
rect 612 122 624 174
rect 566 48 624 122
rect 838 172 896 246
rect 838 120 850 172
rect 884 120 896 172
rect 838 46 896 120
rect 1096 172 1154 246
rect 1096 120 1108 172
rect 1142 120 1154 172
rect 1096 46 1154 120
rect 1354 172 1412 246
rect 1354 120 1366 172
rect 1400 120 1412 172
rect 1354 46 1412 120
<< mvndiffc >>
rect -2362 4712 -2328 4764
rect -2104 4712 -2070 4764
rect -1846 4712 -1812 4764
rect -2362 4418 -2328 4470
rect -2104 4418 -2070 4470
rect -1846 4418 -1812 4470
rect -2362 4124 -2328 4176
rect -2104 4124 -2070 4176
rect -1846 4124 -1812 4176
rect -2362 3830 -2328 3882
rect -2104 3830 -2070 3882
rect -1846 3830 -1812 3882
rect -2362 3536 -2328 3588
rect -2104 3536 -2070 3588
rect -1846 3536 -1812 3588
rect -2362 3242 -2328 3294
rect -2104 3242 -2070 3294
rect -1846 3242 -1812 3294
rect -2362 2948 -2328 3000
rect -2104 2948 -2070 3000
rect 1100 3208 1134 3260
rect 1358 3208 1392 3260
rect 1616 3208 1650 3260
rect -1846 2948 -1812 3000
rect -2362 2654 -2328 2706
rect -2104 2654 -2070 2706
rect -1846 2654 -1812 2706
rect 1100 2914 1134 2966
rect 1358 2914 1392 2966
rect 1616 2914 1650 2966
rect -2362 2360 -2328 2412
rect -2104 2360 -2070 2412
rect -1846 2360 -1812 2412
rect 1100 2620 1134 2672
rect 1358 2620 1392 2672
rect 1616 2620 1650 2672
rect -2362 2066 -2328 2118
rect -2104 2066 -2070 2118
rect -1846 2066 -1812 2118
rect 1100 2326 1134 2378
rect 1358 2326 1392 2378
rect 1616 2326 1650 2378
rect -2362 1772 -2328 1824
rect -2104 1772 -2070 1824
rect -1846 1772 -1812 1824
rect 1100 2032 1134 2084
rect 1358 2032 1392 2084
rect 1616 2032 1650 2084
rect -2362 1478 -2328 1530
rect -2104 1478 -2070 1530
rect -1846 1478 -1812 1530
rect -2362 1184 -2328 1236
rect -2104 1184 -2070 1236
rect -1846 1184 -1812 1236
rect 1758 1284 1792 1336
rect 2016 1284 2050 1336
rect 2274 1284 2308 1336
rect -2362 890 -2328 942
rect -2104 890 -2070 942
rect -1846 890 -1812 942
rect -2362 596 -2328 648
rect -2104 596 -2070 648
rect -1846 596 -1812 648
rect -2362 302 -2328 354
rect -2104 302 -2070 354
rect -1846 302 -1812 354
rect -2362 8 -2328 60
rect -2104 8 -2070 60
rect -1846 8 -1812 60
rect 1758 990 1792 1042
rect 2016 990 2050 1042
rect 2274 990 2308 1042
rect 1758 696 1792 748
rect 2016 696 2050 748
rect 2274 696 2308 748
rect 1758 402 1792 454
rect 2016 402 2050 454
rect 2274 402 2308 454
rect 1758 108 1792 160
rect 2016 108 2050 160
rect 2274 108 2308 160
<< mvpdiffc >>
rect 62 3098 96 3150
rect 320 3098 354 3150
rect 578 3098 612 3150
rect -1450 2770 -1416 2822
rect -1192 2770 -1158 2822
rect -934 2770 -900 2822
rect -676 2770 -642 2822
rect -418 2770 -384 2822
rect 62 2804 96 2856
rect 320 2804 354 2856
rect 578 2804 612 2856
rect -1450 2476 -1416 2528
rect -1192 2476 -1158 2528
rect -934 2476 -900 2528
rect -676 2476 -642 2528
rect -418 2476 -384 2528
rect 62 2510 96 2562
rect 320 2510 354 2562
rect 578 2510 612 2562
rect -1450 2182 -1416 2234
rect -1192 2182 -1158 2234
rect -934 2182 -900 2234
rect -676 2182 -642 2234
rect -418 2182 -384 2234
rect 62 2216 96 2268
rect 320 2216 354 2268
rect 578 2216 612 2268
rect -1450 1888 -1416 1940
rect -1192 1888 -1158 1940
rect -934 1888 -900 1940
rect -676 1888 -642 1940
rect -418 1888 -384 1940
rect 62 1922 96 1974
rect 320 1922 354 1974
rect 578 1922 612 1974
rect -1450 1594 -1416 1646
rect -1192 1594 -1158 1646
rect -934 1594 -900 1646
rect -676 1594 -642 1646
rect -418 1594 -384 1646
rect -1450 1300 -1416 1352
rect -1192 1300 -1158 1352
rect -934 1300 -900 1352
rect -676 1300 -642 1352
rect -418 1300 -384 1352
rect 62 1298 96 1350
rect 320 1298 354 1350
rect 578 1298 612 1350
rect 850 1296 884 1348
rect 1108 1296 1142 1348
rect 1366 1296 1400 1348
rect -1450 1006 -1416 1058
rect -1192 1006 -1158 1058
rect -934 1006 -900 1058
rect -676 1006 -642 1058
rect -418 1006 -384 1058
rect 62 1004 96 1056
rect 320 1004 354 1056
rect 578 1004 612 1056
rect 850 1002 884 1054
rect 1108 1002 1142 1054
rect 1366 1002 1400 1054
rect -1450 712 -1416 764
rect -1192 712 -1158 764
rect -934 712 -900 764
rect -676 712 -642 764
rect -418 712 -384 764
rect 62 710 96 762
rect 320 710 354 762
rect 578 710 612 762
rect 850 708 884 760
rect 1108 708 1142 760
rect 1366 708 1400 760
rect -1450 418 -1416 470
rect -1192 418 -1158 470
rect -934 418 -900 470
rect -676 418 -642 470
rect -418 418 -384 470
rect 62 416 96 468
rect 320 416 354 468
rect 578 416 612 468
rect 850 414 884 466
rect 1108 414 1142 466
rect 1366 414 1400 466
rect -1450 124 -1416 176
rect -1192 124 -1158 176
rect -934 124 -900 176
rect -676 124 -642 176
rect -418 124 -384 176
rect 62 122 96 174
rect 320 122 354 174
rect 578 122 612 174
rect 850 120 884 172
rect 1108 120 1142 172
rect 1366 120 1400 172
<< mvpsubdiff >>
rect -2584 2594 -2450 2676
rect -2584 450 -2560 2594
rect -2482 450 -2450 2594
rect 2432 1222 2602 1280
rect -2584 328 -2450 450
rect 2432 190 2456 1222
rect 2554 190 2602 1222
rect 2432 116 2602 190
<< mvnsubdiff >>
rect -398 3376 -124 3426
rect -398 3054 -378 3376
rect -196 3054 -124 3376
rect -398 3004 -124 3054
rect 1480 960 1576 994
rect 1480 238 1492 960
rect 1564 238 1576 960
rect 1480 210 1576 238
<< mvpsubdiffcont >>
rect -2560 450 -2482 2594
rect 2456 190 2554 1222
<< mvnsubdiffcont >>
rect -378 3054 -196 3376
rect 1492 238 1564 960
<< poly >>
rect -2262 5024 -1908 5090
rect -2262 4922 -2180 5024
rect -2024 4922 -1908 5024
rect -2262 4914 -1908 4922
rect -2260 4864 -1916 4914
rect -2316 4854 -1858 4864
rect -2316 4838 -2116 4854
rect -2058 4838 -1858 4854
rect -2316 4612 -2116 4638
rect -2058 4612 -1858 4638
rect -2286 4570 -2152 4612
rect -2010 4570 -1876 4612
rect -2316 4544 -2116 4570
rect -2058 4544 -1858 4570
rect -2316 4318 -2116 4344
rect -2058 4318 -1858 4344
rect -2296 4276 -2162 4318
rect -2030 4276 -1896 4318
rect -2316 4250 -2116 4276
rect -2058 4250 -1858 4276
rect -2316 4024 -2116 4050
rect -2058 4024 -1858 4050
rect -2292 3982 -2158 4024
rect -2012 3982 -1878 4024
rect -2316 3956 -2116 3982
rect -2058 3956 -1858 3982
rect -2316 3730 -2116 3756
rect -2058 3730 -1858 3756
rect -2276 3688 -2142 3730
rect -2010 3688 -1876 3730
rect -2316 3662 -2116 3688
rect -2058 3662 -1858 3688
rect 1238 3514 1542 3690
rect -2316 3436 -2116 3462
rect -2058 3436 -1858 3462
rect -2282 3394 -2148 3436
rect -2012 3394 -1878 3436
rect -2316 3368 -2116 3394
rect -2058 3368 -1858 3394
rect -2316 3142 -2116 3168
rect -2058 3142 -1858 3168
rect -2282 3100 -2148 3142
rect -2032 3100 -1898 3142
rect -2316 3074 -2116 3100
rect -2058 3074 -1858 3100
rect 190 3352 494 3430
rect 1164 3360 1564 3514
rect 1146 3354 1604 3360
rect 184 3250 510 3352
rect 1146 3334 1346 3354
rect 1404 3334 1604 3354
rect 108 3244 566 3250
rect 108 3224 308 3244
rect 366 3224 566 3244
rect 1146 3108 1346 3134
rect 1404 3108 1604 3134
rect 1166 3066 1302 3108
rect 1442 3066 1578 3108
rect 1146 3040 1346 3066
rect 1404 3040 1604 3066
rect 108 2998 308 3024
rect 366 2998 566 3024
rect 128 2956 284 2998
rect 392 2956 548 2998
rect 108 2930 308 2956
rect 366 2930 566 2956
rect -1404 2896 -1204 2922
rect -1146 2896 -946 2922
rect -888 2896 -688 2922
rect -630 2896 -430 2922
rect -2316 2848 -2116 2874
rect -2058 2848 -1858 2874
rect -2288 2806 -2154 2848
rect -2034 2806 -1900 2848
rect -2316 2780 -2116 2806
rect -2058 2780 -1858 2806
rect 1146 2814 1346 2840
rect 1404 2814 1604 2840
rect 1170 2772 1306 2814
rect 1432 2772 1568 2814
rect 1146 2746 1346 2772
rect 1404 2746 1604 2772
rect 108 2704 308 2730
rect 366 2704 566 2730
rect -1404 2670 -1204 2696
rect -1146 2670 -946 2696
rect -888 2670 -688 2696
rect -630 2670 -430 2696
rect -1382 2628 -1246 2670
rect -1104 2628 -968 2670
rect -854 2628 -718 2670
rect -600 2628 -464 2670
rect 132 2662 288 2704
rect 392 2662 548 2704
rect 108 2636 308 2662
rect 366 2636 566 2662
rect -1404 2602 -1204 2628
rect -1146 2602 -946 2628
rect -888 2602 -688 2628
rect -630 2602 -430 2628
rect -2316 2554 -2116 2580
rect -2058 2554 -1858 2580
rect -2270 2512 -2136 2554
rect -2014 2512 -1880 2554
rect -2316 2486 -2116 2512
rect -2058 2486 -1858 2512
rect 1146 2520 1346 2546
rect 1404 2520 1604 2546
rect 1168 2478 1304 2520
rect 1440 2478 1576 2520
rect 1146 2452 1346 2478
rect 1404 2452 1604 2478
rect 108 2410 308 2436
rect 366 2410 566 2436
rect -1404 2378 -1204 2402
rect -1146 2378 -946 2402
rect -888 2378 -688 2402
rect -630 2378 -430 2402
rect -1404 2376 -430 2378
rect -1364 2334 -466 2376
rect 138 2368 294 2410
rect 400 2368 556 2410
rect 108 2342 308 2368
rect 366 2342 566 2368
rect -1404 2308 -1204 2334
rect -1146 2308 -946 2334
rect -888 2308 -688 2334
rect -630 2308 -430 2334
rect -2316 2260 -2116 2286
rect -2058 2260 -1858 2286
rect -2276 2218 -2142 2260
rect -2044 2218 -1910 2260
rect -2316 2192 -2116 2218
rect -2058 2192 -1858 2218
rect 1146 2226 1346 2252
rect 1404 2226 1604 2252
rect 1168 2184 1304 2226
rect 1436 2184 1572 2226
rect 1146 2158 1346 2184
rect 1404 2158 1604 2184
rect 108 2116 308 2142
rect 366 2116 566 2142
rect -1404 2082 -1204 2108
rect -1146 2082 -946 2108
rect -888 2082 -688 2108
rect -630 2082 -430 2108
rect -1384 2040 -1248 2082
rect -1116 2040 -980 2082
rect -848 2040 -712 2082
rect -582 2040 -446 2082
rect 130 2074 286 2116
rect 406 2074 562 2116
rect 108 2048 308 2074
rect 366 2048 566 2074
rect -1404 2014 -1204 2040
rect -1146 2014 -946 2040
rect -888 2014 -688 2040
rect -630 2014 -430 2040
rect -2316 1966 -2116 1992
rect -2058 1966 -1858 1992
rect -2290 1924 -2156 1966
rect -2002 1924 -1868 1966
rect -2316 1898 -2116 1924
rect -2058 1898 -1858 1924
rect 1146 1932 1346 1958
rect 1404 1932 1604 1958
rect 108 1822 308 1848
rect 366 1822 566 1848
rect -1404 1788 -1204 1814
rect -1146 1788 -946 1814
rect -888 1788 -688 1814
rect -630 1788 -430 1814
rect -1366 1746 -1230 1788
rect -1114 1746 -978 1788
rect -854 1746 -718 1788
rect -600 1746 -464 1788
rect -1404 1720 -1204 1746
rect -1146 1720 -946 1746
rect -888 1720 -688 1746
rect -630 1720 -430 1746
rect -2316 1672 -2116 1698
rect -2058 1672 -1858 1698
rect -2302 1630 -2168 1672
rect -2030 1630 -1896 1672
rect -2316 1604 -2116 1630
rect -2058 1604 -1858 1630
rect -268 1586 -200 1590
rect -268 1584 440 1586
rect -268 1550 1092 1584
rect 1822 1566 2222 1590
rect -1404 1494 -1204 1520
rect -1146 1494 -946 1520
rect -888 1494 -688 1520
rect -630 1496 -430 1520
rect -268 1514 1298 1550
rect -268 1496 -200 1514
rect -630 1494 -200 1496
rect -1378 1452 -1242 1494
rect -1126 1452 -990 1494
rect -860 1452 -724 1494
rect -600 1452 -200 1494
rect -1404 1426 -1204 1452
rect -1146 1426 -946 1452
rect -888 1426 -688 1452
rect -630 1426 -430 1452
rect -268 1442 -200 1452
rect 184 1512 1298 1514
rect 184 1450 510 1512
rect 108 1444 566 1450
rect 972 1448 1298 1512
rect 1822 1498 1940 1566
rect 2086 1498 2222 1566
rect -2316 1378 -2116 1404
rect -2058 1378 -1858 1404
rect -2284 1336 -2150 1378
rect -2022 1336 -1888 1378
rect -2316 1310 -2116 1336
rect -2058 1310 -1858 1336
rect 108 1424 308 1444
rect 366 1424 566 1444
rect 896 1442 1354 1448
rect -1404 1200 -1204 1226
rect -1146 1200 -946 1226
rect -888 1200 -688 1226
rect -630 1200 -430 1226
rect 896 1422 1096 1442
rect 1154 1422 1354 1442
rect 1822 1436 2222 1498
rect 1804 1430 2262 1436
rect -1378 1158 -1242 1200
rect -1092 1158 -956 1200
rect -850 1158 -714 1200
rect -604 1158 -468 1200
rect 108 1198 308 1224
rect 366 1198 566 1224
rect 1804 1410 2004 1430
rect 2062 1410 2262 1430
rect -1404 1132 -1204 1158
rect -1146 1132 -946 1158
rect -888 1132 -688 1158
rect -630 1132 -430 1158
rect 128 1156 284 1198
rect 392 1156 548 1198
rect 896 1196 1096 1222
rect 1154 1196 1354 1222
rect -2316 1084 -2116 1110
rect -2058 1084 -1858 1110
rect -2270 1042 -2136 1084
rect -2024 1042 -1890 1084
rect -2316 1016 -2116 1042
rect -2058 1016 -1858 1042
rect 108 1130 308 1156
rect 366 1130 566 1156
rect 916 1154 1072 1196
rect 1180 1154 1336 1196
rect 1804 1184 2004 1210
rect 2062 1184 2262 1210
rect -1404 906 -1204 932
rect -1146 906 -946 932
rect -888 906 -688 932
rect -630 906 -430 932
rect 896 1128 1096 1154
rect 1154 1128 1354 1154
rect 1824 1142 1960 1184
rect 2100 1142 2236 1184
rect -1380 864 -1244 906
rect -1108 864 -972 906
rect -860 864 -724 906
rect -594 864 -458 906
rect 108 904 308 930
rect 366 904 566 930
rect 1804 1116 2004 1142
rect 2062 1116 2262 1142
rect -1404 838 -1204 864
rect -1146 838 -946 864
rect -888 838 -688 864
rect -630 838 -430 864
rect 132 862 288 904
rect 392 862 548 904
rect 896 902 1096 928
rect 1154 902 1354 928
rect -2316 790 -2116 816
rect -2058 790 -1858 816
rect -2286 748 -2152 790
rect -2010 748 -1876 790
rect -2316 722 -2116 748
rect -2058 722 -1858 748
rect 108 836 308 862
rect 366 836 566 862
rect 920 860 1076 902
rect 1180 860 1336 902
rect -1404 612 -1204 638
rect -1146 612 -946 638
rect -888 612 -688 638
rect -630 612 -430 638
rect 896 834 1096 860
rect 1154 834 1354 860
rect -1378 570 -1242 612
rect -1124 570 -988 612
rect -846 570 -710 612
rect -574 570 -438 612
rect 108 610 308 636
rect 366 610 566 636
rect -1404 544 -1204 570
rect -1146 544 -946 570
rect -888 544 -688 570
rect -630 544 -430 570
rect 138 568 294 610
rect 400 568 556 610
rect 896 608 1096 634
rect 1154 608 1354 634
rect -2316 496 -2116 522
rect -2058 496 -1858 522
rect -2298 454 -2164 496
rect -2004 454 -1870 496
rect -2316 428 -2116 454
rect -2058 428 -1858 454
rect 108 542 308 568
rect 366 542 566 568
rect 926 566 1082 608
rect 1188 566 1344 608
rect -1404 318 -1204 344
rect -1146 318 -946 344
rect -888 318 -688 344
rect -630 318 -430 344
rect 896 540 1096 566
rect 1154 540 1354 566
rect -1376 276 -1240 318
rect -1098 276 -962 318
rect -860 276 -724 318
rect -590 276 -454 318
rect 108 316 308 342
rect 366 316 566 342
rect -1404 250 -1204 276
rect -1146 250 -946 276
rect -888 250 -688 276
rect -630 250 -430 276
rect 130 274 286 316
rect 406 274 562 316
rect 896 314 1096 340
rect 1154 314 1354 340
rect -2316 202 -2116 228
rect -2058 202 -1858 228
rect -2294 160 -2160 202
rect -2026 160 -1892 202
rect -2316 134 -2116 160
rect -2058 134 -1858 160
rect 108 248 308 274
rect 366 248 566 274
rect 918 272 1074 314
rect 1194 272 1350 314
rect -1404 24 -1204 50
rect -1146 24 -946 50
rect -888 24 -688 50
rect -630 24 -430 50
rect 896 246 1096 272
rect 1154 246 1354 272
rect 108 22 308 48
rect 366 22 566 48
rect 1804 890 2004 916
rect 2062 890 2262 916
rect 1828 848 1964 890
rect 2090 848 2226 890
rect 1804 822 2004 848
rect 2062 822 2262 848
rect 1804 596 2004 622
rect 2062 596 2262 622
rect 1826 554 1962 596
rect 2098 554 2234 596
rect 1804 528 2004 554
rect 2062 528 2262 554
rect 1804 302 2004 328
rect 2062 302 2262 328
rect 1826 260 1962 302
rect 2094 260 2230 302
rect 1804 234 2004 260
rect 2062 234 2262 260
rect 126 -6 282 22
rect 896 20 1096 46
rect 1154 20 1354 46
rect 1804 8 2004 34
rect 2062 8 2262 34
rect -2316 -92 -2116 -66
rect -2058 -92 -1858 -66
rect 126 -86 160 -6
rect 236 -86 282 -6
rect 126 -122 282 -86
<< polycont >>
rect -2180 4922 -2024 5024
rect 1940 1498 2086 1566
rect 160 -86 236 -6
<< locali >>
rect -2204 5024 -1988 5048
rect -2204 4922 -2180 5024
rect -2024 4922 -1988 5024
rect -2204 4900 -1988 4922
rect -2362 4764 -2328 4780
rect -2362 4696 -2328 4712
rect -2104 4764 -2070 4780
rect -2104 4696 -2070 4712
rect -1846 4764 -1812 4780
rect -1846 4696 -1812 4712
rect -2362 4470 -2328 4486
rect -2362 4402 -2328 4418
rect -2104 4470 -2070 4486
rect -2104 4402 -2070 4418
rect -1846 4470 -1812 4486
rect -1846 4402 -1812 4418
rect -2362 4176 -2328 4192
rect -2362 4108 -2328 4124
rect -2104 4176 -2070 4192
rect -2104 4108 -2070 4124
rect -1846 4176 -1812 4192
rect -1846 4108 -1812 4124
rect -2362 3882 -2328 3898
rect -2362 3814 -2328 3830
rect -2104 3882 -2070 3898
rect -2104 3814 -2070 3830
rect -1846 3882 -1812 3898
rect -1846 3814 -1812 3830
rect -2362 3588 -2328 3604
rect -2362 3520 -2328 3536
rect -2104 3588 -2070 3604
rect -2104 3520 -2070 3536
rect -1846 3588 -1812 3604
rect -1846 3520 -1812 3536
rect -408 3376 -134 3416
rect -2362 3294 -2328 3310
rect -2362 3226 -2328 3242
rect -2104 3294 -2070 3310
rect -2104 3226 -2070 3242
rect -1846 3294 -1812 3310
rect -1846 3226 -1812 3242
rect -408 3054 -378 3376
rect -196 3054 -134 3376
rect 1100 3260 1134 3276
rect 1100 3192 1134 3208
rect 1358 3260 1392 3276
rect 1358 3192 1392 3208
rect 1616 3260 1650 3276
rect 1616 3192 1650 3208
rect 62 3150 96 3166
rect 62 3082 96 3098
rect 320 3150 354 3166
rect 320 3082 354 3098
rect 578 3150 612 3166
rect 578 3082 612 3098
rect -2362 3000 -2328 3016
rect -2362 2932 -2328 2948
rect -2104 3000 -2070 3016
rect -2104 2932 -2070 2948
rect -1846 3000 -1812 3016
rect -408 3000 -134 3054
rect -1846 2932 -1812 2948
rect 1100 2966 1134 2982
rect 1100 2898 1134 2914
rect 1358 2966 1392 2982
rect 1358 2898 1392 2914
rect 1616 2966 1650 2982
rect 1616 2898 1650 2914
rect 62 2856 96 2872
rect -1450 2822 -1416 2838
rect -1450 2754 -1416 2770
rect -1192 2822 -1158 2838
rect -1192 2754 -1158 2770
rect -934 2822 -900 2838
rect -934 2754 -900 2770
rect -676 2822 -642 2838
rect -676 2754 -642 2770
rect -418 2822 -384 2838
rect 62 2788 96 2804
rect 320 2856 354 2872
rect 320 2788 354 2804
rect 578 2856 612 2872
rect 578 2788 612 2804
rect -418 2754 -384 2770
rect -2362 2706 -2328 2722
rect -2584 2594 -2450 2676
rect -2362 2638 -2328 2654
rect -2104 2706 -2070 2722
rect -2104 2638 -2070 2654
rect -1846 2706 -1812 2722
rect -1846 2638 -1812 2654
rect 1100 2672 1134 2688
rect 1100 2604 1134 2620
rect 1358 2672 1392 2688
rect 1358 2604 1392 2620
rect 1616 2672 1650 2688
rect 1616 2604 1650 2620
rect -2584 450 -2560 2594
rect -2482 450 -2450 2594
rect 62 2562 96 2578
rect -1450 2528 -1416 2544
rect -1450 2460 -1416 2476
rect -1192 2528 -1158 2544
rect -1192 2460 -1158 2476
rect -934 2528 -900 2544
rect -934 2460 -900 2476
rect -676 2528 -642 2544
rect -676 2460 -642 2476
rect -418 2528 -384 2544
rect 62 2494 96 2510
rect 320 2562 354 2578
rect 320 2494 354 2510
rect 578 2562 612 2578
rect 578 2494 612 2510
rect -418 2460 -384 2476
rect -2362 2412 -2328 2428
rect -2362 2344 -2328 2360
rect -2104 2412 -2070 2428
rect -2104 2344 -2070 2360
rect -1846 2412 -1812 2428
rect -1846 2344 -1812 2360
rect 1100 2378 1134 2394
rect 1100 2310 1134 2326
rect 1358 2378 1392 2394
rect 1358 2310 1392 2326
rect 1616 2378 1650 2394
rect 1616 2310 1650 2326
rect 62 2268 96 2284
rect -1450 2234 -1416 2250
rect -1450 2166 -1416 2182
rect -1192 2234 -1158 2250
rect -1192 2166 -1158 2182
rect -934 2234 -900 2250
rect -934 2166 -900 2182
rect -676 2234 -642 2250
rect -676 2166 -642 2182
rect -418 2234 -384 2250
rect 62 2200 96 2216
rect 320 2268 354 2284
rect 320 2200 354 2216
rect 578 2268 612 2284
rect 578 2200 612 2216
rect -418 2166 -384 2182
rect -2362 2118 -2328 2134
rect -2362 2050 -2328 2066
rect -2104 2118 -2070 2134
rect -2104 2050 -2070 2066
rect -1846 2118 -1812 2134
rect -1846 2050 -1812 2066
rect 1100 2084 1134 2100
rect 1100 2016 1134 2032
rect 1358 2084 1392 2100
rect 1358 2016 1392 2032
rect 1616 2084 1650 2100
rect 1616 2016 1650 2032
rect 62 1974 96 1990
rect -1450 1940 -1416 1956
rect -1450 1872 -1416 1888
rect -1192 1940 -1158 1956
rect -1192 1872 -1158 1888
rect -934 1940 -900 1956
rect -934 1872 -900 1888
rect -676 1940 -642 1956
rect -676 1872 -642 1888
rect -418 1940 -384 1956
rect 62 1906 96 1922
rect 320 1974 354 1990
rect 320 1906 354 1922
rect 578 1974 612 1990
rect 578 1906 612 1922
rect -418 1872 -384 1888
rect -2362 1824 -2328 1840
rect -2362 1756 -2328 1772
rect -2104 1824 -2070 1840
rect -2104 1756 -2070 1772
rect -1846 1824 -1812 1840
rect -1846 1756 -1812 1772
rect -1450 1646 -1416 1662
rect -1450 1578 -1416 1594
rect -1192 1646 -1158 1662
rect -1192 1578 -1158 1594
rect -934 1646 -900 1662
rect -934 1578 -900 1594
rect -676 1646 -642 1662
rect -676 1578 -642 1594
rect -418 1646 -384 1662
rect -418 1578 -384 1594
rect 1916 1566 2118 1578
rect -2362 1530 -2328 1546
rect -2362 1462 -2328 1478
rect -2104 1530 -2070 1546
rect -2104 1462 -2070 1478
rect -1846 1530 -1812 1546
rect 1916 1498 1940 1566
rect 2086 1498 2118 1566
rect 1916 1478 2118 1498
rect -1846 1462 -1812 1478
rect -1450 1352 -1416 1368
rect -1450 1284 -1416 1300
rect -1192 1352 -1158 1368
rect -1192 1284 -1158 1300
rect -934 1352 -900 1368
rect -934 1284 -900 1300
rect -676 1352 -642 1368
rect -676 1284 -642 1300
rect -418 1352 -384 1368
rect -418 1284 -384 1300
rect 62 1350 96 1366
rect 62 1282 96 1298
rect 320 1350 354 1366
rect 320 1282 354 1298
rect 578 1350 612 1366
rect 578 1282 612 1298
rect 850 1348 884 1364
rect 850 1280 884 1296
rect 1108 1348 1142 1364
rect 1108 1280 1142 1296
rect 1366 1348 1400 1364
rect 1366 1280 1400 1296
rect 1758 1336 1792 1352
rect 1758 1268 1792 1284
rect 2016 1336 2050 1352
rect 2016 1268 2050 1284
rect 2274 1336 2308 1352
rect 2274 1268 2308 1284
rect -2362 1236 -2328 1252
rect -2362 1168 -2328 1184
rect -2104 1236 -2070 1252
rect -2104 1168 -2070 1184
rect -1846 1236 -1812 1252
rect -1846 1168 -1812 1184
rect 2432 1222 2602 1280
rect -1450 1058 -1416 1074
rect -1450 990 -1416 1006
rect -1192 1058 -1158 1074
rect -1192 990 -1158 1006
rect -934 1058 -900 1074
rect -934 990 -900 1006
rect -676 1058 -642 1074
rect -676 990 -642 1006
rect -418 1058 -384 1074
rect -418 990 -384 1006
rect 62 1056 96 1072
rect 62 988 96 1004
rect 320 1056 354 1072
rect 320 988 354 1004
rect 578 1056 612 1072
rect 578 988 612 1004
rect 850 1054 884 1070
rect 850 986 884 1002
rect 1108 1054 1142 1070
rect 1108 986 1142 1002
rect 1366 1054 1400 1070
rect 1366 986 1400 1002
rect 1758 1042 1792 1058
rect 1480 960 1576 994
rect 1758 974 1792 990
rect 2016 1042 2050 1058
rect 2016 974 2050 990
rect 2274 1042 2308 1058
rect 2274 974 2308 990
rect -2362 942 -2328 958
rect -2362 874 -2328 890
rect -2104 942 -2070 958
rect -2104 874 -2070 890
rect -1846 942 -1812 958
rect -1846 874 -1812 890
rect -1450 764 -1416 780
rect -1450 696 -1416 712
rect -1192 764 -1158 780
rect -1192 696 -1158 712
rect -934 764 -900 780
rect -934 696 -900 712
rect -676 764 -642 780
rect -676 696 -642 712
rect -418 764 -384 780
rect -418 696 -384 712
rect 62 762 96 778
rect 62 694 96 710
rect 320 762 354 778
rect 320 694 354 710
rect 578 762 612 778
rect 578 694 612 710
rect 850 760 884 776
rect 850 692 884 708
rect 1108 760 1142 776
rect 1108 692 1142 708
rect 1366 760 1400 776
rect 1366 692 1400 708
rect -2362 648 -2328 664
rect -2362 580 -2328 596
rect -2104 648 -2070 664
rect -2104 580 -2070 596
rect -1846 648 -1812 664
rect -1846 580 -1812 596
rect -2584 328 -2450 450
rect -1450 470 -1416 486
rect -1450 402 -1416 418
rect -1192 470 -1158 486
rect -1192 402 -1158 418
rect -934 470 -900 486
rect -934 402 -900 418
rect -676 470 -642 486
rect -676 402 -642 418
rect -418 470 -384 486
rect -418 402 -384 418
rect 62 468 96 484
rect 62 400 96 416
rect 320 468 354 484
rect 320 400 354 416
rect 578 468 612 484
rect 578 400 612 416
rect 850 466 884 482
rect 850 398 884 414
rect 1108 466 1142 482
rect 1108 398 1142 414
rect 1366 466 1400 482
rect 1366 398 1400 414
rect -2362 354 -2328 370
rect -2362 286 -2328 302
rect -2104 354 -2070 370
rect -2104 286 -2070 302
rect -1846 354 -1812 370
rect -1846 286 -1812 302
rect 1480 238 1492 960
rect 1564 238 1576 960
rect 1758 748 1792 764
rect 1758 680 1792 696
rect 2016 748 2050 764
rect 2016 680 2050 696
rect 2274 748 2308 764
rect 2274 680 2308 696
rect 1758 454 1792 470
rect 1758 386 1792 402
rect 2016 454 2050 470
rect 2016 386 2050 402
rect 2274 454 2308 470
rect 2274 386 2308 402
rect 1480 210 1576 238
rect -1450 176 -1416 192
rect -1450 108 -1416 124
rect -1192 176 -1158 192
rect -1192 108 -1158 124
rect -934 176 -900 192
rect -934 108 -900 124
rect -676 176 -642 192
rect -676 108 -642 124
rect -418 176 -384 192
rect 2432 190 2456 1222
rect 2554 190 2602 1222
rect -418 108 -384 124
rect 62 174 96 190
rect 62 106 96 122
rect 320 174 354 190
rect 320 106 354 122
rect 578 174 612 190
rect 578 106 612 122
rect 850 172 884 188
rect 850 104 884 120
rect 1108 172 1142 188
rect 1108 104 1142 120
rect 1366 172 1400 188
rect 1366 104 1400 120
rect 1758 160 1792 176
rect 1758 92 1792 108
rect 2016 160 2050 176
rect 2016 92 2050 108
rect 2274 160 2308 176
rect 2432 116 2602 190
rect 2274 92 2308 108
rect -2362 60 -2328 76
rect -2362 -8 -2328 8
rect -2104 60 -2070 76
rect -2104 -8 -2070 8
rect -1846 60 -1812 76
rect -1846 -8 -1812 8
rect 144 -6 262 22
rect 144 -86 160 -6
rect 236 -86 262 -6
rect 144 -104 262 -86
<< viali >>
rect -2180 4922 -2024 5024
rect -2362 4712 -2328 4764
rect -2104 4712 -2070 4764
rect -1846 4712 -1812 4764
rect -2362 4418 -2328 4470
rect -2104 4418 -2070 4470
rect -1846 4418 -1812 4470
rect -2362 4124 -2328 4176
rect -2104 4124 -2070 4176
rect -1846 4124 -1812 4176
rect -2362 3830 -2328 3882
rect -2104 3830 -2070 3882
rect -1846 3830 -1812 3882
rect -2362 3536 -2328 3588
rect -2104 3536 -2070 3588
rect -1846 3536 -1812 3588
rect -2362 3242 -2328 3294
rect -2104 3242 -2070 3294
rect -1846 3242 -1812 3294
rect -378 3054 -196 3376
rect 1100 3208 1134 3260
rect 1358 3208 1392 3260
rect 1616 3208 1650 3260
rect 62 3098 96 3150
rect 320 3098 354 3150
rect 578 3098 612 3150
rect -2362 2948 -2328 3000
rect -2104 2948 -2070 3000
rect -1846 2948 -1812 3000
rect 1100 2914 1134 2966
rect 1358 2914 1392 2966
rect 1616 2914 1650 2966
rect -1450 2770 -1416 2822
rect -1192 2770 -1158 2822
rect -934 2770 -900 2822
rect -676 2770 -642 2822
rect -418 2770 -384 2822
rect 62 2804 96 2856
rect 320 2804 354 2856
rect 578 2804 612 2856
rect -2362 2654 -2328 2706
rect -2104 2654 -2070 2706
rect -1846 2654 -1812 2706
rect 1100 2620 1134 2672
rect 1358 2620 1392 2672
rect 1616 2620 1650 2672
rect -2554 528 -2486 2562
rect -1450 2476 -1416 2528
rect -1192 2476 -1158 2528
rect -934 2476 -900 2528
rect -676 2476 -642 2528
rect -418 2476 -384 2528
rect 62 2510 96 2562
rect 320 2510 354 2562
rect 578 2510 612 2562
rect -2362 2360 -2328 2412
rect -2104 2360 -2070 2412
rect -1846 2360 -1812 2412
rect 1100 2326 1134 2378
rect 1358 2326 1392 2378
rect 1616 2326 1650 2378
rect -1450 2182 -1416 2234
rect -1192 2182 -1158 2234
rect -934 2182 -900 2234
rect -676 2182 -642 2234
rect -418 2182 -384 2234
rect 62 2216 96 2268
rect 320 2216 354 2268
rect 578 2216 612 2268
rect -2362 2066 -2328 2118
rect -2104 2066 -2070 2118
rect -1846 2066 -1812 2118
rect 1100 2032 1134 2084
rect 1358 2032 1392 2084
rect 1616 2032 1650 2084
rect -1450 1888 -1416 1940
rect -1192 1888 -1158 1940
rect -934 1888 -900 1940
rect -676 1888 -642 1940
rect -418 1888 -384 1940
rect 62 1922 96 1974
rect 320 1922 354 1974
rect 578 1922 612 1974
rect -2362 1772 -2328 1824
rect -2104 1772 -2070 1824
rect -1846 1772 -1812 1824
rect -1450 1594 -1416 1646
rect -1192 1594 -1158 1646
rect -934 1594 -900 1646
rect -676 1594 -642 1646
rect -418 1594 -384 1646
rect -2362 1478 -2328 1530
rect -2104 1478 -2070 1530
rect -1846 1478 -1812 1530
rect 1960 1506 2062 1558
rect -1450 1300 -1416 1352
rect -1192 1300 -1158 1352
rect -934 1300 -900 1352
rect -676 1300 -642 1352
rect -418 1300 -384 1352
rect 62 1298 96 1350
rect 320 1298 354 1350
rect 578 1298 612 1350
rect 850 1296 884 1348
rect 1108 1296 1142 1348
rect 1366 1296 1400 1348
rect 1758 1284 1792 1336
rect 2016 1284 2050 1336
rect 2274 1284 2308 1336
rect -2362 1184 -2328 1236
rect -2104 1184 -2070 1236
rect -1846 1184 -1812 1236
rect -1450 1006 -1416 1058
rect -1192 1006 -1158 1058
rect -934 1006 -900 1058
rect -676 1006 -642 1058
rect -418 1006 -384 1058
rect 62 1004 96 1056
rect 320 1004 354 1056
rect 578 1004 612 1056
rect 850 1002 884 1054
rect 1108 1002 1142 1054
rect 1366 1002 1400 1054
rect 1758 990 1792 1042
rect 2016 990 2050 1042
rect 2274 990 2308 1042
rect -2362 890 -2328 942
rect -2104 890 -2070 942
rect -1846 890 -1812 942
rect -1450 712 -1416 764
rect -1192 712 -1158 764
rect -934 712 -900 764
rect -676 712 -642 764
rect -418 712 -384 764
rect 62 710 96 762
rect 320 710 354 762
rect 578 710 612 762
rect 850 708 884 760
rect 1108 708 1142 760
rect 1366 708 1400 760
rect -2362 596 -2328 648
rect -2104 596 -2070 648
rect -1846 596 -1812 648
rect -1450 418 -1416 470
rect -1192 418 -1158 470
rect -934 418 -900 470
rect -676 418 -642 470
rect -418 418 -384 470
rect 62 416 96 468
rect 320 416 354 468
rect 578 416 612 468
rect 850 414 884 466
rect 1108 414 1142 466
rect 1366 414 1400 466
rect -2362 302 -2328 354
rect -2104 302 -2070 354
rect -1846 302 -1812 354
rect 1498 268 1552 922
rect 1758 696 1792 748
rect 2016 696 2050 748
rect 2274 696 2308 748
rect 1758 402 1792 454
rect 2016 402 2050 454
rect 2274 402 2308 454
rect -1450 124 -1416 176
rect -1192 124 -1158 176
rect -934 124 -900 176
rect -676 124 -642 176
rect 2456 190 2554 1222
rect -418 124 -384 176
rect 62 122 96 174
rect 320 122 354 174
rect 578 122 612 174
rect 850 120 884 172
rect 1108 120 1142 172
rect 1366 120 1400 172
rect 1758 108 1792 160
rect 2016 108 2050 160
rect 2274 108 2308 160
rect -2362 8 -2328 60
rect -2104 8 -2070 60
rect -1846 8 -1812 60
rect 160 -86 236 -6
<< metal1 >>
rect -2204 5024 -1988 5048
rect -1770 5024 -1760 5082
rect -2204 4922 -2180 5024
rect -2024 4958 -1760 5024
rect -2024 4922 -1988 4958
rect -1770 4928 -1760 4958
rect -1590 4928 -1580 5082
rect -2204 4900 -1988 4922
rect -2374 4830 -1792 4844
rect -2642 4686 -2632 4810
rect -2528 4780 -2518 4810
rect -2376 4808 -1792 4830
rect -2376 4780 -2326 4808
rect -2528 4776 -2326 4780
rect -1858 4776 -1812 4808
rect -2528 4764 -2322 4776
rect -2528 4712 -2362 4764
rect -2328 4740 -2322 4764
rect -2110 4764 -2064 4776
rect -2328 4712 -2320 4740
rect -2528 4702 -2320 4712
rect -2528 4686 -2518 4702
rect -2370 4470 -2320 4702
rect -2110 4712 -2104 4764
rect -2070 4756 -2064 4764
rect -1858 4764 -1806 4776
rect -2070 4712 -2056 4756
rect -1858 4734 -1846 4764
rect -2110 4700 -2056 4712
rect -2106 4482 -2056 4700
rect -2370 4418 -2362 4470
rect -2328 4418 -2320 4470
rect -2370 4176 -2320 4418
rect -2110 4470 -2056 4482
rect -2110 4418 -2104 4470
rect -2070 4418 -2056 4470
rect -2110 4406 -2056 4418
rect -2106 4188 -2056 4406
rect -2370 4124 -2362 4176
rect -2328 4124 -2320 4176
rect -2370 3882 -2320 4124
rect -2110 4176 -2056 4188
rect -2110 4124 -2104 4176
rect -2070 4124 -2056 4176
rect -2110 4112 -2056 4124
rect -2106 3894 -2056 4112
rect -2370 3830 -2362 3882
rect -2328 3830 -2320 3882
rect -2370 3588 -2320 3830
rect -2110 3882 -2056 3894
rect -2110 3830 -2104 3882
rect -2070 3830 -2056 3882
rect -2110 3818 -2056 3830
rect -2106 3600 -2056 3818
rect -2370 3536 -2362 3588
rect -2328 3536 -2320 3588
rect -2370 3294 -2320 3536
rect -2110 3588 -2056 3600
rect -2110 3536 -2104 3588
rect -2070 3536 -2056 3588
rect -2110 3524 -2056 3536
rect -2106 3306 -2056 3524
rect -2370 3242 -2362 3294
rect -2328 3242 -2320 3294
rect -2370 3000 -2320 3242
rect -2110 3294 -2056 3306
rect -2110 3242 -2104 3294
rect -2070 3242 -2056 3294
rect -2110 3230 -2056 3242
rect -2106 3012 -2056 3230
rect -2370 2948 -2362 3000
rect -2328 2948 -2320 3000
rect -2370 2706 -2320 2948
rect -2110 3000 -2056 3012
rect -2110 2948 -2104 3000
rect -2070 2948 -2056 3000
rect -2110 2936 -2056 2948
rect -2106 2718 -2056 2936
rect -2584 2562 -2450 2676
rect -2584 528 -2554 2562
rect -2486 528 -2450 2562
rect -2584 328 -2450 528
rect -2370 2654 -2362 2706
rect -2328 2654 -2320 2706
rect -2370 2412 -2320 2654
rect -2110 2706 -2056 2718
rect -2110 2654 -2104 2706
rect -2070 2654 -2056 2706
rect -2110 2642 -2056 2654
rect -2106 2424 -2056 2642
rect -2370 2360 -2362 2412
rect -2328 2360 -2320 2412
rect -2370 2118 -2320 2360
rect -2110 2412 -2056 2424
rect -2110 2360 -2104 2412
rect -2070 2360 -2056 2412
rect -2110 2348 -2056 2360
rect -2106 2130 -2056 2348
rect -2370 2066 -2362 2118
rect -2328 2066 -2320 2118
rect -2370 1824 -2320 2066
rect -2110 2118 -2056 2130
rect -2110 2066 -2104 2118
rect -2070 2066 -2056 2118
rect -2110 2054 -2056 2066
rect -2106 1836 -2056 2054
rect -2370 1772 -2362 1824
rect -2328 1772 -2320 1824
rect -2370 1530 -2320 1772
rect -2110 1824 -2056 1836
rect -2110 1772 -2104 1824
rect -2070 1772 -2056 1824
rect -2110 1760 -2056 1772
rect -2106 1542 -2056 1760
rect -2370 1478 -2362 1530
rect -2328 1478 -2320 1530
rect -2370 1236 -2320 1478
rect -2110 1530 -2056 1542
rect -2110 1478 -2104 1530
rect -2070 1478 -2056 1530
rect -2110 1466 -2056 1478
rect -2106 1248 -2056 1466
rect -2370 1184 -2362 1236
rect -2328 1184 -2320 1236
rect -2370 942 -2320 1184
rect -2110 1236 -2056 1248
rect -2110 1184 -2104 1236
rect -2070 1184 -2056 1236
rect -2110 1172 -2056 1184
rect -2106 954 -2056 1172
rect -2370 890 -2362 942
rect -2328 890 -2320 942
rect -2370 648 -2320 890
rect -2110 942 -2056 954
rect -2110 890 -2104 942
rect -2070 890 -2056 942
rect -2110 878 -2056 890
rect -2106 660 -2056 878
rect -2370 596 -2362 648
rect -2328 596 -2320 648
rect -2370 354 -2320 596
rect -2110 648 -2056 660
rect -2110 596 -2104 648
rect -2070 596 -2056 648
rect -2110 584 -2056 596
rect -2106 366 -2056 584
rect -2558 -214 -2490 328
rect -2370 302 -2362 354
rect -2328 302 -2320 354
rect -2370 60 -2320 302
rect -2110 354 -2056 366
rect -2110 302 -2104 354
rect -2070 302 -2056 354
rect -2110 290 -2056 302
rect -2106 72 -2056 290
rect -2370 18 -2362 60
rect -2368 8 -2362 18
rect -2328 18 -2320 60
rect -2110 60 -2056 72
rect -2110 58 -2104 60
rect -2328 8 -2322 18
rect -2368 -4 -2322 8
rect -2112 8 -2104 58
rect -2070 34 -2056 60
rect -1856 4712 -1846 4734
rect -1812 4712 -1806 4764
rect -1514 4750 2742 5148
rect -1856 4470 -1806 4712
rect -1856 4418 -1846 4470
rect -1812 4418 -1806 4470
rect -1856 4176 -1806 4418
rect -1856 4124 -1846 4176
rect -1812 4124 -1806 4176
rect -1856 3882 -1806 4124
rect -1856 3830 -1846 3882
rect -1812 3830 -1806 3882
rect -1856 3588 -1806 3830
rect -1856 3536 -1846 3588
rect -1812 3536 -1806 3588
rect -1856 3294 -1806 3536
rect -1856 3242 -1846 3294
rect -1812 3242 -1806 3294
rect -1856 3000 -1806 3242
rect -1856 2948 -1846 3000
rect -1812 2948 -1806 3000
rect -1856 2706 -1806 2948
rect -1430 4738 2742 4750
rect -1430 2918 -1258 4738
rect -328 3416 -250 4738
rect 42 4732 88 4738
rect 956 4732 1004 4738
rect 1048 3814 1058 3954
rect 1208 3814 1218 3954
rect -408 3376 -134 3416
rect -408 3054 -378 3376
rect -196 3054 -134 3376
rect 1092 3342 1146 3814
rect 1608 3342 1656 3344
rect 1072 3304 1674 3342
rect 1082 3260 1146 3304
rect 46 3224 610 3230
rect 46 3220 618 3224
rect 28 3192 618 3220
rect 1082 3208 1100 3260
rect 1134 3220 1146 3260
rect 1352 3260 1398 3272
rect 1352 3226 1358 3260
rect 1134 3208 1140 3220
rect 1082 3192 1140 3208
rect 28 3162 98 3192
rect 28 3150 102 3162
rect 28 3114 62 3150
rect 50 3110 62 3114
rect -408 3000 -134 3054
rect 52 3098 62 3110
rect 96 3134 102 3150
rect 314 3150 360 3162
rect 96 3098 106 3134
rect -952 2918 -894 2920
rect -1460 2906 -378 2918
rect -1460 2872 -366 2906
rect -1460 2822 -1402 2872
rect -1460 2808 -1450 2822
rect -1856 2654 -1846 2706
rect -1812 2654 -1806 2706
rect -1856 2412 -1806 2654
rect -1856 2360 -1846 2412
rect -1812 2360 -1806 2412
rect -1856 2118 -1806 2360
rect -1856 2066 -1846 2118
rect -1812 2066 -1806 2118
rect -1856 1824 -1806 2066
rect -1856 1772 -1846 1824
rect -1812 1772 -1806 1824
rect -1856 1530 -1806 1772
rect -1856 1478 -1846 1530
rect -1812 1478 -1806 1530
rect -1856 1236 -1806 1478
rect -1856 1184 -1846 1236
rect -1812 1184 -1806 1236
rect -1856 942 -1806 1184
rect -1856 890 -1846 942
rect -1812 890 -1806 942
rect -1856 648 -1806 890
rect -1856 596 -1846 648
rect -1812 596 -1806 648
rect -1856 354 -1806 596
rect -1856 302 -1846 354
rect -1812 302 -1806 354
rect -1856 60 -1806 302
rect -1464 2770 -1450 2808
rect -1416 2800 -1402 2822
rect -1198 2822 -1152 2834
rect -1198 2812 -1192 2822
rect -1416 2770 -1408 2800
rect -1464 2528 -1408 2770
rect -1464 2476 -1450 2528
rect -1416 2476 -1408 2528
rect -1464 2234 -1408 2476
rect -1464 2182 -1450 2234
rect -1416 2182 -1408 2234
rect -1464 1940 -1408 2182
rect -1464 1888 -1450 1940
rect -1416 1888 -1408 1940
rect -1464 1646 -1408 1888
rect -1464 1594 -1450 1646
rect -1416 1594 -1408 1646
rect -1464 1352 -1408 1594
rect -1464 1300 -1450 1352
rect -1416 1300 -1408 1352
rect -1464 1058 -1408 1300
rect -1464 1006 -1450 1058
rect -1416 1006 -1408 1058
rect -1464 764 -1408 1006
rect -1464 712 -1450 764
rect -1416 712 -1408 764
rect -1464 470 -1408 712
rect -1464 418 -1450 470
rect -1416 418 -1408 470
rect -1464 176 -1408 418
rect -1200 2770 -1192 2812
rect -1158 2812 -1152 2822
rect -952 2822 -894 2872
rect -1158 2770 -1144 2812
rect -952 2802 -934 2822
rect -1200 2528 -1144 2770
rect -1200 2476 -1192 2528
rect -1158 2476 -1144 2528
rect -1200 2234 -1144 2476
rect -1200 2182 -1192 2234
rect -1158 2182 -1144 2234
rect -1200 1940 -1144 2182
rect -1200 1888 -1192 1940
rect -1158 1888 -1144 1940
rect -1200 1646 -1144 1888
rect -1200 1594 -1192 1646
rect -1158 1594 -1144 1646
rect -1200 1352 -1144 1594
rect -1200 1300 -1192 1352
rect -1158 1300 -1144 1352
rect -1200 1058 -1144 1300
rect -1200 1006 -1192 1058
rect -1158 1006 -1144 1058
rect -1200 764 -1144 1006
rect -1200 712 -1192 764
rect -1158 712 -1144 764
rect -1200 470 -1144 712
rect -1200 418 -1192 470
rect -1158 418 -1144 470
rect -1200 190 -1144 418
rect -1464 144 -1450 176
rect -1456 124 -1450 144
rect -1416 144 -1408 176
rect -1210 176 -1144 190
rect -1416 124 -1410 144
rect -1456 112 -1410 124
rect -1210 124 -1192 176
rect -1158 124 -1144 176
rect -944 2770 -934 2802
rect -900 2808 -894 2822
rect -682 2822 -636 2834
rect -682 2810 -676 2822
rect -900 2770 -888 2808
rect -944 2528 -888 2770
rect -688 2770 -676 2810
rect -642 2810 -636 2822
rect -424 2822 -366 2872
rect 52 2866 106 3098
rect -642 2770 -632 2810
rect -688 2632 -632 2770
rect -424 2770 -418 2822
rect -384 2788 -366 2822
rect 36 2856 106 2866
rect 36 2804 62 2856
rect 96 2804 106 2856
rect -384 2770 -368 2788
rect 36 2774 106 2804
rect -944 2476 -934 2528
rect -900 2476 -888 2528
rect -944 2234 -888 2476
rect -718 2434 -708 2632
rect -606 2434 -596 2632
rect -424 2528 -368 2770
rect 52 2660 106 2774
rect 314 3098 320 3150
rect 354 3118 360 3150
rect 570 3150 618 3192
rect 354 3098 368 3118
rect 570 3110 578 3150
rect 314 2856 368 3098
rect 572 3098 578 3110
rect 612 3142 618 3150
rect 612 3098 628 3142
rect 572 3086 628 3098
rect 574 2868 628 3086
rect 314 2804 320 2856
rect 354 2804 368 2856
rect -424 2476 -418 2528
rect -384 2476 -368 2528
rect -944 2182 -934 2234
rect -900 2182 -888 2234
rect -944 1940 -888 2182
rect -944 1888 -934 1940
rect -900 1888 -888 1940
rect -944 1646 -888 1888
rect -944 1594 -934 1646
rect -900 1594 -888 1646
rect -944 1352 -888 1594
rect -944 1300 -934 1352
rect -900 1300 -888 1352
rect -944 1058 -888 1300
rect -944 1006 -934 1058
rect -900 1006 -888 1058
rect -944 764 -888 1006
rect -944 712 -934 764
rect -900 712 -888 764
rect -944 470 -888 712
rect -944 418 -934 470
rect -900 418 -888 470
rect -944 176 -888 418
rect -688 2234 -632 2434
rect -688 2182 -676 2234
rect -642 2182 -632 2234
rect -688 1940 -632 2182
rect -688 1888 -676 1940
rect -642 1888 -632 1940
rect -688 1646 -632 1888
rect -688 1594 -676 1646
rect -642 1594 -632 1646
rect -688 1352 -632 1594
rect -688 1300 -676 1352
rect -642 1300 -632 1352
rect -688 1058 -632 1300
rect -688 1006 -676 1058
rect -642 1006 -632 1058
rect -688 764 -632 1006
rect -688 712 -676 764
rect -642 712 -632 764
rect -688 470 -632 712
rect -688 418 -676 470
rect -642 418 -632 470
rect -688 184 -632 418
rect -424 2234 -368 2476
rect -30 2466 -20 2660
rect 148 2466 158 2660
rect 314 2562 368 2804
rect 572 2856 628 2868
rect 572 2804 578 2856
rect 612 2804 628 2856
rect 572 2792 628 2804
rect 574 2574 628 2792
rect 314 2510 320 2562
rect 354 2510 368 2562
rect -424 2182 -418 2234
rect -384 2182 -368 2234
rect -424 1940 -368 2182
rect 52 2268 106 2466
rect 52 2216 62 2268
rect 96 2216 106 2268
rect 52 1974 106 2216
rect 314 2268 368 2510
rect 572 2562 628 2574
rect 572 2510 578 2562
rect 612 2510 628 2562
rect 572 2498 628 2510
rect 574 2280 628 2498
rect 314 2216 320 2268
rect 354 2216 368 2268
rect 314 1974 368 2216
rect 572 2268 628 2280
rect 572 2216 578 2268
rect 612 2216 628 2268
rect 572 2204 628 2216
rect 574 1986 628 2204
rect 1090 2966 1140 3192
rect 1090 2914 1100 2966
rect 1134 2914 1140 2966
rect 1090 2672 1140 2914
rect 1090 2620 1100 2672
rect 1134 2620 1140 2672
rect 1090 2378 1140 2620
rect 1090 2326 1100 2378
rect 1134 2326 1140 2378
rect 1090 2084 1140 2326
rect 1090 2046 1100 2084
rect 1094 2032 1100 2046
rect 1134 2032 1140 2084
rect 1350 3208 1358 3226
rect 1392 3226 1398 3260
rect 1608 3260 1656 3304
rect 1392 3208 1400 3226
rect 1350 2966 1400 3208
rect 1608 3208 1616 3260
rect 1650 3228 1656 3260
rect 1650 3208 1662 3228
rect 1608 3202 1662 3208
rect 1610 3196 1662 3202
rect 1612 3148 1662 3196
rect 1612 3086 1708 3148
rect 1612 2978 1662 3086
rect 1350 2914 1358 2966
rect 1392 2914 1400 2966
rect 1350 2672 1400 2914
rect 1610 2966 1662 2978
rect 1610 2914 1616 2966
rect 1650 2914 1662 2966
rect 1610 2902 1662 2914
rect 1612 2684 1662 2902
rect 1350 2620 1358 2672
rect 1392 2620 1400 2672
rect 1350 2378 1400 2620
rect 1610 2672 1662 2684
rect 1610 2620 1616 2672
rect 1650 2620 1662 2672
rect 1610 2608 1662 2620
rect 1612 2390 1662 2608
rect 1350 2326 1358 2378
rect 1392 2326 1400 2378
rect 1350 2084 1400 2326
rect 1610 2378 1662 2390
rect 1610 2326 1616 2378
rect 1650 2326 1662 2378
rect 1610 2314 1662 2326
rect 1612 2096 1662 2314
rect 1350 2048 1358 2084
rect 1094 2020 1140 2032
rect 1352 2032 1358 2048
rect 1392 2048 1400 2084
rect 1610 2084 1662 2096
rect 1392 2032 1398 2048
rect 1352 2020 1398 2032
rect 1610 2032 1616 2084
rect 1650 2050 1662 2084
rect 1650 2032 1656 2050
rect 1610 2020 1656 2032
rect 52 1942 62 1974
rect -424 1888 -418 1940
rect -384 1888 -368 1940
rect 56 1922 62 1942
rect 96 1942 106 1974
rect 96 1922 102 1942
rect 56 1910 102 1922
rect 312 1922 320 1974
rect 354 1948 368 1974
rect 572 1974 628 1986
rect 354 1922 366 1948
rect -424 1646 -368 1888
rect 312 1846 366 1922
rect 572 1922 578 1974
rect 612 1950 628 1974
rect 612 1922 618 1950
rect 572 1910 618 1922
rect 1352 1944 1394 2020
rect 1352 1878 2466 1944
rect 1494 1846 1550 1878
rect 312 1792 1558 1846
rect 1494 1784 1550 1792
rect -424 1594 -418 1646
rect -384 1594 -368 1646
rect -424 1352 -368 1594
rect 1676 1486 1686 1600
rect 1758 1550 1768 1600
rect 1916 1558 2118 1578
rect 1916 1550 1960 1558
rect 1758 1506 1960 1550
rect 2062 1506 2118 1558
rect 1758 1504 2118 1506
rect 1758 1486 1768 1504
rect 1916 1478 2118 1504
rect 46 1424 610 1430
rect 834 1424 1398 1428
rect 46 1422 1398 1424
rect 1494 1422 1560 1452
rect 46 1392 1560 1422
rect 2012 1418 2042 1478
rect 2266 1418 2314 1420
rect -424 1300 -418 1352
rect -384 1300 -368 1352
rect 50 1362 98 1392
rect 554 1390 1560 1392
rect 554 1382 908 1390
rect 570 1378 908 1382
rect 50 1350 102 1362
rect 50 1310 62 1350
rect -424 1216 -368 1300
rect 52 1298 62 1310
rect 96 1334 102 1350
rect 314 1350 360 1362
rect 96 1298 106 1334
rect 52 1216 106 1298
rect -424 1176 106 1216
rect -424 1058 -368 1176
rect -424 1006 -418 1058
rect -384 1006 -368 1058
rect -424 764 -368 1006
rect -424 712 -418 764
rect -384 712 -368 764
rect -424 470 -368 712
rect -424 418 -418 470
rect -384 418 -368 470
rect -944 144 -934 176
rect -2070 8 -2064 34
rect -1856 32 -1846 60
rect -2112 -4 -2064 8
rect -1852 8 -1846 32
rect -1812 8 -1806 60
rect -1210 72 -1144 124
rect -940 124 -934 144
rect -900 144 -888 176
rect -696 176 -630 184
rect -900 124 -894 144
rect -940 112 -894 124
rect -696 124 -676 176
rect -642 124 -630 176
rect -696 72 -630 124
rect -424 176 -368 418
rect -424 124 -418 176
rect -384 154 -368 176
rect 52 1056 106 1176
rect 52 1004 62 1056
rect 96 1004 106 1056
rect 52 762 106 1004
rect 52 710 62 762
rect 96 710 106 762
rect 52 468 106 710
rect 52 416 62 468
rect 96 416 106 468
rect 52 174 106 416
rect 314 1298 320 1350
rect 354 1318 360 1350
rect 570 1350 618 1378
rect 354 1298 368 1318
rect 570 1310 578 1350
rect 314 1056 368 1298
rect 572 1298 578 1310
rect 612 1342 618 1350
rect 838 1348 908 1378
rect 612 1298 628 1342
rect 838 1308 850 1348
rect 572 1286 628 1298
rect 574 1068 628 1286
rect 314 1004 320 1056
rect 354 1004 368 1056
rect 314 762 368 1004
rect 572 1056 628 1068
rect 572 1004 578 1056
rect 612 1004 628 1056
rect 572 992 628 1004
rect 574 774 628 992
rect 314 710 320 762
rect 354 710 368 762
rect 314 468 368 710
rect 572 762 628 774
rect 572 710 578 762
rect 612 710 628 762
rect 572 698 628 710
rect 574 480 628 698
rect 314 416 320 468
rect 354 416 368 468
rect 314 178 368 416
rect 572 468 628 480
rect 572 416 578 468
rect 612 416 628 468
rect 572 404 628 416
rect 574 186 628 404
rect -384 124 -378 154
rect 52 142 62 174
rect -424 112 -378 124
rect 56 122 62 142
rect 96 142 106 174
rect 308 174 378 178
rect 96 122 102 142
rect 56 110 102 122
rect 308 122 320 174
rect 354 122 378 174
rect -1210 28 -622 72
rect -696 22 -630 28
rect -1852 -4 -1806 8
rect 144 -2 262 22
rect 308 -2 378 122
rect 572 174 628 186
rect 572 122 578 174
rect 612 150 628 174
rect 840 1296 850 1308
rect 884 1324 908 1348
rect 1102 1348 1148 1360
rect 884 1296 894 1324
rect 840 1054 894 1296
rect 840 1002 850 1054
rect 884 1002 894 1054
rect 840 760 894 1002
rect 840 708 850 760
rect 884 708 894 760
rect 840 466 894 708
rect 840 414 850 466
rect 884 414 894 466
rect 840 172 894 414
rect 1102 1296 1108 1348
rect 1142 1316 1148 1348
rect 1358 1348 1406 1390
rect 1466 1360 1560 1390
rect 1730 1380 2332 1418
rect 1142 1296 1156 1316
rect 1358 1308 1366 1348
rect 1102 1054 1156 1296
rect 1360 1296 1366 1308
rect 1400 1340 1406 1348
rect 1400 1296 1416 1340
rect 1360 1284 1416 1296
rect 1362 1066 1416 1284
rect 1102 1002 1108 1054
rect 1142 1002 1156 1054
rect 1102 760 1156 1002
rect 1360 1054 1416 1066
rect 1360 1002 1366 1054
rect 1400 1002 1416 1054
rect 1360 990 1416 1002
rect 1494 994 1560 1360
rect 1740 1336 1802 1380
rect 1740 1284 1758 1336
rect 1792 1302 1802 1336
rect 2010 1336 2056 1348
rect 2010 1302 2016 1336
rect 1792 1284 1798 1302
rect 1740 1268 1798 1284
rect 1748 1042 1798 1268
rect 1362 772 1416 990
rect 1102 708 1108 760
rect 1142 708 1156 760
rect 1102 466 1156 708
rect 1360 760 1416 772
rect 1360 708 1366 760
rect 1400 708 1416 760
rect 1360 696 1416 708
rect 1362 478 1416 696
rect 1102 414 1108 466
rect 1142 414 1156 466
rect 1102 212 1156 414
rect 1360 466 1416 478
rect 1360 414 1366 466
rect 1400 414 1416 466
rect 1360 402 1416 414
rect 612 122 618 150
rect 840 140 850 172
rect 572 110 618 122
rect 844 120 850 140
rect 884 140 894 172
rect 1080 172 1182 212
rect 1362 184 1416 402
rect 1480 922 1576 994
rect 1480 268 1498 922
rect 1552 268 1576 922
rect 1480 210 1576 268
rect 1748 990 1758 1042
rect 1792 990 1798 1042
rect 1748 748 1798 990
rect 1748 696 1758 748
rect 1792 696 1798 748
rect 1748 454 1798 696
rect 1748 402 1758 454
rect 1792 402 1798 454
rect 884 120 890 140
rect 844 108 890 120
rect 1080 120 1108 172
rect 1142 120 1182 172
rect -2112 -214 -2068 -4
rect 144 -6 378 -2
rect 144 -86 160 -6
rect 236 -24 378 -6
rect 1080 60 1182 120
rect 1360 172 1416 184
rect 1360 120 1366 172
rect 1400 148 1416 172
rect 1748 166 1798 402
rect 2008 1284 2016 1302
rect 2050 1302 2056 1336
rect 2266 1336 2314 1380
rect 2050 1284 2058 1302
rect 2008 1042 2058 1284
rect 2266 1284 2274 1336
rect 2308 1304 2314 1336
rect 2308 1284 2320 1304
rect 2266 1278 2320 1284
rect 2268 1272 2320 1278
rect 2270 1054 2320 1272
rect 2008 990 2016 1042
rect 2050 990 2058 1042
rect 2008 748 2058 990
rect 2268 1042 2320 1054
rect 2268 990 2274 1042
rect 2308 990 2320 1042
rect 2268 978 2320 990
rect 2270 760 2320 978
rect 2008 696 2016 748
rect 2050 696 2058 748
rect 2008 454 2058 696
rect 2268 748 2320 760
rect 2268 696 2274 748
rect 2308 696 2320 748
rect 2268 684 2320 696
rect 2270 466 2320 684
rect 2008 402 2016 454
rect 2050 402 2058 454
rect 2008 178 2058 402
rect 2268 454 2320 466
rect 2432 1222 2602 1280
rect 2432 464 2456 1222
rect 2268 402 2274 454
rect 2308 402 2320 454
rect 2268 390 2320 402
rect 1720 160 1810 166
rect 1400 120 1406 148
rect 1360 108 1406 120
rect 1720 108 1758 160
rect 1792 108 1810 160
rect 1720 60 1810 108
rect 1080 -16 1810 60
rect 1720 -18 1810 -16
rect 2000 160 2058 178
rect 2270 172 2320 390
rect 2000 108 2016 160
rect 2050 124 2058 160
rect 2268 160 2320 172
rect 2050 108 2056 124
rect 2000 96 2056 108
rect 2268 108 2274 160
rect 2308 126 2320 160
rect 2426 190 2456 464
rect 2554 190 2602 1222
rect 2308 108 2314 126
rect 2268 96 2314 108
rect 2426 116 2602 190
rect 236 -50 366 -24
rect 236 -86 262 -50
rect 144 -104 262 -86
rect 2000 -214 2052 96
rect 2426 -214 2588 116
rect -2558 -630 2676 -214
<< via1 >>
rect -1760 4928 -1590 5082
rect -2632 4686 -2528 4810
rect 1058 3814 1208 3954
rect -708 2528 -606 2632
rect -708 2476 -676 2528
rect -676 2476 -642 2528
rect -642 2476 -606 2528
rect -708 2434 -606 2476
rect -20 2562 148 2660
rect -20 2510 62 2562
rect 62 2510 96 2562
rect 96 2510 148 2562
rect -20 2466 148 2510
rect 1686 1486 1758 1600
<< metal2 >>
rect -1760 5082 -1590 5092
rect -1760 4918 -1590 4928
rect -2632 4810 -2528 4820
rect -2632 4676 -2528 4686
rect -1668 1558 -1596 4918
rect 1058 3954 1208 3964
rect 1058 3804 1208 3814
rect -20 2660 148 2670
rect -708 2632 -606 2642
rect -606 2516 -20 2562
rect -20 2456 148 2466
rect -708 2424 -606 2434
rect 1686 1600 1758 1610
rect -1670 1498 1686 1558
rect -1668 1480 -1596 1498
rect 1686 1476 1758 1486
<< via2 >>
rect -2632 4686 -2528 4810
rect 1058 3814 1208 3954
<< metal3 >>
rect -2642 4810 -2518 4815
rect -2642 4686 -2632 4810
rect -2528 4686 -2518 4810
rect -2642 4681 -2518 4686
rect -2588 4598 -2528 4681
rect 114 4598 912 4600
rect 1084 4598 1158 4602
rect -2590 4530 1158 4598
rect 114 4528 912 4530
rect 1084 3959 1158 4530
rect 1048 3954 1218 3959
rect 1048 3814 1058 3954
rect 1208 3814 1218 3954
rect 1048 3809 1218 3814
<< labels >>
flabel metal1 -612 4962 -612 4962 0 FreeSans 1600 0 0 0 vdda
flabel metal1 332 4 332 4 0 FreeSans 1600 0 0 0 Iin
flabel metal1 2208 1902 2208 1904 0 FreeSans 1600 0 0 0 vc
flabel poly 1326 3494 1326 3494 0 FreeSans 1600 0 0 0 out2
flabel poly 282 3362 282 3362 0 FreeSans 1600 0 0 0 out1
flabel metal3 448 4556 448 4556 0 FreeSans 1600 0 0 0 nc
flabel metal2 -248 2538 -248 2538 0 FreeSans 1600 0 0 0 pc
flabel metal1 1832 1526 1832 1526 0 FreeSans 1600 0 0 0 dg
flabel metal1 -2098 -144 -2098 -144 0 FreeSans 1600 0 0 0 vssa
<< end >>
