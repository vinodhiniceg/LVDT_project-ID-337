magic
tech sky130A
timestamp 1634301196
<< error_p >>
rect 1949 19827 1978 20327
rect 2478 19827 2507 20327
rect 3007 19827 3036 20327
rect 1949 19512 1978 19780
rect 2478 19512 2507 19780
rect 3007 19512 3036 19780
rect 1963 629 1992 988
rect 2492 629 2521 988
rect 3021 629 3050 988
rect 1963 82 1992 582
rect 2492 82 2521 582
rect 3021 82 3050 582
<< error_s >>
rect 1949 19280 1978 19512
rect 2478 19280 2507 19512
rect 3007 19280 3036 19512
rect 1949 18733 1978 19233
rect 2478 18733 2507 19233
rect 3007 18733 3036 19233
rect 1949 18186 1978 18686
rect 2478 18186 2507 18686
rect 3007 18186 3036 18686
rect 1949 17639 1978 18139
rect 2478 17639 2507 18139
rect 3007 17639 3036 18139
rect 1949 16919 1978 17419
rect 2478 16919 2507 17419
rect 3007 16919 3036 17419
rect 1949 16372 1978 16872
rect 2478 16372 2507 16872
rect 3007 16372 3036 16872
rect 1949 15825 1978 16325
rect 2478 15825 2507 16325
rect 3007 15825 3036 16325
rect 1949 15278 1978 15778
rect 2478 15278 2507 15778
rect 3007 15278 3036 15778
rect 1949 14731 1978 15231
rect 2478 14731 2507 15231
rect 3007 14731 3036 15231
rect 1949 14002 1978 14502
rect 2478 14002 2507 14502
rect 3007 14002 3036 14502
rect 1949 13455 1978 13955
rect 2478 13455 2507 13955
rect 3007 13455 3036 13955
rect 1949 12908 1978 13408
rect 2478 12908 2507 13408
rect 3007 12908 3036 13408
rect 1949 12361 1978 12861
rect 2478 12361 2507 12861
rect 3007 12361 3036 12861
rect 1949 11814 1978 12314
rect 2478 11814 2507 12314
rect 3007 11814 3036 12314
rect 1949 11084 1978 11584
rect 2478 11084 2507 11584
rect 3007 11084 3036 11584
rect 1949 10537 1978 11037
rect 2478 10537 2507 11037
rect 3007 10537 3036 11037
rect 1949 9990 1978 10490
rect 2478 9990 2507 10490
rect 3007 9990 3036 10490
rect 1949 9443 1978 9943
rect 2478 9443 2507 9943
rect 3007 9443 3036 9943
rect 1949 8896 1978 9396
rect 2478 8896 2507 9396
rect 3007 8896 3036 9396
rect 1949 8152 1978 8652
rect 2478 8152 2507 8652
rect 3007 8152 3036 8652
rect 1949 7605 1978 8105
rect 2478 7605 2507 8105
rect 3007 7605 3036 8105
rect 1949 7058 1978 7558
rect 2478 7058 2507 7558
rect 3007 7058 3036 7558
rect 1949 6511 1978 7011
rect 2478 6511 2507 7011
rect 3007 6511 3036 7011
rect 1949 5964 1978 6464
rect 2478 5964 2507 6464
rect 3007 5964 3036 6464
rect 1954 5224 1983 5724
rect 2483 5224 2512 5724
rect 3012 5224 3041 5724
rect 1954 4677 1983 5177
rect 2483 4677 2512 5177
rect 3012 4677 3041 5177
rect 1954 4130 1983 4630
rect 2483 4130 2512 4630
rect 3012 4130 3041 4630
rect 1954 3583 1983 4083
rect 2483 3583 2512 4083
rect 3012 3583 3041 4083
rect 1954 3036 1983 3536
rect 2483 3036 2512 3536
rect 3012 3036 3041 3536
rect 1963 2270 1992 2770
rect 2492 2270 2521 2770
rect 3021 2270 3050 2770
rect 1963 1723 1992 2223
rect 2492 1723 2521 2223
rect 3021 1723 3050 2223
rect 1963 1176 1992 1676
rect 2492 1176 2521 1676
rect 3021 1176 3050 1676
rect 1963 988 1992 1129
rect 2492 988 2521 1129
rect 3021 988 3050 1129
use nmos5555  nmos5555_0
timestamp 1634301196
transform 1 0 376 0 1 69
box -376 -69 2845 2828
use nmos5555  nmos5555_1
timestamp 1634301196
transform 1 0 367 0 1 3023
box -376 -69 2845 2828
use nmos5555  nmos5555_2
timestamp 1634301196
transform 1 0 362 0 1 5951
box -376 -69 2845 2828
use nmos5555  nmos5555_3
timestamp 1634301196
transform 1 0 362 0 1 8883
box -376 -69 2845 2828
use nmos5555  nmos5555_4
timestamp 1634301196
transform 1 0 362 0 1 11801
box -376 -69 2845 2828
use nmos5555  nmos5555_5
timestamp 1634301196
transform 1 0 362 0 1 14718
box -376 -69 2845 2828
use nmos5555  nmos5555_6
timestamp 1634301196
transform 1 0 362 0 1 17626
box -376 -69 2845 2828
<< end >>
