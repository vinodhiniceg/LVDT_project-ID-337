magic
tech sky130A
timestamp 1634044821
<< error_s >>
rect 1873 3786 1902 4786
rect 2902 3786 2931 4786
rect 1873 2739 1902 3739
rect 2902 2739 2931 3739
rect 1873 1692 1902 2692
rect 2902 1692 2931 2692
rect 1873 645 1902 1645
rect 2902 645 2931 1645
rect 1873 -402 1902 598
rect 2902 -402 2931 598
<< pwell >>
rect -717 5029 -209 5050
rect -717 -574 3227 5029
rect -510 -585 3227 -574
<< mvpsubdiff >>
rect -683 3447 -313 3532
rect -683 3300 -640 3447
rect -683 988 -644 3300
rect -372 1135 -313 3447
rect -376 988 -313 1135
rect -683 960 -313 988
<< mvpsubdiffcont >>
rect -640 3300 -372 3447
rect -644 1135 -372 3300
rect -644 988 -376 1135
<< locali >>
rect -683 3447 -313 3532
rect -683 3300 -640 3447
rect -683 988 -644 3300
rect -372 1135 -313 3447
rect -376 988 -313 1135
rect -683 960 -313 988
<< viali >>
rect -584 1358 -435 3204
<< metal1 >>
rect -683 3204 -313 3532
rect -683 1358 -584 3204
rect -435 1358 -313 3204
rect -683 960 -313 1358
use sky130_fd_pr__nfet_g5v0d10v5_C8TC2Y  sky130_fd_pr__nfet_g5v0d10v5_C8TC2Y_0
timestamp 1634044821
transform 1 0 1373 0 1 2192
box -1558 -2607 1558 2607
<< end >>
