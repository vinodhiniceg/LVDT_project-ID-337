magic
tech sky130A
magscale 1 2
timestamp 1634904824
<< nwell >>
rect -745 -1649 745 1649
<< mvpmos >>
rect -487 1223 -287 1423
rect -229 1223 -29 1423
rect 29 1223 229 1423
rect 287 1223 487 1423
rect -487 929 -287 1129
rect -229 929 -29 1129
rect 29 929 229 1129
rect 287 929 487 1129
rect -487 635 -287 835
rect -229 635 -29 835
rect 29 635 229 835
rect 287 635 487 835
rect -487 341 -287 541
rect -229 341 -29 541
rect 29 341 229 541
rect 287 341 487 541
rect -487 47 -287 247
rect -229 47 -29 247
rect 29 47 229 247
rect 287 47 487 247
rect -487 -247 -287 -47
rect -229 -247 -29 -47
rect 29 -247 229 -47
rect 287 -247 487 -47
rect -487 -541 -287 -341
rect -229 -541 -29 -341
rect 29 -541 229 -341
rect 287 -541 487 -341
rect -487 -835 -287 -635
rect -229 -835 -29 -635
rect 29 -835 229 -635
rect 287 -835 487 -635
rect -487 -1129 -287 -929
rect -229 -1129 -29 -929
rect 29 -1129 229 -929
rect 287 -1129 487 -929
rect -487 -1423 -287 -1223
rect -229 -1423 -29 -1223
rect 29 -1423 229 -1223
rect 287 -1423 487 -1223
<< mvpdiff >>
rect -545 1349 -487 1423
rect -545 1297 -533 1349
rect -499 1297 -487 1349
rect -545 1223 -487 1297
rect -287 1349 -229 1423
rect -287 1297 -275 1349
rect -241 1297 -229 1349
rect -287 1223 -229 1297
rect -29 1349 29 1423
rect -29 1297 -17 1349
rect 17 1297 29 1349
rect -29 1223 29 1297
rect 229 1349 287 1423
rect 229 1297 241 1349
rect 275 1297 287 1349
rect 229 1223 287 1297
rect 487 1349 545 1423
rect 487 1297 499 1349
rect 533 1297 545 1349
rect 487 1223 545 1297
rect -545 1055 -487 1129
rect -545 1003 -533 1055
rect -499 1003 -487 1055
rect -545 929 -487 1003
rect -287 1055 -229 1129
rect -287 1003 -275 1055
rect -241 1003 -229 1055
rect -287 929 -229 1003
rect -29 1055 29 1129
rect -29 1003 -17 1055
rect 17 1003 29 1055
rect -29 929 29 1003
rect 229 1055 287 1129
rect 229 1003 241 1055
rect 275 1003 287 1055
rect 229 929 287 1003
rect 487 1055 545 1129
rect 487 1003 499 1055
rect 533 1003 545 1055
rect 487 929 545 1003
rect -545 761 -487 835
rect -545 709 -533 761
rect -499 709 -487 761
rect -545 635 -487 709
rect -287 761 -229 835
rect -287 709 -275 761
rect -241 709 -229 761
rect -287 635 -229 709
rect -29 761 29 835
rect -29 709 -17 761
rect 17 709 29 761
rect -29 635 29 709
rect 229 761 287 835
rect 229 709 241 761
rect 275 709 287 761
rect 229 635 287 709
rect 487 761 545 835
rect 487 709 499 761
rect 533 709 545 761
rect 487 635 545 709
rect -545 467 -487 541
rect -545 415 -533 467
rect -499 415 -487 467
rect -545 341 -487 415
rect -287 467 -229 541
rect -287 415 -275 467
rect -241 415 -229 467
rect -287 341 -229 415
rect -29 467 29 541
rect -29 415 -17 467
rect 17 415 29 467
rect -29 341 29 415
rect 229 467 287 541
rect 229 415 241 467
rect 275 415 287 467
rect 229 341 287 415
rect 487 467 545 541
rect 487 415 499 467
rect 533 415 545 467
rect 487 341 545 415
rect -545 173 -487 247
rect -545 121 -533 173
rect -499 121 -487 173
rect -545 47 -487 121
rect -287 173 -229 247
rect -287 121 -275 173
rect -241 121 -229 173
rect -287 47 -229 121
rect -29 173 29 247
rect -29 121 -17 173
rect 17 121 29 173
rect -29 47 29 121
rect 229 173 287 247
rect 229 121 241 173
rect 275 121 287 173
rect 229 47 287 121
rect 487 173 545 247
rect 487 121 499 173
rect 533 121 545 173
rect 487 47 545 121
rect -545 -121 -487 -47
rect -545 -173 -533 -121
rect -499 -173 -487 -121
rect -545 -247 -487 -173
rect -287 -121 -229 -47
rect -287 -173 -275 -121
rect -241 -173 -229 -121
rect -287 -247 -229 -173
rect -29 -121 29 -47
rect -29 -173 -17 -121
rect 17 -173 29 -121
rect -29 -247 29 -173
rect 229 -121 287 -47
rect 229 -173 241 -121
rect 275 -173 287 -121
rect 229 -247 287 -173
rect 487 -121 545 -47
rect 487 -173 499 -121
rect 533 -173 545 -121
rect 487 -247 545 -173
rect -545 -415 -487 -341
rect -545 -467 -533 -415
rect -499 -467 -487 -415
rect -545 -541 -487 -467
rect -287 -415 -229 -341
rect -287 -467 -275 -415
rect -241 -467 -229 -415
rect -287 -541 -229 -467
rect -29 -415 29 -341
rect -29 -467 -17 -415
rect 17 -467 29 -415
rect -29 -541 29 -467
rect 229 -415 287 -341
rect 229 -467 241 -415
rect 275 -467 287 -415
rect 229 -541 287 -467
rect 487 -415 545 -341
rect 487 -467 499 -415
rect 533 -467 545 -415
rect 487 -541 545 -467
rect -545 -709 -487 -635
rect -545 -761 -533 -709
rect -499 -761 -487 -709
rect -545 -835 -487 -761
rect -287 -709 -229 -635
rect -287 -761 -275 -709
rect -241 -761 -229 -709
rect -287 -835 -229 -761
rect -29 -709 29 -635
rect -29 -761 -17 -709
rect 17 -761 29 -709
rect -29 -835 29 -761
rect 229 -709 287 -635
rect 229 -761 241 -709
rect 275 -761 287 -709
rect 229 -835 287 -761
rect 487 -709 545 -635
rect 487 -761 499 -709
rect 533 -761 545 -709
rect 487 -835 545 -761
rect -545 -1003 -487 -929
rect -545 -1055 -533 -1003
rect -499 -1055 -487 -1003
rect -545 -1129 -487 -1055
rect -287 -1003 -229 -929
rect -287 -1055 -275 -1003
rect -241 -1055 -229 -1003
rect -287 -1129 -229 -1055
rect -29 -1003 29 -929
rect -29 -1055 -17 -1003
rect 17 -1055 29 -1003
rect -29 -1129 29 -1055
rect 229 -1003 287 -929
rect 229 -1055 241 -1003
rect 275 -1055 287 -1003
rect 229 -1129 287 -1055
rect 487 -1003 545 -929
rect 487 -1055 499 -1003
rect 533 -1055 545 -1003
rect 487 -1129 545 -1055
rect -545 -1297 -487 -1223
rect -545 -1349 -533 -1297
rect -499 -1349 -487 -1297
rect -545 -1423 -487 -1349
rect -287 -1297 -229 -1223
rect -287 -1349 -275 -1297
rect -241 -1349 -229 -1297
rect -287 -1423 -229 -1349
rect -29 -1297 29 -1223
rect -29 -1349 -17 -1297
rect 17 -1349 29 -1297
rect -29 -1423 29 -1349
rect 229 -1297 287 -1223
rect 229 -1349 241 -1297
rect 275 -1349 287 -1297
rect 229 -1423 287 -1349
rect 487 -1297 545 -1223
rect 487 -1349 499 -1297
rect 533 -1349 545 -1297
rect 487 -1423 545 -1349
<< mvpdiffc >>
rect -533 1297 -499 1349
rect -275 1297 -241 1349
rect -17 1297 17 1349
rect 241 1297 275 1349
rect 499 1297 533 1349
rect -533 1003 -499 1055
rect -275 1003 -241 1055
rect -17 1003 17 1055
rect 241 1003 275 1055
rect 499 1003 533 1055
rect -533 709 -499 761
rect -275 709 -241 761
rect -17 709 17 761
rect 241 709 275 761
rect 499 709 533 761
rect -533 415 -499 467
rect -275 415 -241 467
rect -17 415 17 467
rect 241 415 275 467
rect 499 415 533 467
rect -533 121 -499 173
rect -275 121 -241 173
rect -17 121 17 173
rect 241 121 275 173
rect 499 121 533 173
rect -533 -173 -499 -121
rect -275 -173 -241 -121
rect -17 -173 17 -121
rect 241 -173 275 -121
rect 499 -173 533 -121
rect -533 -467 -499 -415
rect -275 -467 -241 -415
rect -17 -467 17 -415
rect 241 -467 275 -415
rect 499 -467 533 -415
rect -533 -761 -499 -709
rect -275 -761 -241 -709
rect -17 -761 17 -709
rect 241 -761 275 -709
rect 499 -761 533 -709
rect -533 -1055 -499 -1003
rect -275 -1055 -241 -1003
rect -17 -1055 17 -1003
rect 241 -1055 275 -1003
rect 499 -1055 533 -1003
rect -533 -1349 -499 -1297
rect -275 -1349 -241 -1297
rect -17 -1349 17 -1297
rect 241 -1349 275 -1297
rect 499 -1349 533 -1297
<< mvnsubdiff >>
rect -679 1525 679 1583
rect -679 738 -621 1525
rect -679 -738 -667 738
rect -633 -738 -621 738
rect 621 738 679 1525
rect -679 -1525 -621 -738
rect 621 -738 633 738
rect 667 -738 679 738
rect 621 -1525 679 -738
rect -679 -1583 679 -1525
<< mvnsubdiffcont >>
rect -667 -738 -633 738
rect 633 -738 667 738
<< poly >>
rect -487 1423 -287 1449
rect -229 1423 -29 1449
rect 29 1423 229 1449
rect 287 1423 487 1449
rect -487 1197 -287 1223
rect -229 1197 -29 1223
rect 29 1197 229 1223
rect 287 1197 487 1223
rect -487 1129 -287 1155
rect -229 1129 -29 1155
rect 29 1129 229 1155
rect 287 1129 487 1155
rect -487 903 -287 929
rect -229 903 -29 929
rect 29 903 229 929
rect 287 903 487 929
rect -487 835 -287 861
rect -229 835 -29 861
rect 29 835 229 861
rect 287 835 487 861
rect -487 609 -287 635
rect -229 609 -29 635
rect 29 609 229 635
rect 287 609 487 635
rect -487 541 -287 567
rect -229 541 -29 567
rect 29 541 229 567
rect 287 541 487 567
rect -487 315 -287 341
rect -229 315 -29 341
rect 29 315 229 341
rect 287 315 487 341
rect -487 247 -287 273
rect -229 247 -29 273
rect 29 247 229 273
rect 287 247 487 273
rect -487 21 -287 47
rect -229 21 -29 47
rect 29 21 229 47
rect 287 21 487 47
rect -487 -47 -287 -21
rect -229 -47 -29 -21
rect 29 -47 229 -21
rect 287 -47 487 -21
rect -487 -273 -287 -247
rect -229 -273 -29 -247
rect 29 -273 229 -247
rect 287 -273 487 -247
rect -487 -341 -287 -315
rect -229 -341 -29 -315
rect 29 -341 229 -315
rect 287 -341 487 -315
rect -487 -567 -287 -541
rect -229 -567 -29 -541
rect 29 -567 229 -541
rect 287 -567 487 -541
rect -487 -635 -287 -609
rect -229 -635 -29 -609
rect 29 -635 229 -609
rect 287 -635 487 -609
rect -487 -861 -287 -835
rect -229 -861 -29 -835
rect 29 -861 229 -835
rect 287 -861 487 -835
rect -487 -929 -287 -903
rect -229 -929 -29 -903
rect 29 -929 229 -903
rect 287 -929 487 -903
rect -487 -1155 -287 -1129
rect -229 -1155 -29 -1129
rect 29 -1155 229 -1129
rect 287 -1155 487 -1129
rect -487 -1223 -287 -1197
rect -229 -1223 -29 -1197
rect 29 -1223 229 -1197
rect 287 -1223 487 -1197
rect -487 -1449 -287 -1423
rect -229 -1449 -29 -1423
rect 29 -1449 229 -1423
rect 287 -1449 487 -1423
<< locali >>
rect -533 1349 -499 1365
rect -533 1281 -499 1297
rect -275 1349 -241 1365
rect -275 1281 -241 1297
rect -17 1349 17 1365
rect -17 1281 17 1297
rect 241 1349 275 1365
rect 241 1281 275 1297
rect 499 1349 533 1365
rect 499 1281 533 1297
rect -533 1055 -499 1071
rect -533 987 -499 1003
rect -275 1055 -241 1071
rect -275 987 -241 1003
rect -17 1055 17 1071
rect -17 987 17 1003
rect 241 1055 275 1071
rect 241 987 275 1003
rect 499 1055 533 1071
rect 499 987 533 1003
rect -533 761 -499 777
rect -667 738 -633 754
rect -533 693 -499 709
rect -275 761 -241 777
rect -275 693 -241 709
rect -17 761 17 777
rect -17 693 17 709
rect 241 761 275 777
rect 241 693 275 709
rect 499 761 533 777
rect 499 693 533 709
rect 633 738 667 754
rect -533 467 -499 483
rect -533 399 -499 415
rect -275 467 -241 483
rect -275 399 -241 415
rect -17 467 17 483
rect -17 399 17 415
rect 241 467 275 483
rect 241 399 275 415
rect 499 467 533 483
rect 499 399 533 415
rect -533 173 -499 189
rect -533 105 -499 121
rect -275 173 -241 189
rect -275 105 -241 121
rect -17 173 17 189
rect -17 105 17 121
rect 241 173 275 189
rect 241 105 275 121
rect 499 173 533 189
rect 499 105 533 121
rect -533 -121 -499 -105
rect -533 -189 -499 -173
rect -275 -121 -241 -105
rect -275 -189 -241 -173
rect -17 -121 17 -105
rect -17 -189 17 -173
rect 241 -121 275 -105
rect 241 -189 275 -173
rect 499 -121 533 -105
rect 499 -189 533 -173
rect -533 -415 -499 -399
rect -533 -483 -499 -467
rect -275 -415 -241 -399
rect -275 -483 -241 -467
rect -17 -415 17 -399
rect -17 -483 17 -467
rect 241 -415 275 -399
rect 241 -483 275 -467
rect 499 -415 533 -399
rect 499 -483 533 -467
rect -667 -754 -633 -738
rect -533 -709 -499 -693
rect -533 -777 -499 -761
rect -275 -709 -241 -693
rect -275 -777 -241 -761
rect -17 -709 17 -693
rect -17 -777 17 -761
rect 241 -709 275 -693
rect 241 -777 275 -761
rect 499 -709 533 -693
rect 633 -754 667 -738
rect 499 -777 533 -761
rect -533 -1003 -499 -987
rect -533 -1071 -499 -1055
rect -275 -1003 -241 -987
rect -275 -1071 -241 -1055
rect -17 -1003 17 -987
rect -17 -1071 17 -1055
rect 241 -1003 275 -987
rect 241 -1071 275 -1055
rect 499 -1003 533 -987
rect 499 -1071 533 -1055
rect -533 -1297 -499 -1281
rect -533 -1365 -499 -1349
rect -275 -1297 -241 -1281
rect -275 -1365 -241 -1349
rect -17 -1297 17 -1281
rect -17 -1365 17 -1349
rect 241 -1297 275 -1281
rect 241 -1365 275 -1349
rect 499 -1297 533 -1281
rect 499 -1365 533 -1349
<< viali >>
rect -533 1297 -499 1349
rect -275 1297 -241 1349
rect -17 1297 17 1349
rect 241 1297 275 1349
rect 499 1297 533 1349
rect -533 1003 -499 1055
rect -275 1003 -241 1055
rect -17 1003 17 1055
rect 241 1003 275 1055
rect 499 1003 533 1055
rect -533 709 -499 761
rect -275 709 -241 761
rect -17 709 17 761
rect 241 709 275 761
rect 499 709 533 761
rect -533 415 -499 467
rect -275 415 -241 467
rect -17 415 17 467
rect 241 415 275 467
rect 499 415 533 467
rect -533 121 -499 173
rect -275 121 -241 173
rect -17 121 17 173
rect 241 121 275 173
rect 499 121 533 173
rect -533 -173 -499 -121
rect -275 -173 -241 -121
rect -17 -173 17 -121
rect 241 -173 275 -121
rect 499 -173 533 -121
rect -533 -467 -499 -415
rect -275 -467 -241 -415
rect -17 -467 17 -415
rect 241 -467 275 -415
rect 499 -467 533 -415
rect -533 -761 -499 -709
rect -275 -761 -241 -709
rect -17 -761 17 -709
rect 241 -761 275 -709
rect 499 -761 533 -709
rect -533 -1055 -499 -1003
rect -275 -1055 -241 -1003
rect -17 -1055 17 -1003
rect 241 -1055 275 -1003
rect 499 -1055 533 -1003
rect -533 -1349 -499 -1297
rect -275 -1349 -241 -1297
rect -17 -1349 17 -1297
rect 241 -1349 275 -1297
rect 499 -1349 533 -1297
<< metal1 >>
rect -539 1349 -493 1361
rect -539 1297 -533 1349
rect -499 1297 -493 1349
rect -539 1285 -493 1297
rect -281 1349 -235 1361
rect -281 1297 -275 1349
rect -241 1297 -235 1349
rect -281 1285 -235 1297
rect -23 1349 23 1361
rect -23 1297 -17 1349
rect 17 1297 23 1349
rect -23 1285 23 1297
rect 235 1349 281 1361
rect 235 1297 241 1349
rect 275 1297 281 1349
rect 235 1285 281 1297
rect 493 1349 539 1361
rect 493 1297 499 1349
rect 533 1297 539 1349
rect 493 1285 539 1297
rect -539 1055 -493 1067
rect -539 1003 -533 1055
rect -499 1003 -493 1055
rect -539 991 -493 1003
rect -281 1055 -235 1067
rect -281 1003 -275 1055
rect -241 1003 -235 1055
rect -281 991 -235 1003
rect -23 1055 23 1067
rect -23 1003 -17 1055
rect 17 1003 23 1055
rect -23 991 23 1003
rect 235 1055 281 1067
rect 235 1003 241 1055
rect 275 1003 281 1055
rect 235 991 281 1003
rect 493 1055 539 1067
rect 493 1003 499 1055
rect 533 1003 539 1055
rect 493 991 539 1003
rect -539 761 -493 773
rect -539 709 -533 761
rect -499 709 -493 761
rect -539 697 -493 709
rect -281 761 -235 773
rect -281 709 -275 761
rect -241 709 -235 761
rect -281 697 -235 709
rect -23 761 23 773
rect -23 709 -17 761
rect 17 709 23 761
rect -23 697 23 709
rect 235 761 281 773
rect 235 709 241 761
rect 275 709 281 761
rect 235 697 281 709
rect 493 761 539 773
rect 493 709 499 761
rect 533 709 539 761
rect 493 697 539 709
rect -539 467 -493 479
rect -539 415 -533 467
rect -499 415 -493 467
rect -539 403 -493 415
rect -281 467 -235 479
rect -281 415 -275 467
rect -241 415 -235 467
rect -281 403 -235 415
rect -23 467 23 479
rect -23 415 -17 467
rect 17 415 23 467
rect -23 403 23 415
rect 235 467 281 479
rect 235 415 241 467
rect 275 415 281 467
rect 235 403 281 415
rect 493 467 539 479
rect 493 415 499 467
rect 533 415 539 467
rect 493 403 539 415
rect -539 173 -493 185
rect -539 121 -533 173
rect -499 121 -493 173
rect -539 109 -493 121
rect -281 173 -235 185
rect -281 121 -275 173
rect -241 121 -235 173
rect -281 109 -235 121
rect -23 173 23 185
rect -23 121 -17 173
rect 17 121 23 173
rect -23 109 23 121
rect 235 173 281 185
rect 235 121 241 173
rect 275 121 281 173
rect 235 109 281 121
rect 493 173 539 185
rect 493 121 499 173
rect 533 121 539 173
rect 493 109 539 121
rect -539 -121 -493 -109
rect -539 -173 -533 -121
rect -499 -173 -493 -121
rect -539 -185 -493 -173
rect -281 -121 -235 -109
rect -281 -173 -275 -121
rect -241 -173 -235 -121
rect -281 -185 -235 -173
rect -23 -121 23 -109
rect -23 -173 -17 -121
rect 17 -173 23 -121
rect -23 -185 23 -173
rect 235 -121 281 -109
rect 235 -173 241 -121
rect 275 -173 281 -121
rect 235 -185 281 -173
rect 493 -121 539 -109
rect 493 -173 499 -121
rect 533 -173 539 -121
rect 493 -185 539 -173
rect -539 -415 -493 -403
rect -539 -467 -533 -415
rect -499 -467 -493 -415
rect -539 -479 -493 -467
rect -281 -415 -235 -403
rect -281 -467 -275 -415
rect -241 -467 -235 -415
rect -281 -479 -235 -467
rect -23 -415 23 -403
rect -23 -467 -17 -415
rect 17 -467 23 -415
rect -23 -479 23 -467
rect 235 -415 281 -403
rect 235 -467 241 -415
rect 275 -467 281 -415
rect 235 -479 281 -467
rect 493 -415 539 -403
rect 493 -467 499 -415
rect 533 -467 539 -415
rect 493 -479 539 -467
rect -539 -709 -493 -697
rect -539 -761 -533 -709
rect -499 -761 -493 -709
rect -539 -773 -493 -761
rect -281 -709 -235 -697
rect -281 -761 -275 -709
rect -241 -761 -235 -709
rect -281 -773 -235 -761
rect -23 -709 23 -697
rect -23 -761 -17 -709
rect 17 -761 23 -709
rect -23 -773 23 -761
rect 235 -709 281 -697
rect 235 -761 241 -709
rect 275 -761 281 -709
rect 235 -773 281 -761
rect 493 -709 539 -697
rect 493 -761 499 -709
rect 533 -761 539 -709
rect 493 -773 539 -761
rect -539 -1003 -493 -991
rect -539 -1055 -533 -1003
rect -499 -1055 -493 -1003
rect -539 -1067 -493 -1055
rect -281 -1003 -235 -991
rect -281 -1055 -275 -1003
rect -241 -1055 -235 -1003
rect -281 -1067 -235 -1055
rect -23 -1003 23 -991
rect -23 -1055 -17 -1003
rect 17 -1055 23 -1003
rect -23 -1067 23 -1055
rect 235 -1003 281 -991
rect 235 -1055 241 -1003
rect 275 -1055 281 -1003
rect 235 -1067 281 -1055
rect 493 -1003 539 -991
rect 493 -1055 499 -1003
rect 533 -1055 539 -1003
rect 493 -1067 539 -1055
rect -539 -1297 -493 -1285
rect -539 -1349 -533 -1297
rect -499 -1349 -493 -1297
rect -539 -1361 -493 -1349
rect -281 -1297 -235 -1285
rect -281 -1349 -275 -1297
rect -241 -1349 -235 -1297
rect -281 -1361 -235 -1349
rect -23 -1297 23 -1285
rect -23 -1349 -17 -1297
rect 17 -1349 23 -1297
rect -23 -1361 23 -1349
rect 235 -1297 281 -1285
rect 235 -1349 241 -1297
rect 275 -1349 281 -1297
rect 235 -1361 281 -1349
rect 493 -1297 539 -1285
rect 493 -1349 499 -1297
rect 533 -1349 539 -1297
rect 493 -1361 539 -1349
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string FIXED_BBOX -650 -1554 650 1554
string parameters w 1 l 1 m 10 nf 4 diffcov 30 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 50 rlcov 50 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 30 viadrn 30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
