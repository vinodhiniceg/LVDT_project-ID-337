magic
tech sky130A
timestamp 1634132563
<< mvnmos >>
rect -808 544 -508 844
rect -479 544 -179 844
rect -150 544 150 844
rect 179 544 479 844
rect 508 544 808 844
rect -808 197 -508 497
rect -479 197 -179 497
rect -150 197 150 497
rect 179 197 479 497
rect 508 197 808 497
rect -808 -150 -508 150
rect -479 -150 -179 150
rect -150 -150 150 150
rect 179 -150 479 150
rect 508 -150 808 150
rect -808 -497 -508 -197
rect -479 -497 -179 -197
rect -150 -497 150 -197
rect 179 -497 479 -197
rect 508 -497 808 -197
rect -808 -844 -508 -544
rect -479 -844 -179 -544
rect -150 -844 150 -544
rect 179 -844 479 -544
rect 508 -844 808 -544
<< mvndiff >>
rect -837 737 -808 844
rect -837 651 -831 737
rect -814 651 -808 737
rect -837 544 -808 651
rect -508 737 -479 844
rect -508 651 -502 737
rect -485 651 -479 737
rect -508 544 -479 651
rect -179 737 -150 844
rect -179 651 -173 737
rect -156 651 -150 737
rect -179 544 -150 651
rect 150 737 179 844
rect 150 651 156 737
rect 173 651 179 737
rect 150 544 179 651
rect 479 737 508 844
rect 479 651 485 737
rect 502 651 508 737
rect 479 544 508 651
rect 808 737 837 844
rect 808 651 814 737
rect 831 651 837 737
rect 808 544 837 651
rect -837 390 -808 497
rect -837 304 -831 390
rect -814 304 -808 390
rect -837 197 -808 304
rect -508 390 -479 497
rect -508 304 -502 390
rect -485 304 -479 390
rect -508 197 -479 304
rect -179 390 -150 497
rect -179 304 -173 390
rect -156 304 -150 390
rect -179 197 -150 304
rect 150 390 179 497
rect 150 304 156 390
rect 173 304 179 390
rect 150 197 179 304
rect 479 390 508 497
rect 479 304 485 390
rect 502 304 508 390
rect 479 197 508 304
rect 808 390 837 497
rect 808 304 814 390
rect 831 304 837 390
rect 808 197 837 304
rect -837 43 -808 150
rect -837 -43 -831 43
rect -814 -43 -808 43
rect -837 -150 -808 -43
rect -508 43 -479 150
rect -508 -43 -502 43
rect -485 -43 -479 43
rect -508 -150 -479 -43
rect -179 43 -150 150
rect -179 -43 -173 43
rect -156 -43 -150 43
rect -179 -150 -150 -43
rect 150 43 179 150
rect 150 -43 156 43
rect 173 -43 179 43
rect 150 -150 179 -43
rect 479 43 508 150
rect 479 -43 485 43
rect 502 -43 508 43
rect 479 -150 508 -43
rect 808 43 837 150
rect 808 -43 814 43
rect 831 -43 837 43
rect 808 -150 837 -43
rect -837 -304 -808 -197
rect -837 -390 -831 -304
rect -814 -390 -808 -304
rect -837 -497 -808 -390
rect -508 -304 -479 -197
rect -508 -390 -502 -304
rect -485 -390 -479 -304
rect -508 -497 -479 -390
rect -179 -304 -150 -197
rect -179 -390 -173 -304
rect -156 -390 -150 -304
rect -179 -497 -150 -390
rect 150 -304 179 -197
rect 150 -390 156 -304
rect 173 -390 179 -304
rect 150 -497 179 -390
rect 479 -304 508 -197
rect 479 -390 485 -304
rect 502 -390 508 -304
rect 479 -497 508 -390
rect 808 -304 837 -197
rect 808 -390 814 -304
rect 831 -390 837 -304
rect 808 -497 837 -390
rect -837 -651 -808 -544
rect -837 -737 -831 -651
rect -814 -737 -808 -651
rect -837 -844 -808 -737
rect -508 -651 -479 -544
rect -508 -737 -502 -651
rect -485 -737 -479 -651
rect -508 -844 -479 -737
rect -179 -651 -150 -544
rect -179 -737 -173 -651
rect -156 -737 -150 -651
rect -179 -844 -150 -737
rect 150 -651 179 -544
rect 150 -737 156 -651
rect 173 -737 179 -651
rect 150 -844 179 -737
rect 479 -651 508 -544
rect 479 -737 485 -651
rect 502 -737 508 -651
rect 479 -844 508 -737
rect 808 -651 837 -544
rect 808 -737 814 -651
rect 831 -737 837 -651
rect 808 -844 837 -737
<< mvndiffc >>
rect -831 651 -814 737
rect -502 651 -485 737
rect -173 651 -156 737
rect 156 651 173 737
rect 485 651 502 737
rect 814 651 831 737
rect -831 304 -814 390
rect -502 304 -485 390
rect -173 304 -156 390
rect 156 304 173 390
rect 485 304 502 390
rect 814 304 831 390
rect -831 -43 -814 43
rect -502 -43 -485 43
rect -173 -43 -156 43
rect 156 -43 173 43
rect 485 -43 502 43
rect 814 -43 831 43
rect -831 -390 -814 -304
rect -502 -390 -485 -304
rect -173 -390 -156 -304
rect 156 -390 173 -304
rect 485 -390 502 -304
rect 814 -390 831 -304
rect -831 -737 -814 -651
rect -502 -737 -485 -651
rect -173 -737 -156 -651
rect 156 -737 173 -651
rect 485 -737 502 -651
rect 814 -737 831 -651
<< poly >>
rect -808 844 -508 857
rect -479 844 -179 857
rect -150 844 150 857
rect 179 844 479 857
rect 508 844 808 857
rect -808 531 -508 544
rect -479 531 -179 544
rect -150 531 150 544
rect 179 531 479 544
rect 508 531 808 544
rect -808 497 -508 510
rect -479 497 -179 510
rect -150 497 150 510
rect 179 497 479 510
rect 508 497 808 510
rect -808 184 -508 197
rect -479 184 -179 197
rect -150 184 150 197
rect 179 184 479 197
rect 508 184 808 197
rect -808 150 -508 163
rect -479 150 -179 163
rect -150 150 150 163
rect 179 150 479 163
rect 508 150 808 163
rect -808 -163 -508 -150
rect -479 -163 -179 -150
rect -150 -163 150 -150
rect 179 -163 479 -150
rect 508 -163 808 -150
rect -808 -197 -508 -184
rect -479 -197 -179 -184
rect -150 -197 150 -184
rect 179 -197 479 -184
rect 508 -197 808 -184
rect -808 -510 -508 -497
rect -479 -510 -179 -497
rect -150 -510 150 -497
rect 179 -510 479 -497
rect 508 -510 808 -497
rect -808 -544 -508 -531
rect -479 -544 -179 -531
rect -150 -544 150 -531
rect 179 -544 479 -531
rect 508 -544 808 -531
rect -808 -857 -508 -844
rect -479 -857 -179 -844
rect -150 -857 150 -844
rect 179 -857 479 -844
rect 508 -857 808 -844
<< locali >>
rect -831 737 -814 745
rect -831 643 -814 651
rect -502 737 -485 745
rect -502 643 -485 651
rect -173 737 -156 745
rect -173 643 -156 651
rect 156 737 173 745
rect 156 643 173 651
rect 485 737 502 745
rect 485 643 502 651
rect 814 737 831 745
rect 814 643 831 651
rect -831 390 -814 398
rect -831 296 -814 304
rect -502 390 -485 398
rect -502 296 -485 304
rect -173 390 -156 398
rect -173 296 -156 304
rect 156 390 173 398
rect 156 296 173 304
rect 485 390 502 398
rect 485 296 502 304
rect 814 390 831 398
rect 814 296 831 304
rect -831 43 -814 51
rect -831 -51 -814 -43
rect -502 43 -485 51
rect -502 -51 -485 -43
rect -173 43 -156 51
rect -173 -51 -156 -43
rect 156 43 173 51
rect 156 -51 173 -43
rect 485 43 502 51
rect 485 -51 502 -43
rect 814 43 831 51
rect 814 -51 831 -43
rect -831 -304 -814 -296
rect -831 -398 -814 -390
rect -502 -304 -485 -296
rect -502 -398 -485 -390
rect -173 -304 -156 -296
rect -173 -398 -156 -390
rect 156 -304 173 -296
rect 156 -398 173 -390
rect 485 -304 502 -296
rect 485 -398 502 -390
rect 814 -304 831 -296
rect 814 -398 831 -390
rect -831 -651 -814 -643
rect -831 -745 -814 -737
rect -502 -651 -485 -643
rect -502 -745 -485 -737
rect -173 -651 -156 -643
rect -173 -745 -156 -737
rect 156 -651 173 -643
rect 156 -745 173 -737
rect 485 -651 502 -643
rect 485 -745 502 -737
rect 814 -651 831 -643
rect 814 -745 831 -737
<< viali >>
rect -831 651 -814 737
rect -502 651 -485 737
rect -173 651 -156 737
rect 156 651 173 737
rect 485 651 502 737
rect 814 651 831 737
rect -831 304 -814 390
rect -502 304 -485 390
rect -173 304 -156 390
rect 156 304 173 390
rect 485 304 502 390
rect 814 304 831 390
rect -831 -43 -814 43
rect -502 -43 -485 43
rect -173 -43 -156 43
rect 156 -43 173 43
rect 485 -43 502 43
rect 814 -43 831 43
rect -831 -390 -814 -304
rect -502 -390 -485 -304
rect -173 -390 -156 -304
rect 156 -390 173 -304
rect 485 -390 502 -304
rect 814 -390 831 -304
rect -831 -737 -814 -651
rect -502 -737 -485 -651
rect -173 -737 -156 -651
rect 156 -737 173 -651
rect 485 -737 502 -651
rect 814 -737 831 -651
<< metal1 >>
rect -834 737 -811 743
rect -834 651 -831 737
rect -814 651 -811 737
rect -834 645 -811 651
rect -505 737 -482 743
rect -505 651 -502 737
rect -485 651 -482 737
rect -505 645 -482 651
rect -176 737 -153 743
rect -176 651 -173 737
rect -156 651 -153 737
rect -176 645 -153 651
rect 153 737 176 743
rect 153 651 156 737
rect 173 651 176 737
rect 153 645 176 651
rect 482 737 505 743
rect 482 651 485 737
rect 502 651 505 737
rect 482 645 505 651
rect 811 737 834 743
rect 811 651 814 737
rect 831 651 834 737
rect 811 645 834 651
rect -834 390 -811 396
rect -834 304 -831 390
rect -814 304 -811 390
rect -834 298 -811 304
rect -505 390 -482 396
rect -505 304 -502 390
rect -485 304 -482 390
rect -505 298 -482 304
rect -176 390 -153 396
rect -176 304 -173 390
rect -156 304 -153 390
rect -176 298 -153 304
rect 153 390 176 396
rect 153 304 156 390
rect 173 304 176 390
rect 153 298 176 304
rect 482 390 505 396
rect 482 304 485 390
rect 502 304 505 390
rect 482 298 505 304
rect 811 390 834 396
rect 811 304 814 390
rect 831 304 834 390
rect 811 298 834 304
rect -834 43 -811 49
rect -834 -43 -831 43
rect -814 -43 -811 43
rect -834 -49 -811 -43
rect -505 43 -482 49
rect -505 -43 -502 43
rect -485 -43 -482 43
rect -505 -49 -482 -43
rect -176 43 -153 49
rect -176 -43 -173 43
rect -156 -43 -153 43
rect -176 -49 -153 -43
rect 153 43 176 49
rect 153 -43 156 43
rect 173 -43 176 43
rect 153 -49 176 -43
rect 482 43 505 49
rect 482 -43 485 43
rect 502 -43 505 43
rect 482 -49 505 -43
rect 811 43 834 49
rect 811 -43 814 43
rect 831 -43 834 43
rect 811 -49 834 -43
rect -834 -304 -811 -298
rect -834 -390 -831 -304
rect -814 -390 -811 -304
rect -834 -396 -811 -390
rect -505 -304 -482 -298
rect -505 -390 -502 -304
rect -485 -390 -482 -304
rect -505 -396 -482 -390
rect -176 -304 -153 -298
rect -176 -390 -173 -304
rect -156 -390 -153 -304
rect -176 -396 -153 -390
rect 153 -304 176 -298
rect 153 -390 156 -304
rect 173 -390 176 -304
rect 153 -396 176 -390
rect 482 -304 505 -298
rect 482 -390 485 -304
rect 502 -390 505 -304
rect 482 -396 505 -390
rect 811 -304 834 -298
rect 811 -390 814 -304
rect 831 -390 834 -304
rect 811 -396 834 -390
rect -834 -651 -811 -645
rect -834 -737 -831 -651
rect -814 -737 -811 -651
rect -834 -743 -811 -737
rect -505 -651 -482 -645
rect -505 -737 -502 -651
rect -485 -737 -482 -651
rect -505 -743 -482 -737
rect -176 -651 -153 -645
rect -176 -737 -173 -651
rect -156 -737 -153 -651
rect -176 -743 -153 -737
rect 153 -651 176 -645
rect 153 -737 156 -651
rect 173 -737 176 -651
rect 153 -743 176 -737
rect 482 -651 505 -645
rect 482 -737 485 -651
rect 502 -737 505 -651
rect 482 -743 505 -737
rect 811 -651 834 -645
rect 811 -737 814 -651
rect 831 -737 834 -651
rect 811 -743 834 -737
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string parameters w 3 l 3 m 5 nf 5 diffcov 30 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 30 viadrn 30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
