magic
tech sky130A
timestamp 1634186000
<< mvnsubdiff >>
rect 79 279 357 8202
rect 12877 7766 13155 8132
rect 12877 6387 12956 7766
rect 13068 6387 13155 7766
rect 12877 5819 13155 6387
rect 12877 4558 12962 5819
rect 13075 4558 13155 5819
rect 12877 3839 13155 4558
rect 12877 2493 12943 3839
rect 13075 2493 13155 3839
rect 12877 1615 13155 2493
rect 12877 546 12949 1615
rect 13081 546 13155 1615
rect 12877 209 13155 546
<< mvnsubdiffcont >>
rect 12956 6387 13068 7766
rect 12962 4558 13075 5819
rect 12943 2493 13075 3839
rect 12949 546 13081 1615
<< poly >>
rect 6281 8064 6908 8214
rect 1898 3966 1899 3981
rect 3996 3955 3997 3976
rect 6234 3956 6235 3971
rect 8332 3945 8333 3966
rect 10528 3928 10529 3943
rect 12626 3917 12627 3938
<< polycont >>
rect 2171 8018 2313 8090
rect 10844 7976 11045 8049
<< locali >>
rect 2156 8090 2328 8098
rect 2156 8018 2171 8090
rect 2313 8018 2328 8090
rect 2156 8009 2328 8018
rect 2208 7915 2275 8009
rect 4149 7965 4211 7991
rect 3828 7888 4211 7965
rect 4149 7826 4211 7888
rect 4744 7867 4822 8141
rect 4149 7743 4615 7826
rect 8470 7758 8584 8209
rect 10807 8049 11078 8063
rect 10807 7976 10844 8049
rect 11045 7976 11078 8049
rect 10807 7968 11078 7976
rect 10880 7882 11005 7968
rect 12776 7914 12828 7929
rect 12440 7846 12828 7914
rect 12776 7769 12828 7846
rect 12923 7769 13101 7799
rect 12771 7766 13112 7769
rect 12771 7675 12956 7766
rect 12923 6387 12956 7675
rect 13068 7675 13112 7766
rect 13068 6387 13101 7675
rect 12923 6340 13101 6387
rect 4465 5740 4677 6035
rect 12929 5819 13108 5885
rect 12929 4558 12962 5819
rect 13075 4558 13108 5819
rect 12929 4466 13108 4558
rect 12923 3839 13101 3872
rect 12923 2493 12943 3839
rect 13075 2493 13101 3839
rect 12923 2427 13101 2493
rect 12903 1615 13114 1655
rect 12903 546 12949 1615
rect 13081 546 13114 1615
rect 12903 473 13114 546
<< viali >>
rect 2201 8033 2291 8085
rect 10868 7981 11019 8043
rect 12962 6433 13055 7707
rect 12989 4585 13055 5779
rect 12969 2598 13048 3780
rect 12976 599 13035 1556
<< metal1 >>
rect 2156 8085 2328 8098
rect 2156 8033 2201 8085
rect 2291 8033 2328 8085
rect 2156 8009 2328 8033
rect 10807 8043 11078 8063
rect 10807 7981 10868 8043
rect 11019 7981 11078 8043
rect 10807 7968 11078 7981
rect 12923 7707 13101 7799
rect 12923 6433 12962 7707
rect 13055 6433 13101 7707
rect 12923 6340 13101 6433
rect 12929 5779 13108 5885
rect 12929 4585 12989 5779
rect 13055 4585 13108 5779
rect 12929 4466 13108 4585
rect 12923 3780 13101 3872
rect 12923 2598 12969 3780
rect 13048 2598 13101 3780
rect 12923 2427 13101 2598
rect 12903 1556 13114 1655
rect 12903 599 12976 1556
rect 13035 599 13114 1556
rect 12903 473 13114 599
use pmos331020  pmos331020_0
timestamp 1634181701
transform 1 0 113 0 1 50
box -113 -50 4688 8286
use pmos331020  pmos331020_1
timestamp 1634181701
transform 1 0 4449 0 1 40
box -113 -50 4688 8286
use pmos331020  pmos331020_2
timestamp 1634181701
transform 1 0 8743 0 1 12
box -113 -50 4688 8286
<< labels >>
flabel locali 4765 8043 4765 8043 0 FreeSans 800 0 0 0 d
flabel locali 8512 8064 8512 8064 0 FreeSans 800 0 0 0 s
flabel locali 4522 5926 4522 5926 0 FreeSans 800 0 0 0 sub
flabel poly 6530 8136 6530 8136 0 FreeSans 800 0 0 0 g
<< end >>
