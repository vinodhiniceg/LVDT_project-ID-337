magic
tech sky130A
magscale 1 2
timestamp 1634273660
<< nwell >>
rect -218 22778 3696 23614
rect -218 22726 3700 22778
rect -216 19150 3700 22726
rect -216 18976 2396 19150
rect 2526 18976 3700 19150
rect -216 -22 3700 18976
<< poly >>
rect 1032 23422 2962 23520
rect 902 22568 980 22782
rect 1350 22568 1428 22782
rect 2098 22560 2170 22792
rect 2650 22554 2722 22786
rect 906 18792 1012 19098
rect 1314 18792 1420 19098
rect 2022 18798 2128 19104
rect 2624 18792 2730 19098
rect 926 15018 1032 15324
rect 1360 15014 1466 15320
rect 2080 15012 2186 15318
rect 2664 15012 2770 15318
rect 896 11260 1002 11566
rect 1270 11250 1376 11556
rect 2042 11248 2148 11554
rect 2660 11254 2766 11560
rect 910 7470 1006 7794
rect 1378 7472 1474 7796
rect 1988 7468 2084 7792
rect 2678 7466 2774 7790
rect 934 3698 1030 4022
rect 1362 3694 1458 4018
rect 2038 3690 2134 4014
rect 2700 3690 2796 4014
<< locali >>
rect 1820 23358 1918 23366
rect 3142 23358 3218 23362
rect 516 23354 3218 23358
rect 512 23256 3218 23354
rect 512 23018 566 23256
rect 1820 23138 1918 23256
rect 3142 23112 3218 23256
rect 484 22384 576 23018
rect 1156 22938 1234 23074
rect 2474 23044 2552 23064
rect 2450 23030 2552 23044
rect 2450 22940 2556 23030
rect 2336 22938 2556 22940
rect 1156 22862 2556 22938
rect 1156 22860 2352 22862
rect 1168 22858 2352 22860
rect 2476 22854 2556 22862
rect 472 18588 538 19450
rect 2446 19150 2504 19216
rect 464 14844 546 15710
rect 476 11074 536 11986
rect 476 7236 552 8304
rect 484 3448 560 4516
<< metal1 >>
rect 2428 22680 2554 23072
rect 2426 22648 2554 22680
rect 2426 22614 2526 22648
rect 2428 22220 2526 22614
rect 2454 22218 2526 22220
rect 2450 18438 2534 19384
rect 2426 14626 2550 15624
rect 2448 10856 2524 11924
rect 2448 7086 2524 8154
rect 2448 3306 2524 4374
use pmos3345  pmos3345_0 ~/layout test
timestamp 1634272161
transform 1 0 450 0 1 192
box -450 -192 2936 3588
use pmos3345  pmos3345_1
timestamp 1634272161
transform 1 0 446 0 1 3964
box -450 -192 2936 3588
use pmos3345  pmos3345_2
timestamp 1634272161
transform 1 0 446 0 1 7740
box -450 -192 2936 3588
use pmos3345  pmos3345_3
timestamp 1634272161
transform 1 0 446 0 1 11504
box -450 -192 2936 3588
use pmos3345  pmos3345_4
timestamp 1634272161
transform 1 0 446 0 1 15274
box -450 -192 2936 3588
use pmos3345  pmos3345_5
timestamp 1634272161
transform 1 0 450 0 1 19050
box -450 -192 2936 3588
use sky130_fd_pr__pfet_g5v0d10v5_6STA4Z  sky130_fd_pr__pfet_g5v0d10v5_6STA4Z_0 ~/layout test
timestamp 1634272774
transform 1 0 1859 0 1 23102
box -1411 -366 1411 366
<< end >>
