magic
tech sky130A
timestamp 1634301196
<< pwell >>
rect 12764 21313 42868 21326
rect 12764 20657 42883 21313
rect 12788 20391 42883 20657
rect 12788 20237 32589 20391
rect 32639 20237 32734 20391
rect 32833 20237 42883 20391
rect 12788 17445 42883 20237
rect 12788 17429 30994 17445
rect 12788 17398 24554 17429
rect 24598 17414 30994 17429
rect 31156 17414 42883 17445
rect 24598 17398 42883 17414
rect 12788 8897 42883 17398
rect 12788 8839 20496 8897
rect 22649 8839 42883 8897
rect 12788 3042 42883 8839
rect 12788 2863 23728 3042
rect 25965 2863 42883 3042
rect 12788 -748 42883 2863
rect 12788 -1375 42910 -748
rect 42543 -1390 42883 -1375
<< mvpsubdiff >>
rect 12764 21313 42868 21326
rect 12764 20657 42883 21313
rect 12788 -748 13615 20657
rect 42543 19586 42883 20657
rect 42529 19496 42883 19586
rect 42529 18712 42550 19496
rect 42682 18712 42883 19496
rect 42529 18643 42883 18712
rect 42543 16527 42883 18643
rect 42543 15833 42606 16527
rect 42710 15833 42883 16527
rect 42543 13558 42883 15833
rect 42543 12823 42585 13558
rect 42751 12823 42883 13558
rect 42543 10735 42883 12823
rect 42543 9958 42571 10735
rect 42696 9958 42883 10735
rect 42543 7842 42883 9958
rect 42543 7100 42613 7842
rect 42710 7100 42883 7842
rect 42543 4881 42883 7100
rect 42543 4194 42613 4881
rect 42731 4194 42883 4881
rect 42543 1967 42883 4194
rect 42543 1280 42606 1967
rect 42689 1280 42883 1967
rect 42543 -748 42883 1280
rect 12788 -1375 42910 -748
rect 42543 -1390 42883 -1375
<< mvpsubdiffcont >>
rect 42550 18712 42682 19496
rect 42606 15833 42710 16527
rect 42585 12823 42751 13558
rect 42571 9958 42696 10735
rect 42613 7100 42710 7842
rect 42613 4194 42731 4881
rect 42606 1280 42689 1967
<< poly >>
rect 24718 20555 31683 20609
rect 34223 20578 41188 20631
rect 24718 20544 31785 20555
rect 34223 20549 37539 20578
rect 15843 20478 21213 20521
rect 15843 20459 18289 20478
rect 15526 20413 18289 20459
rect 18384 20459 21213 20478
rect 24502 20461 31785 20544
rect 18384 20413 21495 20459
rect 15526 20410 21495 20413
rect 15526 20340 16044 20410
rect 18079 20338 18597 20410
rect 20977 20340 21495 20410
rect 24502 20335 25042 20461
rect 27817 20335 28357 20461
rect 31245 20346 31785 20461
rect 34009 20483 37539 20549
rect 34009 20340 34549 20483
rect 37371 20446 37539 20483
rect 37751 20571 41188 20578
rect 37751 20483 41499 20571
rect 37751 20446 37911 20483
rect 37371 20359 37911 20446
rect 40959 20362 41499 20483
rect 14008 17419 14091 17618
rect 14455 17423 14538 17622
rect 14970 17421 15053 17620
rect 15487 17427 15570 17626
rect 16004 17417 16087 17616
rect 17231 17587 19556 17619
rect 18340 17427 18504 17587
rect 20493 17572 22621 17623
rect 21905 17434 21983 17572
rect 23771 17523 26010 17617
rect 24562 17429 24711 17523
rect 27030 17515 29179 17624
rect 30272 17526 32517 17628
rect 33506 17527 35751 17627
rect 24598 17407 24711 17429
rect 27801 17424 27950 17515
rect 30999 17445 31148 17526
rect 34277 17424 34426 17527
rect 36816 17501 39045 17638
rect 40046 17562 42343 17644
rect 38003 17447 38152 17501
rect 40634 17432 40747 17562
rect 14042 14512 14125 14711
rect 14459 14512 14542 14711
rect 15008 14508 15091 14707
rect 15508 14510 15591 14709
rect 16040 14512 16123 14711
rect 17238 14668 19544 14712
rect 18327 14514 18513 14668
rect 20494 14645 22765 14715
rect 22142 14517 22224 14645
rect 23742 14604 25982 14708
rect 27020 14620 29260 14716
rect 30266 14627 32510 14720
rect 24373 14484 24522 14604
rect 27772 14513 27921 14620
rect 30987 14513 31136 14627
rect 33509 14623 35751 14719
rect 36788 14635 39038 14730
rect 34306 14507 34455 14623
rect 37871 14518 38020 14635
rect 40063 14615 42296 14737
rect 40618 14517 40731 14615
rect 14042 11597 14125 11796
rect 14404 11593 14487 11792
rect 14927 11595 15010 11794
rect 15442 11595 15525 11794
rect 16014 11595 16097 11794
rect 17234 11758 19539 11795
rect 18464 11596 18501 11758
rect 20493 11718 22707 11798
rect 21733 11596 21844 11718
rect 23829 11681 25978 11791
rect 27021 11694 29261 11800
rect 30267 11699 32512 11802
rect 33507 11717 35759 11801
rect 36788 11718 39038 11813
rect 24379 11584 24528 11681
rect 27909 11589 28058 11694
rect 31194 11569 31375 11699
rect 34448 11584 34561 11717
rect 37417 11579 37530 11718
rect 40085 11708 42322 11820
rect 40575 11595 40688 11708
rect 14063 8665 14171 8877
rect 14447 8663 14555 8875
rect 14970 8661 15078 8873
rect 15489 8663 15597 8875
rect 15959 8663 16067 8875
rect 17238 8853 19581 8877
rect 18288 8647 18378 8853
rect 20496 8771 22627 8881
rect 21704 8662 21776 8771
rect 23763 8761 25913 8874
rect 26963 8779 29202 8879
rect 30238 8780 32483 8883
rect 33505 8787 35755 8885
rect 36739 8801 38989 8896
rect 24320 8655 24423 8761
rect 27977 8657 28080 8779
rect 31256 8660 31359 8780
rect 34464 8647 34577 8787
rect 37428 8663 37541 8801
rect 40043 8789 42280 8901
rect 40591 8685 40704 8789
rect 14048 5736 14156 5948
rect 14432 5731 14540 5943
rect 14953 5731 15061 5943
rect 15478 5736 15586 5948
rect 16038 5734 16146 5946
rect 17243 5898 19521 5945
rect 18301 5729 18391 5898
rect 20514 5867 22748 5950
rect 21621 5731 21705 5867
rect 23740 5828 25890 5941
rect 27053 5842 29198 5950
rect 30267 5846 32513 5951
rect 24285 5709 24388 5828
rect 28014 5728 28117 5842
rect 31235 5738 31338 5846
rect 33501 5844 35750 5952
rect 36815 5865 39053 5963
rect 34469 5736 34582 5844
rect 37761 5742 37874 5865
rect 40057 5859 42294 5971
rect 40570 5742 40683 5859
rect 14070 2772 14203 3020
rect 14440 2772 14573 3020
rect 15004 2774 15137 3022
rect 15463 2770 15596 3018
rect 16046 2768 16179 3016
rect 17215 2974 19491 3017
rect 18335 2778 18425 2974
rect 20510 2960 22788 3021
rect 21566 2783 21671 2960
rect 23796 2878 26025 3012
rect 27009 2927 29156 3020
rect 24333 2764 24436 2878
rect 28041 2775 28144 2927
rect 30301 2910 32547 3024
rect 33525 2911 35773 3023
rect 36812 2934 39050 3036
rect 40088 2944 42324 3042
rect 31227 2777 31330 2910
rect 34007 2767 34120 2911
rect 37315 2788 37428 2934
rect 40527 2783 40640 2944
<< polycont >>
rect 18289 20413 18384 20478
rect 37539 20446 37751 20578
<< locali >>
rect 37491 20578 37799 20612
rect 18272 20478 18409 20497
rect 13719 2614 13787 20423
rect 18272 20413 18289 20478
rect 18384 20413 18409 20478
rect 18272 20393 18409 20413
rect 16384 20291 16452 20305
rect 15850 20168 17088 20291
rect 18303 20248 18360 20393
rect 19076 20248 20477 20286
rect 22891 20280 22933 20285
rect 19053 20222 20477 20248
rect 16384 2496 16452 20168
rect 16982 2454 17050 20168
rect 19637 20121 19708 20222
rect 19635 20113 19708 20121
rect 19635 20096 19701 20113
rect 19648 2530 19701 20096
rect 20234 3230 20278 20222
rect 22355 20213 22933 20280
rect 22885 20103 22933 20213
rect 23235 20147 23461 20427
rect 28866 20287 28869 20296
rect 30070 20287 30200 20296
rect 23506 20218 23518 20279
rect 25594 20207 26884 20276
rect 28849 20191 30304 20287
rect 31995 20191 32160 20282
rect 32616 20165 32788 20549
rect 37491 20446 37539 20578
rect 37751 20446 37799 20578
rect 37491 20417 37799 20446
rect 33198 20191 33329 20282
rect 35355 20230 36714 20279
rect 37585 20248 37683 20417
rect 42438 20300 42487 20338
rect 38653 20241 40012 20290
rect 22885 14975 22932 20103
rect 32643 19975 32725 20165
rect 35892 19887 35957 20230
rect 39179 19897 39244 20241
rect 41912 20209 42487 20300
rect 42438 20042 42487 20209
rect 42529 19496 42731 19586
rect 42529 18712 42550 19496
rect 42682 18712 42731 19496
rect 42529 18643 42731 18712
rect 23477 17264 23543 17968
rect 26116 17171 26182 17875
rect 26749 17305 26815 18009
rect 29986 17865 30047 17969
rect 29389 17153 29455 17857
rect 29986 17841 30052 17865
rect 29989 17173 30052 17841
rect 32648 17166 32711 17858
rect 33245 17216 33308 17908
rect 35885 17174 35948 17866
rect 36538 17208 36604 17912
rect 39189 17209 39237 17878
rect 39795 17242 39843 17911
rect 42435 17176 42483 17845
rect 42564 16527 42765 16652
rect 42564 15833 42606 16527
rect 42710 15833 42765 16527
rect 42564 15688 42765 15833
rect 22885 14271 22954 14975
rect 23484 14364 23550 15068
rect 22885 12042 22932 14271
rect 26138 14230 26204 14934
rect 26738 14383 26804 15087
rect 29378 14226 29444 14930
rect 29989 14304 30052 14996
rect 32641 14276 32704 14968
rect 33245 14269 33308 14961
rect 35885 14234 35948 14926
rect 36526 14301 36592 15005
rect 39185 14292 39233 14961
rect 39770 14939 39836 15013
rect 39770 14309 39851 14939
rect 42439 14292 42487 14961
rect 42557 13558 42779 13655
rect 42557 12823 42585 13558
rect 42751 12823 42779 13558
rect 42557 12677 42779 12823
rect 22884 11338 22950 12042
rect 23469 11442 23535 12146
rect 26134 11345 26200 12049
rect 26746 11446 26812 12150
rect 20234 2526 20300 3230
rect 22885 3223 22932 11338
rect 29393 11330 29456 12022
rect 29989 11386 30052 12078
rect 32641 11295 32704 11987
rect 33245 11336 33308 12028
rect 35885 11350 35948 12042
rect 36534 11453 36600 12157
rect 39182 11361 39230 12030
rect 39803 11494 39851 12163
rect 42442 11383 42490 12052
rect 42550 10735 42731 10867
rect 42550 9958 42571 10735
rect 42696 9958 42731 10735
rect 42550 9819 42731 9958
rect 23469 8456 23535 9177
rect 26108 8408 26174 9112
rect 26727 8535 26793 9239
rect 29386 8397 29449 9089
rect 29997 8503 30060 9195
rect 32641 8397 32704 9089
rect 33238 8472 33301 9164
rect 35885 8417 35948 9109
rect 36538 8453 36604 9157
rect 39193 8426 39241 9095
rect 39776 8453 39839 9145
rect 42446 8448 42494 9117
rect 42578 7842 42765 7953
rect 42578 7100 42613 7842
rect 42710 7100 42765 7842
rect 42578 6961 42765 7100
rect 23484 5571 23550 6275
rect 26138 5486 26204 6190
rect 26749 5594 26815 6298
rect 29386 5437 29449 6129
rect 29989 5542 30052 6234
rect 32648 5458 32711 6150
rect 33252 5546 33315 6238
rect 35892 5434 35955 6126
rect 36528 5556 36591 6248
rect 39179 5584 39242 6276
rect 39783 5598 39846 6290
rect 42455 5514 42518 6206
rect 42585 4881 42765 4957
rect 42585 4194 42613 4881
rect 42731 4194 42765 4881
rect 42585 4111 42765 4194
rect 23491 3301 23526 3318
rect 26751 3305 26798 3360
rect 39790 3337 39852 3354
rect 22885 2527 22954 3223
rect 23491 2597 23557 3301
rect 22888 2519 22954 2527
rect 26119 2515 26185 3219
rect 26746 2601 26812 3305
rect 29393 2519 29456 3211
rect 29997 2589 30060 3281
rect 32655 2547 32718 3239
rect 33238 2613 33301 3305
rect 35892 2473 35955 3165
rect 36535 2617 36598 3309
rect 39200 2505 39263 3197
rect 39790 2645 39853 3337
rect 42448 2526 42511 3218
rect 42564 1967 42738 2016
rect 42564 1280 42606 1967
rect 42689 1280 42738 1967
rect 42564 1197 42738 1280
rect 26015 90 27526 192
rect 29277 95 30775 224
rect 35941 131 41124 234
<< viali >>
rect 18301 20433 18372 20464
rect 37575 20470 37697 20554
rect 42550 18712 42682 19496
rect 42606 15833 42710 16527
rect 42585 12823 42751 13558
rect 42571 9958 42696 10735
rect 42613 7100 42710 7842
rect 42613 4194 42731 4881
rect 42606 1280 42689 1967
<< metal1 >>
rect 37491 20554 37799 20612
rect 18272 20464 18409 20497
rect 18272 20433 18301 20464
rect 18372 20433 18409 20464
rect 18272 20393 18409 20433
rect 37491 20470 37575 20554
rect 37697 20470 37799 20554
rect 37491 20417 37799 20470
rect 42529 19496 42731 19586
rect 42529 18712 42550 19496
rect 42682 18712 42731 19496
rect 42529 18643 42731 18712
rect 42564 16527 42765 16652
rect 42564 15833 42606 16527
rect 42710 15833 42765 16527
rect 42564 15688 42765 15833
rect 42557 13558 42779 13655
rect 42557 12823 42585 13558
rect 42751 12823 42779 13558
rect 42557 12677 42779 12823
rect 42550 10735 42731 10867
rect 42550 9958 42571 10735
rect 42696 9958 42731 10735
rect 42550 9819 42731 9958
rect 42578 7842 42765 7953
rect 42578 7100 42613 7842
rect 42710 7100 42765 7842
rect 42578 6961 42765 7100
rect 42585 4881 42765 4957
rect 42585 4194 42613 4881
rect 42731 4194 42765 4881
rect 42585 4111 42765 4194
rect 42564 1967 42738 2016
rect 42564 1280 42606 1967
rect 42689 1280 42738 1967
rect 42564 1197 42738 1280
use nmos55535  nmos55535_4
timestamp 1634301196
transform 1 0 13375 0 1 -14
box -14 0 3221 20454
use nmos55535  nmos55535_5
timestamp 1634301196
transform 1 0 16632 0 1 -10
box -14 0 3221 20454
use nmos55535  nmos55535_6
timestamp 1634301196
transform 1 0 19885 0 1 -6
box -14 0 3221 20454
use nmos55535  nmos55535_7
timestamp 1634301196
transform 1 0 23130 0 1 -14
box -14 0 3221 20454
use nmos55535  nmos55535_8
timestamp 1634301196
transform 1 0 26391 0 1 -6
box -14 0 3221 20454
use nmos55535  nmos55535_0
timestamp 1634301196
transform 1 0 29646 0 1 -3
box -14 0 3221 20454
use nmos55535  nmos55535_1
timestamp 1634301196
transform 1 0 32891 0 1 -3
box -14 0 3221 20454
use nmos55535  nmos55535_2
timestamp 1634301196
transform 1 0 36185 0 1 8
box -14 0 3221 20454
use nmos55535  nmos55535_3
timestamp 1634301196
transform 1 0 39442 0 1 15
box -14 0 3221 20454
<< labels >>
flabel poly 28014 20518 28014 20518 0 FreeSans 1600 0 0 0 g
flabel locali 32680 20414 32680 20414 0 FreeSans 1600 0 0 0 S
flabel locali 23293 20251 23293 20251 0 FreeSans 1600 0 0 0 D
<< end >>
