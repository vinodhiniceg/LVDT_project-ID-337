magic
tech sky130A
magscale 1 2
timestamp 1634206384
<< error_p >>
rect -2216 -2600 -2156 2600
rect -2136 -2600 -2076 2600
rect 2076 -2600 2136 2600
rect 2156 -2600 2216 2600
<< metal3 >>
rect -6428 2572 -2156 2600
rect -6428 -2572 -2240 2572
rect -2176 -2572 -2156 2572
rect -6428 -2600 -2156 -2572
rect -2136 2572 2136 2600
rect -2136 -2572 2052 2572
rect 2116 -2572 2136 2572
rect -2136 -2600 2136 -2572
rect 2156 2572 6428 2600
rect 2156 -2572 6344 2572
rect 6408 -2572 6428 2572
rect 2156 -2600 6428 -2572
<< via3 >>
rect -2240 -2572 -2176 2572
rect 2052 -2572 2116 2572
rect 6344 -2572 6408 2572
<< mimcap >>
rect -6328 2460 -2328 2500
rect -6328 -2460 -4916 2460
rect -3740 -2460 -2328 2460
rect -6328 -2500 -2328 -2460
rect -2036 2460 1964 2500
rect -2036 -2460 -624 2460
rect 552 -2460 1964 2460
rect -2036 -2500 1964 -2460
rect 2256 2460 6256 2500
rect 2256 -2460 3668 2460
rect 4844 -2460 6256 2460
rect 2256 -2500 6256 -2460
<< mimcapcontact >>
rect -4916 -2460 -3740 2460
rect -624 -2460 552 2460
rect 3668 -2460 4844 2460
<< metal4 >>
rect -2256 2572 -2160 2588
rect -4917 2460 -3739 2461
rect -4917 -2460 -4916 2460
rect -3740 -2460 -3739 2460
rect -4917 -2461 -3739 -2460
rect -2256 -2572 -2240 2572
rect -2176 -2572 -2160 2572
rect 2036 2572 2132 2588
rect -625 2460 553 2461
rect -625 -2460 -624 2460
rect 552 -2460 553 2460
rect -625 -2461 553 -2460
rect -2256 -2588 -2160 -2572
rect 2036 -2572 2052 2572
rect 2116 -2572 2132 2572
rect 6328 2572 6424 2588
rect 3667 2460 4845 2461
rect 3667 -2460 3668 2460
rect 4844 -2460 4845 2460
rect 3667 -2461 4845 -2460
rect 2036 -2588 2132 -2572
rect 6328 -2572 6344 2572
rect 6408 -2572 6424 2572
rect 6328 -2588 6424 -2572
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX 2156 -2600 6356 2600
string parameters w 20.00 l 25.00 val 1.017k carea 2.00 cperi 0.19 nx 3 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 30
string library sky130
<< end >>
