* NGSPICE file created from colpitts4_flat.ext - technology: sky130A


* Top level circuit colpitts4_flat

X0 vout2.t1 vout1.t2 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+06u l=3e+06u
X1 bot bot bot bot sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+06u l=3e+06u M=138
X2 vout2 vout1 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+06u l=3e+06u M=199
X3 bot bot bot bot sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=5e+06u M=1450
X4 vdda vdda vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+06u l=3e+06u M=1016
X5 vcap.t0 vin1 vout.t0 bot sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=5e+06u
X6 bot vout1.t3 vout2.t0 bot sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+06u l=3e+06u
X7 vout vin1 vcap bot sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=5e+06u M=524
X8 vout1.t0 vout.t1 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+06u l=3e+06u
X9 vout1 vout vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+06u l=3e+06u M=183
X10 bot vin2 vcap.t1 bot sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=5e+06u
X11 vout3.t1 vout2.t2 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+06u l=3e+06u
X12 vcap vin2 bot bot sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=5e+06u M=199
X13 vdda vout2 vout3 vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+06u l=3e+06u M=123
X14 vout3.t0 vout2.t3 bot bot sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+06u l=3e+06u
X15 vout2 vout1 bot bot sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+06u l=3e+06u M=24
X16 bot vout.t2 vout1.t1 bot sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+06u l=3e+06u
X17 vout1 vout bot bot sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+06u l=3e+06u M=19
X18 vout3 vout2 bot bot sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+06u l=3e+06u M=23
X19 a_85326_53811# a_83611_53805# a_85147_53811# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X20 vout3.t2 bot sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2.5e+07u
X21 a_84193_53900# a_83611_53805# a_83724_53900# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X22 vout2.t4 bot sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2.5e+07u
X23 a_85659_53375# vdda bot bot sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X24 a_83611_53805# a_83302_53375.t2 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X25 vdda clkin a_83302_53375.t1 vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X26 vout1.t4 bot sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2.5e+07u
X27 a_84391_53774# a_84193_53900# bot bot sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X28 vdda a_85147_53811# a_85921_53475# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X29 a_84363_53441# a_83611_53805# a_84193_53900# bot sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X30 bot a_85368_53685# a_85361_53375# bot sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X31 dfout a_85921_53475# bot bot sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X32 a_84391_53774# a_84193_53900# vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X33 bot a_85147_53811# a_85921_53475# bot sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X34 vdda vdda a_83724_53900# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X35 a_84349_53900# a_83302_53375.t3 a_84193_53900# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X36 a_84193_53900# vdda vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X37 vdda a_85368_53685# a_85326_53811# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X38 a_83611_53805# a_83302_53375.t4 bot bot sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X39 vout3 bot sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2.5e+07u
X40 bot clkin a_83302_53375.t0 bot sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X41 a_83909_53441# vdda bot bot sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X42 vdda a_84391_53774# a_84349_53900# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X43 a_85147_53811# a_83302_53375.t5 a_84391_53774# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X44 vout2 bot sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2.5e+07u
X45 a_83724_53900# vout3.t3 a_83909_53441# bot sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X46 vout1 bot sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2.5e+07u
X47 vout2 bot sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2.5e+07u
X48 bot vdda a_84505_53441# bot sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X49 a_83724_53900# vout3.t4 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X50 vdda a_85147_53811# a_85368_53685# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X51 a_85368_53685# vdda vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X52 a_85361_53375# a_83302_53375.t6 a_85147_53811# bot sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X53 a_85368_53685# a_85147_53811# a_85659_53375# bot sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X54 vout1 bot sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2.5e+07u
X55 a_84193_53900# a_83302_53375.t7 a_83724_53900# bot sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X56 a_85147_53811# a_83611_53805# a_84391_53774# bot sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X57 vout1 bot sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2.5e+07u
X58 vout1 bot sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2.5e+07u
X59 dfout a_85921_53475# vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X60 a_84505_53441# a_84391_53774# a_84363_53441# bot sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
R0 vout1.n0 vout1.t1 1554.43
R1 vout1 vout1.n279 1537.99
R2 vout1.n280 vout1 703.239
R3 vout1.n246 vout1.n245 381.257
R4 vout1.n159 vout1.n153 368.573
R5 vout1.n153 vout1.n95 368.573
R6 vout1.n248 vout1.n247 368.573
R7 vout1.n247 vout1.n246 363.643
R8 vout1.n248 vout1.n43 325.302
R9 vout1.n240 vout1.n239 317.928
R10 vout1.n159 vout1.n158 305.036
R11 vout1.n239 vout1.n233 271.976
R12 vout1.n280 vout1.t0 265.444
R13 vout1.n223 vout1.n222 257.825
R14 vout1.n212 vout1.n95 237.666
R15 vout1.n222 vout1.n221 235.213
R16 vout1.n89 vout1.n54 223.973
R17 vout1.n254 vout1.n38 159.889
R18 vout1.n170 vout1.n169 153.573
R19 vout1.n171 vout1.n119 153.566
R20 vout1.n107 vout1.n106 153.547
R21 vout1.n101 vout1.n100 153.516
R22 vout1.n148 vout1.n141 153.482
R23 vout1.n164 vout1.n163 152.655
R24 vout1.n207 vout1.n206 152.572
R25 vout1.n201 vout1.n200 152.572
R26 vout1.n33 vout1.n21 152.45
R27 vout1.n27 vout1.n26 152.394
R28 vout1.n260 vout1.n259 152.34
R29 vout1.n60 vout1.n59 152.321
R30 vout1.n44 vout1.n38 152.125
R31 vout1.n16 vout1.n10 151.673
R32 vout1.n39 vout1.n32 151.635
R33 vout1.n54 vout1.n53 151.612
R34 vout1.n266 vout1.n265 151.533
R35 vout1.n267 vout1.n4 151.363
R36 vout1.n254 vout1.n253 151.312
R37 vout1.n76 vout1.n75 151.061
R38 vout1.n177 vout1.n113 149.481
R39 vout1.n171 vout1.n107 148.934
R40 vout1.n132 vout1.n113 147.855
R41 vout1.n177 vout1.n176 147.764
R42 vout1.n188 vout1.n187 147.623
R43 vout1.n164 vout1.n147 147.017
R44 vout1.n195 vout1.n194 146.994
R45 vout1.n142 vout1.n131 146.873
R46 vout1.n154 vout1.n147 146.862
R47 vout1.n84 vout1.n83 145.868
R48 vout1.n266 vout1.n10 145.648
R49 vout1.n188 vout1.n177 145.647
R50 vout1.n90 vout1.n89 145.564
R51 vout1.n78 vout1.n77 144.95
R52 vout1.n260 vout1.n21 144.004
R53 vout1.n126 vout1.n125 141.082
R54 vout1.n141 vout1.n101 137.431
R55 vout1.n60 vout1.n21 135.788
R56 vout1.n171 vout1.n170 135.24
R57 vout1.n77 vout1.n76 134.398
R58 vout1.n54 vout1.n38 124.834
R59 vout1.n76 vout1.n10 124.833
R60 vout1.n164 vout1.n141 120.452
R61 vout1.n83 vout1.n60 117.987
R62 vout1.n125 vout1.n113 105.335
R63 vout1.n200 vout1.n107 105.116
R64 vout1.n206 vout1.n101 102.377
R65 vout1.n242 vout1.n212 102.349
R66 vout1.n170 vout1.n131 100.305
R67 vout1.n260 vout1.n26 99.639
R68 vout1.n267 vout1.n266 98.542
R69 vout1.n194 vout1.n188 95.256
R70 vout1.n254 vout1.n32 85.397
R71 vout1.n245 vout1.n244 84.164
R72 vout1.n225 vout1.n224 48.2
R73 vout1.n226 vout1.n225 48.2
R74 vout1.n227 vout1.n226 48.2
R75 vout1.n228 vout1.n227 48.2
R76 vout1.n218 vout1.t3 48.2
R77 vout1.n219 vout1.n218 48.2
R78 vout1.n220 vout1.n219 48.2
R79 vout1.n221 vout1.n220 48.2
R80 vout1.n214 vout1.n213 48.2
R81 vout1.n215 vout1.n214 48.2
R82 vout1.n216 vout1.n215 48.2
R83 vout1.n217 vout1.n216 48.2
R84 vout1.n230 vout1.n229 48.2
R85 vout1.n231 vout1.n230 48.2
R86 vout1.n232 vout1.n231 48.2
R87 vout1.n233 vout1.n232 48.2
R88 vout1.n235 vout1.n234 48.2
R89 vout1.n236 vout1.n235 48.2
R90 vout1.n237 vout1.n236 48.2
R91 vout1.n238 vout1.n237 48.2
R92 vout1.n152 vout1.n151 48.2
R93 vout1.n151 vout1.n150 48.2
R94 vout1.n150 vout1.n149 48.2
R95 vout1.n149 vout1.n148 48.2
R96 vout1.n121 vout1.n120 48.2
R97 vout1.n122 vout1.n121 48.2
R98 vout1.n123 vout1.n122 48.2
R99 vout1.n124 vout1.n123 48.2
R100 vout1.n146 vout1.n145 48.2
R101 vout1.n145 vout1.n144 48.2
R102 vout1.n144 vout1.n143 48.2
R103 vout1.n143 vout1.n142 48.2
R104 vout1.n130 vout1.n129 48.2
R105 vout1.n129 vout1.n128 48.2
R106 vout1.n128 vout1.n127 48.2
R107 vout1.n127 vout1.n126 48.2
R108 vout1.n109 vout1.n108 48.2
R109 vout1.n110 vout1.n109 48.2
R110 vout1.n111 vout1.n110 48.2
R111 vout1.n112 vout1.n111 48.2
R112 vout1.n136 vout1.n135 48.2
R113 vout1.n135 vout1.n134 48.2
R114 vout1.n134 vout1.n133 48.2
R115 vout1.n133 vout1.n132 48.2
R116 vout1.n115 vout1.n114 48.2
R117 vout1.n116 vout1.n115 48.2
R118 vout1.n117 vout1.n116 48.2
R119 vout1.n118 vout1.n117 48.2
R120 vout1.n173 vout1.n172 48.2
R121 vout1.n174 vout1.n173 48.2
R122 vout1.n175 vout1.n174 48.2
R123 vout1.n176 vout1.n175 48.2
R124 vout1.n179 vout1.n178 48.2
R125 vout1.n180 vout1.n179 48.2
R126 vout1.n181 vout1.n180 48.2
R127 vout1.n182 vout1.n181 48.2
R128 vout1.n184 vout1.n183 48.2
R129 vout1.n185 vout1.n184 48.2
R130 vout1.n186 vout1.n185 48.2
R131 vout1.n187 vout1.n186 48.2
R132 vout1.n190 vout1.n189 48.2
R133 vout1.n191 vout1.n190 48.2
R134 vout1.n192 vout1.n191 48.2
R135 vout1.n193 vout1.n192 48.2
R136 vout1.n196 vout1.n195 48.2
R137 vout1.n197 vout1.n196 48.2
R138 vout1.n198 vout1.n197 48.2
R139 vout1.n199 vout1.n198 48.2
R140 vout1.n211 vout1.n210 48.2
R141 vout1.n210 vout1.n209 48.2
R142 vout1.n209 vout1.n208 48.2
R143 vout1.n208 vout1.n207 48.2
R144 vout1.n205 vout1.n204 48.2
R145 vout1.n204 vout1.n203 48.2
R146 vout1.n203 vout1.n202 48.2
R147 vout1.n202 vout1.n201 48.2
R148 vout1.n106 vout1.n105 48.2
R149 vout1.n105 vout1.n104 48.2
R150 vout1.n104 vout1.n103 48.2
R151 vout1.n103 vout1.n102 48.2
R152 vout1.n97 vout1.n96 48.2
R153 vout1.n98 vout1.n97 48.2
R154 vout1.n99 vout1.n98 48.2
R155 vout1.n100 vout1.n99 48.2
R156 vout1.n140 vout1.n139 48.2
R157 vout1.n139 vout1.n138 48.2
R158 vout1.n138 vout1.n137 48.2
R159 vout1.n137 vout1.n119 48.2
R160 vout1.n169 vout1.n168 48.2
R161 vout1.n168 vout1.n167 48.2
R162 vout1.n167 vout1.n166 48.2
R163 vout1.n166 vout1.n165 48.2
R164 vout1.n161 vout1.n160 48.2
R165 vout1.t2 vout1.n161 48.2
R166 vout1.n162 vout1.t2 48.2
R167 vout1.n163 vout1.n162 48.2
R168 vout1.n155 vout1.n154 48.2
R169 vout1.n156 vout1.n155 48.2
R170 vout1.n157 vout1.n156 48.2
R171 vout1.n158 vout1.n157 48.2
R172 vout1.n48 vout1.n47 48.2
R173 vout1.n47 vout1.n46 48.2
R174 vout1.n46 vout1.n45 48.2
R175 vout1.n45 vout1.n44 48.2
R176 vout1.n62 vout1.n61 48.2
R177 vout1.n63 vout1.n62 48.2
R178 vout1.n64 vout1.n63 48.2
R179 vout1.n65 vout1.n64 48.2
R180 vout1.n88 vout1.n87 48.2
R181 vout1.n87 vout1.n86 48.2
R182 vout1.n86 vout1.n85 48.2
R183 vout1.n85 vout1.n84 48.2
R184 vout1.n82 vout1.n81 48.2
R185 vout1.n81 vout1.n80 48.2
R186 vout1.n80 vout1.n79 48.2
R187 vout1.n79 vout1.n78 48.2
R188 vout1.n67 vout1.n66 48.2
R189 vout1.n68 vout1.n67 48.2
R190 vout1.n69 vout1.n68 48.2
R191 vout1.n70 vout1.n69 48.2
R192 vout1.n72 vout1.n71 48.2
R193 vout1.n73 vout1.n72 48.2
R194 vout1.n74 vout1.n73 48.2
R195 vout1.n75 vout1.n74 48.2
R196 vout1.n6 vout1.n5 48.2
R197 vout1.n7 vout1.n6 48.2
R198 vout1.n8 vout1.n7 48.2
R199 vout1.n9 vout1.n8 48.2
R200 vout1.n20 vout1.n19 48.2
R201 vout1.n19 vout1.n18 48.2
R202 vout1.n18 vout1.n17 48.2
R203 vout1.n17 vout1.n16 48.2
R204 vout1.n12 vout1.n11 48.2
R205 vout1.n13 vout1.n12 48.2
R206 vout1.n14 vout1.n13 48.2
R207 vout1.n15 vout1.n14 48.2
R208 vout1.n265 vout1.n264 48.2
R209 vout1.n264 vout1.n263 48.2
R210 vout1.n263 vout1.n262 48.2
R211 vout1.n262 vout1.n261 48.2
R212 vout1.n259 vout1.n258 48.2
R213 vout1.n258 vout1.n257 48.2
R214 vout1.n257 vout1.n256 48.2
R215 vout1.n256 vout1.n255 48.2
R216 vout1.n250 vout1.n249 48.2
R217 vout1.n251 vout1.n250 48.2
R218 vout1.n252 vout1.n251 48.2
R219 vout1.n253 vout1.n252 48.2
R220 vout1.n37 vout1.n36 48.2
R221 vout1.n36 vout1.n35 48.2
R222 vout1.n35 vout1.n34 48.2
R223 vout1.n34 vout1.n33 48.2
R224 vout1.n59 vout1.n58 48.2
R225 vout1.n58 vout1.n57 48.2
R226 vout1.n57 vout1.n56 48.2
R227 vout1.n56 vout1.n55 48.2
R228 vout1.n50 vout1.n49 48.2
R229 vout1.n51 vout1.n50 48.2
R230 vout1.n52 vout1.n51 48.2
R231 vout1.n53 vout1.n52 48.2
R232 vout1.n91 vout1.n90 48.2
R233 vout1.n92 vout1.n91 48.2
R234 vout1.n93 vout1.n92 48.2
R235 vout1.n94 vout1.n93 48.2
R236 vout1.n43 vout1.n42 48.2
R237 vout1.n42 vout1.n41 48.2
R238 vout1.n41 vout1.n40 48.2
R239 vout1.n40 vout1.n39 48.2
R240 vout1.n31 vout1.n30 48.2
R241 vout1.n30 vout1.n29 48.2
R242 vout1.n29 vout1.n28 48.2
R243 vout1.n28 vout1.n27 48.2
R244 vout1.n25 vout1.n24 48.2
R245 vout1.n24 vout1.n23 48.2
R246 vout1.n23 vout1.n22 48.2
R247 vout1.n22 vout1.n4 48.2
R248 vout1.n269 vout1.n268 48.2
R249 vout1.n270 vout1.n269 48.2
R250 vout1.n271 vout1.n270 48.2
R251 vout1.n272 vout1.n271 48.2
R252 vout1.n279 vout1.n0 38.407
R253 vout1.n125 vout1.n124 31.66
R254 vout1.n77 vout1.n65 31.659
R255 vout1.n147 vout1.n146 31.658
R256 vout1.n89 vout1.n88 31.658
R257 vout1.n131 vout1.n130 31.605
R258 vout1.n83 vout1.n82 31.604
R259 vout1.n273 vout1.n272 29.507
R260 vout1.n240 vout1.n228 24.101
R261 vout1.n222 vout1.n217 24.1
R262 vout1.n239 vout1.n238 24.1
R263 vout1.n153 vout1.n152 24.1
R264 vout1.n113 vout1.n112 24.1
R265 vout1.n170 vout1.n136 24.1
R266 vout1.n177 vout1.n118 24.1
R267 vout1.n172 vout1.n171 24.1
R268 vout1.n188 vout1.n182 24.1
R269 vout1.n183 vout1.n107 24.1
R270 vout1.n194 vout1.n193 24.1
R271 vout1.n200 vout1.n199 24.1
R272 vout1.n212 vout1.n211 24.1
R273 vout1.n206 vout1.n205 24.1
R274 vout1.n102 vout1.n101 24.1
R275 vout1.n96 vout1.n95 24.1
R276 vout1.n141 vout1.n140 24.1
R277 vout1.n165 vout1.n164 24.1
R278 vout1.n160 vout1.n159 24.1
R279 vout1.n247 vout1.n48 24.1
R280 vout1.n76 vout1.n70 24.1
R281 vout1.n71 vout1.n60 24.1
R282 vout1.n10 vout1.n9 24.1
R283 vout1.n21 vout1.n20 24.1
R284 vout1.n266 vout1.n15 24.1
R285 vout1.n261 vout1.n260 24.1
R286 vout1.n255 vout1.n254 24.1
R287 vout1.n249 vout1.n248 24.1
R288 vout1.n38 vout1.n37 24.1
R289 vout1.n55 vout1.n54 24.1
R290 vout1.n246 vout1.n49 24.1
R291 vout1.n245 vout1.n94 24.1
R292 vout1.n32 vout1.n31 24.1
R293 vout1.n26 vout1.n25 24.1
R294 vout1.n268 vout1.n267 24.1
R295 vout1 vout1.n243 16.936
R296 vout1 vout1.n280 15.857
R297 vout1.n0 vout1 15.369
R298 vout1.n244 vout1 14.763
R299 vout1.n244 vout1.n243 10.666
R300 vout1.n242 vout1.n241 9.703
R301 vout1.n241 vout1.n223 7.158
R302 vout1.n279 vout1.n278 2.446
R303 vout1.n223 vout1 1.285
R304 vout1.n277 vout1.t4 0.557
R305 vout1.n274 vout1.n273 0.443
R306 vout1 vout1.n274 0.371
R307 vout1.n241 vout1.n240 0.34
R308 vout1.n243 vout1.n242 0.246
R309 vout1.n278 vout1.n275 0.219
R310 vout1.n278 vout1.n277 0.18
R311 vout1.n273 vout1.n3 0.163
R312 vout1.n274 vout1.n2 0.157
R313 vout1.n275 vout1.n1 0.157
R314 vout1.n277 vout1.n276 0.157
R315 vout1.n275 vout1 0.035
R316 vout2 vout2.t1 1131.96
R317 vout2.n188 vout2 905.362
R318 vout2 vout2.t0 623.923
R319 vout2.n185 vout2.n184 472.435
R320 vout2 vout2.n187 346.183
R321 vout2.n122 vout2 307.132
R322 vout2.n183 vout2.n182 298.282
R323 vout2.n124 vout2.n123 285.127
R324 vout2.n120 vout2.n119 273.61
R325 vout2.n120 vout2.n34 260.13
R326 vout2.n16 vout2.n15 213.521
R327 vout2.n87 vout2.n64 213.472
R328 vout2.n148 vout2.n147 213.146
R329 vout2.n10 vout2.n9 212.536
R330 vout2.n154 vout2.n153 211.221
R331 vout2.n82 vout2.n81 209.659
R332 vout2.n90 vout2.n89 208.583
R333 vout2.n184 vout2 207.793
R334 vout2.n74 vout2.n73 207.463
R335 vout2.n117 vout2.n40 204.444
R336 vout2.n119 vout2.n118 203.761
R337 vout2.n95 vout2.n21 199.205
R338 vout2.n35 vout2.n33 196.871
R339 vout2.n118 vout2.n117 196.473
R340 vout2.n112 vout2.n111 196.214
R341 vout2.n130 vout2.n129 194.849
R342 vout2.n28 vout2.n27 194.708
R343 vout2.n48 vout2.n47 192.937
R344 vout2.n136 vout2.n135 192.895
R345 vout2.n187 vout2 192.394
R346 vout2.n102 vout2.n53 191.785
R347 vout2.n97 vout2.n96 191.725
R348 vout2.n22 vout2.n21 191.691
R349 vout2.n142 vout2.n141 190.12
R350 vout2.n105 vout2.n104 188.993
R351 vout2.n59 vout2.n58 187.08
R352 vout2.n103 vout2.n27 185.584
R353 vout2.n110 vout2.n33 182.44
R354 vout2.n148 vout2.n15 180.344
R355 vout2.n80 vout2.n9 176.678
R356 vout2.n154 vout2.n9 173.01
R357 vout2.n122 vout2.n121 172.114
R358 vout2.n124 vout2.n34 171.836
R359 vout2.n40 vout2.n39 160.595
R360 vout2.n88 vout2.n15 159.388
R361 vout2.n142 vout2.n21 158.864
R362 vout2.n130 vout2.n33 154.673
R363 vout2.n136 vout2.n27 149.958
R364 vout2.n88 vout2.n87 122.191
R365 vout2.n81 vout2.n80 111.713
R366 vout2.n103 vout2.n102 110.664
R367 vout2.n111 vout2.n110 103.853
R368 vout2 vout2.n183 99.128
R369 vout2.n96 vout2.n95 94.947
R370 vout2 vout2.n188 65.344
R371 vout2.n42 vout2.n40 59.202
R372 vout2.n125 vout2.n124 57.106
R373 vout2.n178 vout2.n177 48.2
R374 vout2.n179 vout2.n178 48.2
R375 vout2.n180 vout2.n179 48.2
R376 vout2.n181 vout2.n180 48.2
R377 vout2.n182 vout2.n181 48.2
R378 vout2.n172 vout2.n171 48.2
R379 vout2.n173 vout2.n172 48.2
R380 vout2.n174 vout2.n173 48.2
R381 vout2.n175 vout2.n174 48.2
R382 vout2.n176 vout2.n175 48.2
R383 vout2.n167 vout2.n166 48.2
R384 vout2.n168 vout2.n167 48.2
R385 vout2.n169 vout2.n168 48.2
R386 vout2.t3 vout2.n169 48.2
R387 vout2.n170 vout2.t3 48.2
R388 vout2.n161 vout2.n160 48.2
R389 vout2.n162 vout2.n161 48.2
R390 vout2.n163 vout2.n162 48.2
R391 vout2.n164 vout2.n163 48.2
R392 vout2.n165 vout2.n164 48.2
R393 vout2.n47 vout2.n46 48.2
R394 vout2.n46 vout2.n45 48.2
R395 vout2.n45 vout2.n44 48.2
R396 vout2.n44 vout2.n43 48.2
R397 vout2.n116 vout2.n115 48.2
R398 vout2.n115 vout2.n114 48.2
R399 vout2.n114 vout2.n113 48.2
R400 vout2.n113 vout2.n112 48.2
R401 vout2.n53 vout2.n52 48.2
R402 vout2.n52 vout2.n51 48.2
R403 vout2.n51 vout2.n50 48.2
R404 vout2.n50 vout2.n41 48.2
R405 vout2.n109 vout2.n108 48.2
R406 vout2.n108 vout2.n107 48.2
R407 vout2.n107 vout2.n106 48.2
R408 vout2.n106 vout2.n105 48.2
R409 vout2.n58 vout2.n57 48.2
R410 vout2.n57 vout2.n56 48.2
R411 vout2.n56 vout2.n55 48.2
R412 vout2.n55 vout2.n49 48.2
R413 vout2.n101 vout2.n100 48.2
R414 vout2.n100 vout2.n99 48.2
R415 vout2.n99 vout2.n98 48.2
R416 vout2.n98 vout2.n97 48.2
R417 vout2.n64 vout2.n63 48.2
R418 vout2.n63 vout2.n62 48.2
R419 vout2.n62 vout2.n61 48.2
R420 vout2.n61 vout2.n54 48.2
R421 vout2.n94 vout2.n93 48.2
R422 vout2.n93 vout2.n92 48.2
R423 vout2.n92 vout2.n91 48.2
R424 vout2.n91 vout2.n90 48.2
R425 vout2.n73 vout2.n72 48.2
R426 vout2.n72 vout2.n71 48.2
R427 vout2.n71 vout2.n70 48.2
R428 vout2.n70 vout2.n60 48.2
R429 vout2.n86 vout2.n85 48.2
R430 vout2.n85 vout2.n84 48.2
R431 vout2.n84 vout2.n83 48.2
R432 vout2.n83 vout2.n82 48.2
R433 vout2.n66 vout2.n65 48.2
R434 vout2.n67 vout2.n66 48.2
R435 vout2.n68 vout2.n67 48.2
R436 vout2.n69 vout2.n68 48.2
R437 vout2.n76 vout2.n75 48.2
R438 vout2.n77 vout2.n76 48.2
R439 vout2.n78 vout2.n77 48.2
R440 vout2.n79 vout2.n78 48.2
R441 vout2.n5 vout2.n4 48.2
R442 vout2.n6 vout2.n5 48.2
R443 vout2.n7 vout2.n6 48.2
R444 vout2.n8 vout2.n7 48.2
R445 vout2.n11 vout2.n10 48.2
R446 vout2.n12 vout2.n11 48.2
R447 vout2.n13 vout2.n12 48.2
R448 vout2.n14 vout2.n13 48.2
R449 vout2.n17 vout2.n16 48.2
R450 vout2.n18 vout2.n17 48.2
R451 vout2.n19 vout2.n18 48.2
R452 vout2.n20 vout2.n19 48.2
R453 vout2.n23 vout2.n22 48.2
R454 vout2.n24 vout2.n23 48.2
R455 vout2.n25 vout2.n24 48.2
R456 vout2.n26 vout2.n25 48.2
R457 vout2.n29 vout2.n28 48.2
R458 vout2.n30 vout2.n29 48.2
R459 vout2.n31 vout2.n30 48.2
R460 vout2.n32 vout2.n31 48.2
R461 vout2.n36 vout2.n35 48.2
R462 vout2.t2 vout2.n36 48.2
R463 vout2.n37 vout2.t2 48.2
R464 vout2.n38 vout2.n37 48.2
R465 vout2.n126 vout2.n125 48.2
R466 vout2.n127 vout2.n126 48.2
R467 vout2.n128 vout2.n127 48.2
R468 vout2.n129 vout2.n128 48.2
R469 vout2.n132 vout2.n131 48.2
R470 vout2.n133 vout2.n132 48.2
R471 vout2.n134 vout2.n133 48.2
R472 vout2.n135 vout2.n134 48.2
R473 vout2.n138 vout2.n137 48.2
R474 vout2.n139 vout2.n138 48.2
R475 vout2.n140 vout2.n139 48.2
R476 vout2.n141 vout2.n140 48.2
R477 vout2.n144 vout2.n143 48.2
R478 vout2.n145 vout2.n144 48.2
R479 vout2.n146 vout2.n145 48.2
R480 vout2.n147 vout2.n146 48.2
R481 vout2.n150 vout2.n149 48.2
R482 vout2.n151 vout2.n150 48.2
R483 vout2.n152 vout2.n151 48.2
R484 vout2.n153 vout2.n152 48.2
R485 vout2.n156 vout2.n155 48.2
R486 vout2.n157 vout2.n156 48.2
R487 vout2.n158 vout2.n157 48.2
R488 vout2.n159 vout2.n158 48.2
R489 vout2.n42 vout2 33.53
R490 vout2.n186 vout2.n159 26.731
R491 vout2.n185 vout2.n165 24.344
R492 vout2.n183 vout2.n176 24.1
R493 vout2.n184 vout2.n170 24.1
R494 vout2.n43 vout2.n42 24.1
R495 vout2.n119 vout2.n39 24.1
R496 vout2.n117 vout2.n116 24.1
R497 vout2.n111 vout2.n41 24.1
R498 vout2.n110 vout2.n109 24.1
R499 vout2.n103 vout2.n49 24.1
R500 vout2.n102 vout2.n101 24.1
R501 vout2.n96 vout2.n54 24.1
R502 vout2.n95 vout2.n94 24.1
R503 vout2.n88 vout2.n60 24.1
R504 vout2.n87 vout2.n86 24.1
R505 vout2.n81 vout2.n69 24.1
R506 vout2.n80 vout2.n79 24.1
R507 vout2.n9 vout2.n8 24.1
R508 vout2.n15 vout2.n14 24.1
R509 vout2.n21 vout2.n20 24.1
R510 vout2.n27 vout2.n26 24.1
R511 vout2.n33 vout2.n32 24.1
R512 vout2.n123 vout2.n38 24.1
R513 vout2.n121 vout2.n120 24.1
R514 vout2.n131 vout2.n130 24.1
R515 vout2.n137 vout2.n136 24.1
R516 vout2.n143 vout2.n142 24.1
R517 vout2.n149 vout2.n148 24.1
R518 vout2.n155 vout2.n154 24.1
R519 vout2.n104 vout2 18.267
R520 vout2.n74 vout2 18.069
R521 vout2.n89 vout2 17.808
R522 vout2.n48 vout2 16.443
R523 vout2.n123 vout2.n122 13.621
R524 vout2.n59 vout2 10.595
R525 vout2.n187 vout2.n186 8.052
R526 vout2.n89 vout2.n88 5.988
R527 vout2.n104 vout2.n103 5.089
R528 vout2.n80 vout2.n74 4.755
R529 vout2.n186 vout2.n185 3.567
R530 vout2.n110 vout2.n48 2.739
R531 vout2.n188 vout2.n3 2.727
R532 vout2.n95 vout2.n59 1.079
R533 vout2 vout2.n0 0.65
R534 vout2.n3 vout2.t4 0.608
R535 vout2.n2 vout2.n1 0.166
R536 vout2.n3 vout2.n2 0.033
R537 vout2.n2 vout2 0.014
R538 vout.n5 vout 1325.3
R539 vout.n6 vout.n5 1307.19
R540 vout vout.n284 1306.49
R541 vout.n8 vout.n7 1300.31
R542 vout.n0 vout 1297.81
R543 vout.n9 vout.n8 1289.42
R544 vout.n7 vout.n6 1286.35
R545 vout.n1 vout.n0 1281.21
R546 vout.n3 vout.n2 1278.32
R547 vout vout.n9 1277.28
R548 vout.n2 vout.n1 1275.19
R549 vout.n281 vout.n280 1275.03
R550 vout.n284 vout.n283 1273.91
R551 vout.n4 vout.n3 1272.1
R552 vout.n280 vout.n279 1270.16
R553 vout.n10 vout.n4 1255.59
R554 vout.n279 vout.n278 1214.9
R555 vout.n11 vout 706.558
R556 vout.n283 vout.n282 661.999
R557 vout.n10 vout 640.059
R558 vout.n282 vout.n281 631.752
R559 vout.n219 vout.n215 410.193
R560 vout.n226 vout.n225 409.266
R561 vout.n231 vout.n230 377.75
R562 vout.n239 vout.n238 372.189
R563 vout.n243 vout.n29 368.481
R564 vout.n247 vout.n17 366.628
R565 vout.n254 vout.n253 348.089
R566 vout.n142 vout.n135 345.308
R567 vout.n181 vout.n14 330.477
R568 vout.n197 vout.n39 327.696
R569 vout.n135 vout.n53 326.77
R570 vout.n201 vout.n45 325.843
R571 vout.n189 vout.n72 324.916
R572 vout.n115 vout.n90 321.208
R573 vout.n111 vout.n80 319.355
R574 vout.n173 vout.n172 316.034
R575 vout.n174 vout.n173 316.034
R576 vout.n178 vout.n174 316.034
R577 vout.n178 vout.n177 316.034
R578 vout.n111 vout.n86 314.72
R579 vout.n193 vout.n68 307.305
R580 vout.n115 vout.n76 302.67
R581 vout.n185 vout.n21 300.816
R582 vout.n131 vout.n60 299.889
R583 vout.n185 vout.n76 298.962
R584 vout.n127 vout.n102 297.108
R585 vout.n119 vout.n94 295.254
R586 vout.n243 vout.n25 293.4
R587 vout.n181 vout.n80 291.546
R588 vout.n201 vout.n60 289.693
R589 vout.n215 vout.n212 288.766
R590 vout.n123 vout.n98 288.766
R591 vout.n253 vout.n14 287.839
R592 vout.n172 vout.n171 286.736
R593 vout.n131 vout.n106 285.985
R594 vout.n239 vout.n33 284.131
R595 vout.n193 vout.n33 275.789
R596 vout.n230 vout.n39 275.788
R597 vout.n119 vout.n72 273.935
R598 vout.n247 vout.n21 273.008
R599 vout.n127 vout.n64 272.081
R600 vout.n123 vout.n68 270.227
R601 vout.n175 vout.n14 269.189
R602 vout.n81 vout.n80 269.161
R603 vout.n255 vout.n254 269.123
R604 vout.n111 vout.n110 269.075
R605 vout.n253 vout.n252 269.036
R606 vout.n181 vout.n180 269.014
R607 vout.n86 vout.n85 269.003
R608 vout.n170 vout.n169 268.657
R609 vout.n205 vout.n53 267.447
R610 vout.n189 vout.n25 266.519
R611 vout.n212 vout.n205 265.592
R612 vout.n226 vout.n45 260.958
R613 vout.n158 vout.n98 255.397
R614 vout.n106 vout.n105 252.315
R615 vout.n45 vout.n44 252.289
R616 vout.n131 vout.n130 252.282
R617 vout.n61 vout.n60 252.261
R618 vout.n201 vout.n200 252.151
R619 vout.n227 vout.n226 251.794
R620 vout.n225 vout.n224 251.722
R621 vout.n151 vout.n150 250.648
R622 vout.n135 vout.n134 250.306
R623 vout.n205 vout.n204 250.278
R624 vout.n57 vout.n53 250.256
R625 vout.n142 vout.n141 250.083
R626 vout.n220 vout.n219 249.928
R627 vout.n212 vout.n211 249.874
R628 vout.n215 vout.n214 249.406
R629 vout.n147 vout.n146 248.579
R630 vout.n257 vout.n12 239.118
R631 vout.n17 vout.n16 235.834
R632 vout.n197 vout.n64 230.37
R633 vout.n150 vout.n106 228.516
R634 vout vout.n12 221.524
R635 vout.n154 vout.n102 219.247
R636 vout.n21 vout.n20 217.516
R637 vout.n185 vout.n184 217.513
R638 vout.n77 vout.n76 217.512
R639 vout.n115 vout.n114 217.503
R640 vout.n248 vout.n247 217.431
R641 vout.n90 vout.n89 217.383
R642 vout.t1 vout.n166 216.609
R643 vout.n102 vout.n101 209.575
R644 vout.n155 vout.n154 208.613
R645 vout.n189 vout.n188 203.416
R646 vout.n123 vout.n122 203.368
R647 vout.n193 vout.n192 203.368
R648 vout.n98 vout.n97 203.368
R649 vout.n244 vout.n243 203.332
R650 vout.n119 vout.n118 203.303
R651 vout.n25 vout.n24 203.295
R652 vout.n33 vout.n32 203.271
R653 vout.n94 vout.n93 203.24
R654 vout.n240 vout.n239 203.22
R655 vout.n69 vout.n68 203.209
R656 vout.n73 vout.n72 203.129
R657 vout.n238 vout.n237 203.014
R658 vout.n29 vout.n28 202.828
R659 vout.n163 vout.n162 202.472
R660 vout.n159 vout.n158 201.492
R661 vout.n127 vout.n126 201.268
R662 vout.n65 vout.n64 201.242
R663 vout.n39 vout.n38 201.133
R664 vout.n230 vout.n41 200.984
R665 vout.n232 vout.n231 200.843
R666 vout.n169 vout.n86 200.708
R667 vout.n197 vout.n196 200.192
R668 vout.n166 vout.n90 190.512
R669 vout.n146 vout.n142 184.95
R670 vout.n162 vout.n94 171.974
R671 vout.n177 vout 94.509
R672 vout.n268 vout 69.482
R673 vout.n278 vout.n11 61.418
R674 vout.n259 vout.n258 48.2
R675 vout.n260 vout.n259 48.2
R676 vout.n261 vout.n260 48.2
R677 vout.n262 vout.n261 48.2
R678 vout.n263 vout.n262 48.2
R679 vout.n264 vout.n263 48.2
R680 vout.n265 vout.n264 48.2
R681 vout.n266 vout.n265 48.2
R682 vout.n267 vout.n266 48.2
R683 vout.n269 vout.n268 48.2
R684 vout.n270 vout.n269 48.2
R685 vout.n271 vout.n270 48.2
R686 vout.n272 vout.n271 48.2
R687 vout.n273 vout.n272 48.2
R688 vout.n274 vout.n273 48.2
R689 vout.n275 vout.n274 48.2
R690 vout.n276 vout.n275 48.2
R691 vout.t2 vout.n276 48.2
R692 vout.n130 vout.n129 48.2
R693 vout.n129 vout.n128 48.2
R694 vout.n122 vout.n121 48.2
R695 vout.n121 vout.n120 48.2
R696 vout.n82 vout.n81 48.2
R697 vout.n44 vout.n43 48.2
R698 vout.n43 vout.n42 48.2
R699 vout.n32 vout.n31 48.2
R700 vout.n31 vout.n30 48.2
R701 vout.n176 vout.n175 48.2
R702 vout.n19 vout.n18 48.2
R703 vout.n20 vout.n19 48.2
R704 vout.n217 vout.n216 48.2
R705 vout.n218 vout.n217 48.2
R706 vout.n222 vout.n221 48.2
R707 vout.n221 vout.n220 48.2
R708 vout.n48 vout.n47 48.2
R709 vout.n49 vout.n48 48.2
R710 vout.n207 vout.n206 48.2
R711 vout.n208 vout.n207 48.2
R712 vout.n214 vout.n213 48.2
R713 vout.n213 vout.n46 48.2
R714 vout.n224 vout.n223 48.2
R715 vout.n223 vout.n35 48.2
R716 vout.n233 vout.n232 48.2
R717 vout.n234 vout.n233 48.2
R718 vout.n41 vout.n40 48.2
R719 vout.n40 vout.n34 48.2
R720 vout.n237 vout.n236 48.2
R721 vout.n236 vout.n235 48.2
R722 vout.n28 vout.n27 48.2
R723 vout.n27 vout.n26 48.2
R724 vout.n15 vout.n13 48.2
R725 vout.n16 vout.n15 48.2
R726 vout.n245 vout.n244 48.2
R727 vout.n246 vout.n245 48.2
R728 vout.n250 vout.n249 48.2
R729 vout.n249 vout.n248 48.2
R730 vout.n23 vout.n22 48.2
R731 vout.n24 vout.n23 48.2
R732 vout.n242 vout.n241 48.2
R733 vout.n241 vout.n240 48.2
R734 vout.n37 vout.n36 48.2
R735 vout.n38 vout.n37 48.2
R736 vout.n229 vout.n228 48.2
R737 vout.n228 vout.n227 48.2
R738 vout.n210 vout.n209 48.2
R739 vout.n211 vout.n210 48.2
R740 vout.n55 vout.n54 48.2
R741 vout.n56 vout.n55 48.2
R742 vout.n203 vout.n202 48.2
R743 vout.n204 vout.n203 48.2
R744 vout.n51 vout.n50 48.2
R745 vout.n52 vout.n51 48.2
R746 vout.n108 vout.n107 48.2
R747 vout.n109 vout.n108 48.2
R748 vout.n58 vout.n57 48.2
R749 vout.n59 vout.n58 48.2
R750 vout.n200 vout.n199 48.2
R751 vout.n199 vout.n198 48.2
R752 vout.n196 vout.n195 48.2
R753 vout.n195 vout.n194 48.2
R754 vout.n66 vout.n65 48.2
R755 vout.n67 vout.n66 48.2
R756 vout.n192 vout.n191 48.2
R757 vout.n191 vout.n190 48.2
R758 vout.n188 vout.n187 48.2
R759 vout.n187 vout.n186 48.2
R760 vout.n74 vout.n73 48.2
R761 vout.n75 vout.n74 48.2
R762 vout.n184 vout.n183 48.2
R763 vout.n183 vout.n182 48.2
R764 vout.n180 vout.n179 48.2
R765 vout.n114 vout.n113 48.2
R766 vout.n113 vout.n112 48.2
R767 vout.n110 vout.n83 48.2
R768 vout.n79 vout.n78 48.2
R769 vout.n78 vout.n77 48.2
R770 vout.n117 vout.n116 48.2
R771 vout.n118 vout.n117 48.2
R772 vout.n71 vout.n70 48.2
R773 vout.n70 vout.n69 48.2
R774 vout.n125 vout.n124 48.2
R775 vout.n126 vout.n125 48.2
R776 vout.n63 vout.n62 48.2
R777 vout.n62 vout.n61 48.2
R778 vout.n133 vout.n132 48.2
R779 vout.n134 vout.n133 48.2
R780 vout.n137 vout.n136 48.2
R781 vout.n138 vout.n137 48.2
R782 vout.n140 vout.n139 48.2
R783 vout.n141 vout.n140 48.2
R784 vout.n144 vout.n143 48.2
R785 vout.n145 vout.n144 48.2
R786 vout.n148 vout.n147 48.2
R787 vout.n149 vout.n148 48.2
R788 vout.n153 vout.n152 48.2
R789 vout.n152 vout.n151 48.2
R790 vout.n105 vout.n104 48.2
R791 vout.n104 vout.n103 48.2
R792 vout.n100 vout.n99 48.2
R793 vout.n101 vout.n100 48.2
R794 vout.n156 vout.n155 48.2
R795 vout.n157 vout.n156 48.2
R796 vout.n161 vout.n160 48.2
R797 vout.n160 vout.n159 48.2
R798 vout.n97 vout.n96 48.2
R799 vout.n96 vout.n95 48.2
R800 vout.n92 vout.n91 48.2
R801 vout.n93 vout.n92 48.2
R802 vout.n164 vout.n163 48.2
R803 vout.n165 vout.n164 48.2
R804 vout.n168 vout.n167 48.2
R805 vout.n167 vout.t1 48.2
R806 vout.n89 vout.n88 48.2
R807 vout.n88 vout.n87 48.2
R808 vout.n85 vout.n84 48.2
R809 vout.n171 vout.n170 48.2
R810 vout.n252 vout.n251 48.2
R811 vout.n256 vout.n255 48.2
R812 vout vout.n267 42.373
R813 vout.n277 vout.t2 27.832
R814 vout.n257 vout.n256 25.813
R815 vout.n128 vout.n127 24.1
R816 vout.n120 vout.n119 24.1
R817 vout.n174 vout.n82 24.1
R818 vout.n42 vout.n39 24.1
R819 vout.n30 vout.n25 24.1
R820 vout.n177 vout.n176 24.1
R821 vout.n18 vout.n14 24.1
R822 vout.n219 vout.n218 24.1
R823 vout.n225 vout.n222 24.1
R824 vout.n215 vout.n49 24.1
R825 vout.n212 vout.n208 24.1
R826 vout.n226 vout.n46 24.1
R827 vout.n231 vout.n35 24.1
R828 vout.n238 vout.n234 24.1
R829 vout.n239 vout.n34 24.1
R830 vout.n235 vout.n29 24.1
R831 vout.n26 vout.n17 24.1
R832 vout.n254 vout.n13 24.1
R833 vout.n247 vout.n246 24.1
R834 vout.n253 vout.n250 24.1
R835 vout.n22 vout.n21 24.1
R836 vout.n243 vout.n242 24.1
R837 vout.n36 vout.n33 24.1
R838 vout.n230 vout.n229 24.1
R839 vout.n209 vout.n45 24.1
R840 vout.n205 vout.n56 24.1
R841 vout.n202 vout.n201 24.1
R842 vout.n53 vout.n52 24.1
R843 vout.n135 vout.n109 24.1
R844 vout.n60 vout.n59 24.1
R845 vout.n198 vout.n197 24.1
R846 vout.n194 vout.n193 24.1
R847 vout.n68 vout.n67 24.1
R848 vout.n190 vout.n189 24.1
R849 vout.n186 vout.n185 24.1
R850 vout.n76 vout.n75 24.1
R851 vout.n182 vout.n181 24.1
R852 vout.n179 vout.n178 24.1
R853 vout.n112 vout.n111 24.1
R854 vout.n173 vout.n83 24.1
R855 vout.n80 vout.n79 24.1
R856 vout.n116 vout.n115 24.1
R857 vout.n72 vout.n71 24.1
R858 vout.n124 vout.n123 24.1
R859 vout.n64 vout.n63 24.1
R860 vout.n132 vout.n131 24.1
R861 vout.n142 vout.n138 24.1
R862 vout.n139 vout.n106 24.1
R863 vout.n146 vout.n145 24.1
R864 vout.n150 vout.n149 24.1
R865 vout.n154 vout.n153 24.1
R866 vout.n103 vout.n102 24.1
R867 vout.n99 vout.n98 24.1
R868 vout.n158 vout.n157 24.1
R869 vout.n162 vout.n161 24.1
R870 vout.n95 vout.n94 24.1
R871 vout.n91 vout.n90 24.1
R872 vout.n166 vout.n165 24.1
R873 vout.n169 vout.n168 24.1
R874 vout.n87 vout.n86 24.1
R875 vout.n172 vout.n84 24.1
R876 vout.n251 vout.n12 24.1
R877 vout.n11 vout 12.891
R878 vout.n4 vout 11.115
R879 vout.n2 vout 10.302
R880 vout vout.n10 10.288
R881 vout.n280 vout 10.031
R882 vout.n0 vout 9.76
R883 vout.n6 vout 9.217
R884 vout.n284 vout 8.675
R885 vout.n279 vout 8.133
R886 vout.n3 vout 8.133
R887 vout.n9 vout 7.048
R888 vout.n8 vout 7.048
R889 vout.n7 vout 7.048
R890 vout.n281 vout 5.964
R891 vout.n283 vout 5.964
R892 vout.n5 vout 5.693
R893 vout.n1 vout 5.151
R894 vout vout.n277 4.084
R895 vout.n282 vout.t0 3.308
R896 vout.n278 vout 1.599
R897 vout.n277 vout.n257 0.575
R898 vcap.n22 vcap 1339.41
R899 vcap.n8 vcap.n7 1337.7
R900 vcap.n4 vcap.n3 1332.37
R901 vcap.n21 vcap.n5 1330.68
R902 vcap vcap.n22 1329.9
R903 vcap vcap.n0 1329.44
R904 vcap.n10 vcap.n9 1329.21
R905 vcap.n3 vcap.n2 1327.01
R906 vcap.n11 vcap.n10 1322.22
R907 vcap.n0 vcap 1321.63
R908 vcap.n5 vcap.n4 1319.78
R909 vcap.n1 vcap 1316.23
R910 vcap.n9 vcap.n8 1314.6
R911 vcap.n7 vcap.n6 1313.42
R912 vcap.n2 vcap.n1 1312.31
R913 vcap.n19 vcap.n11 1297.62
R914 vcap.n12 vcap 1234.9
R915 vcap vcap.n13 1222.32
R916 vcap.n6 vcap 1205.13
R917 vcap vcap.n18 1173.82
R918 vcap.n0 vcap.t0 1166.46
R919 vcap.n17 vcap.n16 1157.45
R920 vcap.n18 vcap.n17 1157.44
R921 vcap.n13 vcap.n12 1157.42
R922 vcap.n16 vcap.n15 870.815
R923 vcap.n14 vcap 681.578
R924 vcap vcap.n21 614.791
R925 vcap vcap.n20 607.702
R926 vcap.n15 vcap.n14 347.985
R927 vcap.n13 vcap 77.494
R928 vcap.n12 vcap 77.494
R929 vcap.n16 vcap 77.494
R930 vcap.n17 vcap 77.494
R931 vcap.n18 vcap 77.494
R932 vcap.n20 vcap.n19 49.009
R933 vcap.n14 vcap 16.076
R934 vcap.n20 vcap 11.818
R935 vcap.n0 vcap 6.1
R936 vcap.n22 vcap 4.575
R937 vcap.n19 vcap 4.572
R938 vcap.n21 vcap 4.397
R939 vcap.n1 vcap 3.812
R940 vcap.n15 vcap.t1 3.308
R941 vcap.n9 vcap 2.541
R942 vcap.n8 vcap 2.541
R943 vcap.n7 vcap 2.541
R944 vcap.n4 vcap 2.541
R945 vcap.n3 vcap 2.541
R946 vcap.n5 vcap 2.033
R947 vcap.n11 vcap 1.897
R948 vcap.n10 vcap 1.817
R949 vcap.n6 vcap 1.817
R950 vcap.n2 vcap 1.817
R951 vout3.n12 vout3.n11 643.741
R952 vout3.n13 vout3.n12 605.267
R953 vout3.n14 vout3.n13 605.248
R954 vout3.n16 vout3.n15 605.176
R955 vout3.n15 vout3.n14 604.644
R956 vout3.n9 vout3.t0 512.965
R957 vout3.n16 vout3.t1 310.422
R958 vout3.n11 vout3 258.793
R959 vout3.n3 vout3.t4 131.932
R960 vout3.n6 vout3.n5 75.994
R961 vout3.n2 vout3.n0 75.23
R962 vout3 vout3.n16 52.953
R963 vout3.n12 vout3 51.789
R964 vout3.n13 vout3 51.789
R965 vout3.n14 vout3 51.789
R966 vout3.n15 vout3 51.789
R967 vout3.n4 vout3.t3 50.61
R968 vout3.n10 vout3.n9 45.76
R969 vout3.n4 vout3.n3 32.776
R970 vout3 vout3.n10 19.454
R971 vout3.n3 vout3.n2 18.482
R972 vout3.n5 vout3.n4 13.653
R973 vout3.n11 vout3 13.309
R974 vout3.n0 vout3 12.498
R975 vout3.n9 vout3 7.05
R976 vout3.n7 vout3.n6 6.362
R977 vout3.n5 vout3.n2 1.556
R978 vout3.n10 vout3.n8 1.18
R979 vout3 vout3.n0 1.11
R980 vout3.n5 vout3 0.739
R981 vout3.n8 vout3.n7 0.394
R982 vout3.n8 vout3.t2 0.168
R983 vout3.n7 vout3.n1 0.098
R984 vout3.n6 vout3.n0 0.026
R985 a_83302_53375.n4 a_83302_53375.n2 454.539
R986 a_83302_53375.n2 a_83302_53375.n0 402.744
R987 a_83302_53375.n1 a_83302_53375.t7 313.3
R988 a_83302_53375.n0 a_83302_53375.t6 159.908
R989 a_83302_53375.n3 a_83302_53375.t4 132.929
R990 a_83302_53375.n5 a_83302_53375.t0 121.39
R991 a_83302_53375.t1 a_83302_53375.n5 105.108
R992 a_83302_53375.n0 a_83302_53375.t5 86.336
R993 a_83302_53375.n3 a_83302_53375.t2 70.758
R994 a_83302_53375.n5 a_83302_53375.n4 57.411
R995 a_83302_53375.n1 a_83302_53375.t3 51.574
R996 a_83302_53375.n2 a_83302_53375.n1 8.836
R997 a_83302_53375.n4 a_83302_53375.n3 5.505
C0 vin2 bot 168.81fF
C1 vcap bot 125.88fF
C2 vin1 bot 369.56fF
C3 vout bot 177.98fF
C4 vout1 bot 228.40fF
C5 vout2 bot 156.89fF
C6 vdda bot 4271.97fF
V1 net1 bot 1.8
V2 vin1 bot 1.2
L1 net2 vout 10m m=1
R2000 net1 net2 68 m=1
C10 vout vcap 47n m=1
C11 vcap bot 0.1u m=1
V3 vin2 bot 0.9
V4 bot GND 0
V5 vdda bot 3.3
.lib /home/vinodhini/open_pdks/sky130/sky130A/libs.tech/ngspice/sky130.lib.spice tt


.tran 1n 10m
.options gmin=1E-11
.save vout vout1 vout2 vout3
.control
run
plot v(vout) v(vout1) v(vout2) v(vout3)
let i=1
let a=unitvec(70)
while i<71
let z=i+1
meas tran te trig V(vout3) val=1.78 rise=i targ  V(vout3) val =1.78 rise=z
let a[i-1]=te
let i=i+1
end
let j=0
while j<70
print a[j]
let j=j+1
end
.endc

**** end user architecture code
**.ends
.GLOBAL GND
** flattened .save nodes


.end

