magic
tech sky130A
magscale 1 2
timestamp 1633948548
<< pwell >>
rect -226 3664 3298 3668
rect -226 -126 3316 3664
rect -234 -226 3316 -126
rect 3204 -230 3316 -226
<< mvpsubdiff >>
rect -226 3664 3298 3668
rect -226 3568 3316 3664
rect -226 1420 -108 3568
rect -226 694 -200 1420
rect -134 694 -108 1420
rect 3204 1568 3316 3568
rect 3204 842 3224 1568
rect 3290 842 3316 1568
rect -226 -126 -108 694
rect 3204 -126 3316 842
rect -234 -226 3316 -126
rect 3204 -230 3316 -226
<< mvpsubdiffcont >>
rect -200 694 -134 1420
rect 3224 842 3290 1568
<< poly >>
rect 220 3418 2816 3498
rect 168 2718 542 2792
rect 930 2720 1304 2794
rect 1764 2722 2138 2796
rect 2518 2724 2892 2798
rect 174 2028 548 2102
rect 940 2028 1314 2102
rect 1754 2024 2128 2098
rect 2498 2024 2872 2098
rect 174 1332 548 1406
rect 952 1328 1326 1402
rect 1732 1332 2106 1406
rect 2530 1328 2904 1402
rect 182 632 556 706
rect 948 636 1322 710
rect 1742 632 2116 706
rect 2534 640 2908 714
<< locali >>
rect -4 3358 2388 3366
rect -4 3304 2396 3358
rect 0 3166 62 3304
rect 776 3150 838 3304
rect 1556 3146 1618 3304
rect 2334 3160 2396 3304
rect -222 1420 -114 1558
rect -222 694 -200 1420
rect -134 694 -114 1420
rect -222 616 -114 694
rect 8 394 48 3104
rect 662 380 712 3086
rect 778 370 828 3076
rect 1442 378 1492 3084
rect 1568 390 1618 3096
rect 2220 388 2270 3094
rect 2340 384 2390 3090
rect 2998 384 3048 3090
rect 3204 1568 3312 1714
rect 3204 842 3224 1568
rect 3290 842 3312 1568
rect 3204 772 3312 842
rect 664 130 726 260
rect 1434 130 1496 282
rect 2214 130 2276 264
rect 2992 130 3054 260
rect 654 68 3054 130
rect 664 62 726 68
rect 2214 66 2276 68
rect 2992 62 3054 68
<< metal1 >>
rect -222 616 -114 1558
rect 3204 772 3312 1714
use sky130_fd_pr__nfet_g5v0d10v5_HTYTG7  sky130_fd_pr__nfet_g5v0d10v5_HTYTG7_0 ~/Documents/colpitts layout
timestamp 1633929031
transform 1 0 1525 0 1 1714
box -1525 -1714 1525 1714
<< end >>
