magic
tech sky130A
magscale 1 2
timestamp 1634564537
<< mvpsubdiffcont >>
rect 22980 54924 23102 55346
rect 24240 44696 25328 44998
rect 38946 44424 42360 45148
rect 68330 43808 68980 43950
<< mvnsubdiffcont >>
rect 280 56666 496 57816
rect 81910 54182 82086 54936
<< poly >>
rect 41738 64334 42170 64424
rect 41738 64098 41814 64334
rect 42072 64098 42170 64334
rect 41738 64030 42170 64098
rect 20700 54660 20840 54740
rect 20792 54424 20840 54660
rect 20700 54364 20840 54424
rect 23258 54734 23408 54810
rect 23258 54418 23294 54734
rect 23382 54418 23408 54734
rect 23258 54332 23408 54418
rect 77304 51022 77728 51078
rect 77304 50826 77348 51022
rect 77656 50826 77728 51022
rect 77304 50774 77728 50826
rect 30102 43952 31230 44070
rect 80846 39538 81140 39582
rect 80846 39410 80866 39538
rect 81116 39410 81140 39538
rect 80846 39390 81140 39410
rect 80178 26206 81252 26704
<< polycont >>
rect 41814 64098 42072 64334
rect 57780 60506 57972 61190
rect 20678 54424 20792 54660
rect 23294 54418 23382 54734
rect 77348 50826 77656 51022
rect 67818 43438 68110 43584
rect 80866 39410 81116 39538
<< locali >>
rect 56852 64504 56966 64938
rect 41772 64334 42106 64372
rect 41772 64098 41814 64334
rect 42072 64098 42106 64334
rect 41772 64076 42106 64098
rect 57706 61190 58040 61298
rect 57706 60506 57780 61190
rect 57972 60506 58040 61190
rect 57706 60396 58040 60506
rect 222 57816 554 57874
rect 222 56666 280 57816
rect 496 57298 554 57816
rect 496 57184 854 57298
rect 496 56666 554 57184
rect 57906 56922 58868 57112
rect 222 56552 554 56666
rect 20464 55532 23774 55614
rect 22916 55346 23202 55376
rect 22916 54924 22980 55346
rect 23102 55070 23202 55346
rect 23102 54924 23484 55070
rect 22916 54892 23484 54924
rect 22916 54860 23202 54892
rect 23278 54734 23414 54780
rect 20658 54660 20824 54672
rect 20658 54424 20678 54660
rect 20792 54424 20824 54660
rect 20658 54392 20824 54424
rect 23278 54418 23294 54734
rect 23382 54418 23414 54734
rect 23278 54366 23414 54418
rect 24498 45070 24856 52002
rect 58938 46504 59118 56840
rect 81894 54946 81928 54954
rect 81894 54936 82128 54946
rect 81894 54918 81910 54936
rect 81896 54182 81910 54918
rect 82086 54182 82128 54936
rect 81896 54108 82128 54182
rect 75934 48690 76256 51190
rect 77322 51022 77690 51054
rect 77322 50826 77348 51022
rect 77656 50826 77690 51022
rect 77322 50798 77690 50826
rect 58938 46342 66184 46504
rect 38714 45148 42794 45178
rect 24024 44998 25442 45070
rect 24024 44696 24240 44998
rect 25328 44696 25442 44998
rect 24024 44582 25442 44696
rect 38714 44424 38946 45148
rect 42360 44424 42794 45148
rect 38714 44308 42794 44424
rect 66242 43426 66422 46248
rect 68276 43950 69060 43984
rect 68276 43808 68330 43950
rect 68980 43808 69060 43950
rect 68276 43782 69060 43808
rect 67732 43614 68038 43628
rect 67732 43584 68228 43614
rect 67732 43438 67818 43584
rect 68110 43438 68228 43584
rect 67732 43396 68228 43438
rect 69568 41790 69838 41896
rect 80846 39538 81140 39582
rect 80846 39410 80866 39538
rect 81116 39410 81140 39538
rect 80846 39390 81140 39410
rect 40322 -496 40566 5796
rect 59718 -184 60160 5936
rect 67706 840 68258 5814
rect 74412 804 74964 5924
<< viali >>
rect 41840 64136 42022 64304
rect 57798 60588 57940 61090
rect 338 56766 438 57716
rect 58868 56840 59184 57288
rect 23006 55000 23088 55346
rect 20690 54456 20770 54624
rect 23316 54452 23374 54720
rect 81924 54218 82048 54890
rect 83382 53640 83448 53700
rect 83970 53550 84020 53606
rect 86270 53586 86316 53630
rect 83870 53460 83920 53498
rect 77384 50850 77634 51008
rect 75734 48226 76396 48690
rect 66184 46248 66696 46524
rect 24382 44696 25184 44984
rect 39408 44424 41694 45004
rect 68426 43844 68848 43922
rect 67844 43482 68066 43584
rect 80908 39444 81068 39522
rect 39836 -1246 41558 -496
rect 59520 -682 60594 -184
rect 67080 -192 69254 840
rect 73674 -228 75848 804
<< metal1 >>
rect 58792 78708 94938 78714
rect 788 76048 94938 78708
rect 3778 69202 4576 76048
rect 56220 73516 56604 76048
rect 58792 75912 94938 76048
rect 70984 72778 71248 75912
rect 77770 73944 77930 75912
rect 3778 68604 4600 69202
rect 3878 65778 4600 68604
rect 38838 65126 38848 65882
rect 39974 65126 39984 65882
rect 39286 64292 39472 65126
rect 41772 64304 42106 64372
rect 41772 64292 41840 64304
rect 39286 64162 41840 64292
rect 41772 64136 41840 64162
rect 42022 64136 42106 64304
rect 41772 64076 42106 64136
rect 57706 61090 58040 61298
rect 57706 60588 57798 61090
rect 57940 60948 58040 61090
rect 59906 60948 60318 60972
rect 57940 60764 60318 60948
rect 57940 60588 58040 60764
rect 57706 60396 58040 60588
rect 222 57716 554 57874
rect 222 56766 338 57716
rect 438 56766 554 57716
rect 58862 57288 59190 57300
rect 58862 56840 58868 57288
rect 59184 57078 59190 57288
rect 59226 57078 59236 57262
rect 59184 56938 59236 57078
rect 59184 56840 59190 56938
rect 59226 56850 59236 56938
rect 59510 56850 59520 57262
rect 58862 56828 59190 56840
rect 222 56552 554 56766
rect 30970 55602 30980 55738
rect 29968 55538 30980 55602
rect 30970 55430 30980 55538
rect 31268 55430 31278 55738
rect 22916 55346 23202 55376
rect 22916 55000 23006 55346
rect 23088 55000 23202 55346
rect 22916 54860 23202 55000
rect 23278 54720 23414 54780
rect 20658 54628 20824 54672
rect 21354 54628 21608 54638
rect 23278 54628 23316 54720
rect 20658 54624 23316 54628
rect 20658 54456 20690 54624
rect 20770 54504 23316 54624
rect 20770 54456 20824 54504
rect 20658 54392 20824 54456
rect 21354 49318 21608 54504
rect 23278 54452 23316 54504
rect 23374 54452 23414 54720
rect 23278 54366 23414 54452
rect 59906 50432 60318 60764
rect 81894 54946 81928 54954
rect 81894 54918 82128 54946
rect 81896 54890 82128 54918
rect 81896 54218 81924 54890
rect 82048 54294 82128 54890
rect 83280 54294 83328 54300
rect 82048 54218 83332 54294
rect 81896 54146 83332 54218
rect 81896 54108 82128 54146
rect 83004 54070 83090 54146
rect 82966 53912 82976 54070
rect 83164 53912 83174 54070
rect 83280 53962 83328 54146
rect 83370 53700 83460 53706
rect 83370 53682 83382 53700
rect 82548 53468 82558 53658
rect 82674 53584 82684 53658
rect 83236 53652 83382 53682
rect 83370 53640 83382 53652
rect 83448 53640 83460 53700
rect 83370 53634 83460 53640
rect 86258 53630 86328 53636
rect 83964 53606 84026 53618
rect 83964 53584 83970 53606
rect 82674 53550 83970 53584
rect 84020 53550 84026 53606
rect 86258 53586 86270 53630
rect 86316 53590 86440 53630
rect 86316 53586 86328 53590
rect 86258 53580 86328 53586
rect 82674 53538 84026 53550
rect 82674 53528 83248 53538
rect 82674 53468 82684 53528
rect 83858 53498 83932 53504
rect 82998 53424 83008 53498
rect 83100 53492 83110 53498
rect 83100 53490 83758 53492
rect 83858 53490 83870 53498
rect 83100 53460 83870 53490
rect 83920 53460 83932 53498
rect 83100 53454 83932 53460
rect 83100 53452 83880 53454
rect 83100 53450 83758 53452
rect 83100 53424 83110 53450
rect 86140 51866 86212 53374
rect 88266 51866 88276 51918
rect 86140 51792 88276 51866
rect 86140 51778 86212 51792
rect 88266 51730 88276 51792
rect 88474 51730 88484 51918
rect 77322 51022 77690 51054
rect 77294 51008 77690 51022
rect 77294 50850 77384 51008
rect 77634 50850 77690 51008
rect 77294 50798 77690 50850
rect 59872 49850 68038 50432
rect 59906 49814 60318 49850
rect 21354 46432 21634 49318
rect 38414 47838 38424 48764
rect 39756 47838 39766 48764
rect 21354 46256 21640 46432
rect 21384 42946 21640 46256
rect 39090 45178 39496 47838
rect 66814 46560 66824 46688
rect 66550 46530 66824 46560
rect 66172 46524 66824 46530
rect 66172 46248 66184 46524
rect 66696 46248 66824 46524
rect 66172 46242 66824 46248
rect 66550 46158 66824 46242
rect 66814 45974 66824 46158
rect 67244 45974 67254 46688
rect 24024 44984 25442 45070
rect 24024 44696 24382 44984
rect 25184 44696 25442 44984
rect 24024 44582 25442 44696
rect 38714 45004 42794 45178
rect 38714 44424 39408 45004
rect 41694 44424 42794 45004
rect 38714 44308 42794 44424
rect 67818 43628 68038 49850
rect 75722 48690 76408 48696
rect 75722 48226 75734 48690
rect 76396 48226 76408 48690
rect 75722 48220 76408 48226
rect 68188 47424 68198 47812
rect 68884 47424 68894 47812
rect 75960 47790 76198 48220
rect 77294 48002 77620 50798
rect 68408 43984 68610 47424
rect 75714 47308 75724 47790
rect 76368 47308 76378 47790
rect 73050 46020 73060 46882
rect 73674 46672 73684 46882
rect 77264 46672 77620 48002
rect 73674 46636 77620 46672
rect 80598 46636 80954 46672
rect 73674 46204 80954 46636
rect 73674 46020 73684 46204
rect 68276 43922 69060 43984
rect 68276 43844 68426 43922
rect 68848 43844 69060 43922
rect 68276 43782 69060 43844
rect 67732 43614 68038 43628
rect 67732 43584 68228 43614
rect 67732 43482 67844 43584
rect 68066 43482 68228 43584
rect 67732 43396 68228 43482
rect 79160 43104 79170 43578
rect 79870 43104 79880 43578
rect 79424 43100 79728 43104
rect 79424 43084 79608 43100
rect 1264 -3192 1560 41416
rect 7722 40838 8018 41824
rect 14216 40876 14512 41602
rect 7722 40536 8496 40838
rect 13786 40574 14512 40876
rect 20748 40840 21044 41712
rect 62116 41292 62296 41604
rect 7722 -3192 8018 40536
rect 14216 -3192 14512 40574
rect 20338 40538 21044 40840
rect 20748 -3192 21044 40538
rect 27278 -3192 27574 40970
rect 33848 -3192 34144 40896
rect 40304 5642 40638 41156
rect 59632 41040 62296 41292
rect 46836 5684 47170 40858
rect 53442 5720 53776 41008
rect 46836 5478 47736 5684
rect 53392 5514 54196 5720
rect 59680 5702 60012 41040
rect 62116 39622 62296 41040
rect 65952 39622 66228 42408
rect 69708 39622 69984 42468
rect 73598 39634 73874 42542
rect 79424 41422 79538 43084
rect 80598 41576 80954 46204
rect 88542 42666 88552 43684
rect 89804 42666 89814 43684
rect 79422 41196 80188 41422
rect 76654 39634 76954 39646
rect 73508 39622 76954 39634
rect 62116 39454 76954 39622
rect 62140 39418 73870 39454
rect 65952 39370 66228 39418
rect 76654 38662 76954 39454
rect 80106 39474 80188 41196
rect 80598 39582 80952 41576
rect 86688 40886 87154 40908
rect 88846 40886 89414 42666
rect 86626 40396 89414 40886
rect 80598 39522 81140 39582
rect 80106 39470 80530 39474
rect 80598 39470 80908 39522
rect 80106 39410 80534 39470
rect 80440 39050 80534 39410
rect 80846 39444 80908 39470
rect 81068 39444 81140 39522
rect 80846 39390 81140 39444
rect 86688 38762 87154 40396
rect 88846 40376 89414 40396
rect 76680 34874 76932 36478
rect 80016 34874 80268 36478
rect 81094 34874 81226 35554
rect 83336 34874 83588 36436
rect 86710 34874 86962 36510
rect 76680 34670 86964 34874
rect 83336 34628 83588 34670
rect 53442 5494 53776 5514
rect 59364 5478 60012 5702
rect 67596 5592 68186 23790
rect 46836 5344 47170 5478
rect 59680 3574 60012 5478
rect 74374 5408 74964 23606
rect 39690 2594 39982 3390
rect 75142 2594 75380 3416
rect 39688 2392 75380 2594
rect 75142 2284 75380 2392
rect 67068 840 69266 846
rect 59508 -184 60606 -178
rect 39824 -496 41570 -490
rect 39824 -1246 39836 -496
rect 41558 -1246 41570 -496
rect 59508 -682 59520 -184
rect 60594 -682 60606 -184
rect 67068 -192 67080 840
rect 69254 -192 69266 840
rect 67068 -198 69266 -192
rect 73662 804 75860 810
rect 59508 -688 60606 -682
rect 39824 -1252 41570 -1246
rect 40284 -3192 40658 -1252
rect 59810 -3192 60142 -688
rect 67632 -3192 68480 -198
rect 73662 -228 73674 804
rect 75848 -228 75860 804
rect 73662 -234 75860 -228
rect 74154 -3192 75258 -234
rect 80820 -3192 81372 23754
rect 87672 3590 88224 23606
rect 87006 3340 88224 3590
rect 87672 -3192 88224 3340
rect 94120 -3192 94672 23348
rect 100788 -3192 101376 22686
rect 101856 -3192 111286 -3176
rect -588 -9218 111286 -3192
rect 101856 -9328 111286 -9218
<< via1 >>
rect 38848 65126 39974 65882
rect 59236 56850 59510 57262
rect 30980 55430 31268 55738
rect 82976 53912 83164 54070
rect 82558 53468 82674 53658
rect 83008 53424 83100 53498
rect 88276 51730 88474 51918
rect 38424 47838 39756 48764
rect 66824 45974 67244 46688
rect 68198 47424 68884 47812
rect 75724 47308 76368 47790
rect 73060 46020 73674 46882
rect 79170 43104 79870 43578
rect 88552 42666 89804 43684
<< metal2 >>
rect 38848 67730 39922 67740
rect 38848 66930 39922 66940
rect 39152 65892 39538 66930
rect 38848 65882 39974 65892
rect 38848 65116 39974 65126
rect 60520 57272 60932 57282
rect 59236 57262 59510 57272
rect 59510 56956 60520 57174
rect 59236 56840 59510 56850
rect 60520 56770 60932 56780
rect 31454 55766 31654 55776
rect 30980 55738 31268 55748
rect 31268 55524 31454 55630
rect 30980 55420 31268 55430
rect 31454 55398 31654 55408
rect 82976 54070 83164 54080
rect 82976 53902 83164 53912
rect 82558 53658 82674 53668
rect 82674 53468 82680 53654
rect 83018 53508 83086 53902
rect 82558 53458 82680 53468
rect 82568 51232 82680 53458
rect 83008 53498 83100 53508
rect 83008 53414 83100 53424
rect 89286 51966 89526 51976
rect 88276 51918 88474 51928
rect 88474 51860 89118 51864
rect 88474 51794 89286 51860
rect 89034 51790 89286 51794
rect 88276 51720 88474 51730
rect 89526 51790 89544 51860
rect 89286 51720 89526 51730
rect 82500 51222 82792 51232
rect 82500 50964 82792 50974
rect 38454 50414 39552 50424
rect 38454 49652 39552 49662
rect 68170 50012 68902 50022
rect 38540 48774 39118 49652
rect 68170 49466 68902 49476
rect 38424 48764 39756 48774
rect 38424 47828 39756 47838
rect 68312 47822 68620 49466
rect 68198 47812 68884 47822
rect 68198 47414 68884 47424
rect 75724 47790 76368 47800
rect 75724 47298 76368 47308
rect 73060 46882 73674 46892
rect 66824 46688 67244 46698
rect 67244 46212 73060 46578
rect 73060 46010 73674 46020
rect 66824 45964 67244 45974
rect 75884 45904 76188 47298
rect 77922 45994 78764 46004
rect 75856 45858 76958 45904
rect 75828 45650 77922 45858
rect 75856 45560 77922 45650
rect 75856 45180 76182 45560
rect 76398 45544 77922 45560
rect 77922 45280 78764 45290
rect 88708 45818 89786 45828
rect 88708 45240 89786 45250
rect 75856 45076 76228 45180
rect 75856 45054 76188 45076
rect 75866 43464 76188 45054
rect 88982 43694 89414 45240
rect 88552 43684 89804 43694
rect 79170 43578 79870 43588
rect 75866 43200 79170 43464
rect 75866 43190 76188 43200
rect 79170 43100 79870 43104
rect 79170 43094 79608 43100
rect 79798 43094 79870 43100
rect 88552 42656 89804 42666
<< via2 >>
rect 38848 66940 39922 67730
rect 60520 56780 60932 57272
rect 31454 55408 31654 55766
rect 89286 51730 89526 51966
rect 82500 50974 82792 51222
rect 38454 49662 39552 50414
rect 68170 49476 68902 50012
rect 77922 45290 78764 45994
rect 88708 45250 89786 45818
<< metal3 >>
rect 39024 68250 39034 69308
rect 39622 68250 39632 69308
rect 39184 67735 39488 68250
rect 38838 67730 39932 67735
rect 38838 66940 38848 67730
rect 39922 66940 39932 67730
rect 38838 66935 39932 66940
rect 60510 57272 60942 57277
rect 60510 56780 60520 57272
rect 60932 57148 60942 57272
rect 61028 57148 61038 57236
rect 60932 56928 61038 57148
rect 60932 56780 60942 56928
rect 61028 56780 61038 56928
rect 61372 56780 61382 57236
rect 60510 56775 60942 56780
rect 31444 55766 31664 55771
rect 31444 55408 31454 55766
rect 31654 55644 31664 55766
rect 31760 55644 31770 55766
rect 31654 55508 31770 55644
rect 31654 55408 31664 55508
rect 31444 55403 31664 55408
rect 31760 55386 31770 55508
rect 32028 55386 32038 55766
rect 68320 53232 68550 55528
rect 38598 50419 38946 51802
rect 38444 50414 39562 50419
rect 38444 49662 38454 50414
rect 39552 49662 39562 50414
rect 68320 50017 68576 53232
rect 89276 51966 89536 51971
rect 89276 51730 89286 51966
rect 89526 51730 89536 51966
rect 89276 51725 89536 51730
rect 89340 51408 89478 51725
rect 82490 51222 82802 51227
rect 82490 50974 82500 51222
rect 82792 50974 82802 51222
rect 82490 50969 82802 50974
rect 82562 50666 82690 50969
rect 82428 50454 82438 50666
rect 82798 50454 82808 50666
rect 38444 49657 39562 49662
rect 68160 50012 68912 50017
rect 68160 49476 68170 50012
rect 68902 49476 68912 50012
rect 68160 49471 68912 49476
rect 89350 47658 89462 51408
rect 83032 47638 88248 47658
rect 88904 47638 89472 47658
rect 83032 47384 89472 47638
rect 83032 47346 88248 47384
rect 77912 45994 78774 45999
rect 77912 45290 77922 45994
rect 78764 45818 78774 45994
rect 81260 45818 81270 46190
rect 78764 45408 81270 45818
rect 78764 45290 78774 45408
rect 77912 45285 78774 45290
rect 81260 45270 81270 45408
rect 81936 45270 81946 46190
rect 88904 45823 89472 47384
rect 88698 45818 89796 45823
rect 88698 45250 88708 45818
rect 89786 45250 89796 45818
rect 88698 45245 89796 45250
<< via3 >>
rect 39034 68250 39622 69308
rect 61038 56780 61372 57236
rect 31770 55386 32028 55766
rect 82438 50454 82798 50666
rect 81270 45270 81936 46190
<< metal4 >>
rect 39033 69308 39623 69309
rect 39033 69224 39034 69308
rect 32146 68754 39034 69224
rect 32162 66334 32516 68754
rect 39033 68250 39034 68754
rect 39622 68250 39623 69308
rect 39033 68249 39623 68250
rect 61037 57236 61373 57237
rect 61037 56780 61038 57236
rect 61372 57130 61373 57236
rect 61372 56928 61942 57130
rect 61372 56780 61373 56928
rect 61037 56779 61373 56780
rect 31769 55766 32029 55767
rect 31769 55386 31770 55766
rect 32028 55624 32029 55766
rect 32028 55494 32408 55624
rect 32028 55386 32029 55494
rect 31769 55385 32029 55386
rect 82437 50666 82799 50667
rect 82437 50454 82438 50666
rect 82798 50454 82799 50666
rect 82437 50453 82799 50454
rect 82546 50030 82702 50453
rect 82462 50010 82908 50030
rect 82462 49486 84228 50010
rect 82462 48376 82908 49486
rect 82446 47596 82908 48376
rect 81269 46190 81937 46191
rect 81269 45270 81270 46190
rect 81936 46092 81937 46190
rect 82462 46092 82908 47596
rect 81936 45686 82908 46092
rect 81936 45642 84208 45686
rect 81936 45270 81937 45642
rect 81269 45269 81937 45270
rect 82462 45144 84208 45642
use nmos551020guard  nmos551020guard_0 ~/layout test
timestamp 1634553547
transform 1 0 60534 0 1 1904
box 0 -60 40992 25660
use nmos3346guard  nmos3346guard_0 ~/layout test
timestamp 1634226173
transform 1 0 76634 0 1 35100
box -198 -464 10640 4940
use pmos33431guard  pmos33431guard_0 ~/layout test
timestamp 1634274673
transform 1 0 70594 0 1 50830
box -52 -1146 11632 24722
use pmos33823guard  pmos33823guard_0 ~/layout test
timestamp 1634123280
transform 0 1 62 -1 0 66356
box 0 -28 19500 21152
use nmos33210guard  nmos33210guard_0 ~/layout test
timestamp 1634117422
transform 0 1 23394 -1 0 57492
box -692 -504 5802 7534
use cap5p  cap5p_0 ~/layout test
timestamp 1634206023
transform 0 -1 38214 -1 0 51430
box -17168 -670 4272 6120
use pmos331020guard  pmos331020guard_0
timestamp 1634186000
transform 0 1 41674 -1 0 74064
box 0 -76 26862 16672
use cap3p  cap3p_0
timestamp 1634206384
transform 0 -1 67632 -1 0 55396
box -8584 -1022 4272 6028
use nmos3355guard  nmos3355guard_0
timestamp 1634141228
transform 1 0 62148 0 1 39920
box -212 -578 12082 4120
use sky130_fd_pr__cap_mim_m3_1_DAF5A5  sky130_fd_pr__cap_mim_m3_1_DAF5A5_0 ~/layout test
timestamp 1634365921
transform 0 1 85636 -1 0 47470
box -4282 -2600 4282 2600
use sky130_fd_sc_hvl__dfrtp_1  sky130_fd_sc_hvl__dfrtp_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1632099954
transform 1 0 83272 0 1 53268
box -66 -43 3138 897
use nmos551535  nmos551535_0 ~/layout test
timestamp 1634301196
transform 1 0 -25528 0 1 2780
box 25528 -2780 85820 42652
<< labels >>
flabel poly 30710 44036 30710 44036 0 FreeSans 4800 0 0 0 vin1
flabel metal1 21456 45972 21456 45972 0 FreeSans 1600 0 0 0 vout
flabel locali 21634 55558 21634 55558 0 FreeSans 1600 0 0 0 vout1
flabel locali 61674 46392 61674 46392 0 FreeSans 1600 0 0 0 vout2
flabel metal1 4286 77500 4286 77500 0 FreeSans 1600 0 0 0 vdda
rlabel metal3 88528 47472 88528 47472 5 bot
flabel locali 76018 49066 76018 49066 0 FreeSans 1600 0 0 0 vout3
flabel metal1 86350 53606 86350 53606 0 FreeSans 800 0 0 0 dfout
flabel metal1 83702 53468 83702 53468 0 FreeSans 800 0 0 0 reset
flabel metal1 83258 53670 83258 53670 0 FreeSans 800 0 0 0 clkin
flabel metal1 1910 -6426 1910 -6426 0 FreeSans 1600 0 0 0 vssa
flabel metal1 46520 2470 46520 2470 0 FreeSans 1600 0 0 0 vcap
flabel poly 80634 26412 80658 26412 0 FreeSans 1600 0 0 0 vin2
<< end >>
