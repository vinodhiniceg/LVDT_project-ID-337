magic
tech sky130A
magscale 1 2
timestamp 1634616792
<< mvnmos >>
rect -287 194 -187 394
rect -129 194 -29 394
rect 29 194 129 394
rect 187 194 287 394
rect -287 -100 -187 100
rect -129 -100 -29 100
rect 29 -100 129 100
rect 187 -100 287 100
rect -287 -394 -187 -194
rect -129 -394 -29 -194
rect 29 -394 129 -194
rect 187 -394 287 -194
<< mvndiff >>
rect -345 320 -287 394
rect -345 268 -333 320
rect -299 268 -287 320
rect -345 194 -287 268
rect -187 320 -129 394
rect -187 268 -175 320
rect -141 268 -129 320
rect -187 194 -129 268
rect -29 320 29 394
rect -29 268 -17 320
rect 17 268 29 320
rect -29 194 29 268
rect 129 320 187 394
rect 129 268 141 320
rect 175 268 187 320
rect 129 194 187 268
rect 287 320 345 394
rect 287 268 299 320
rect 333 268 345 320
rect 287 194 345 268
rect -345 26 -287 100
rect -345 -26 -333 26
rect -299 -26 -287 26
rect -345 -100 -287 -26
rect -187 26 -129 100
rect -187 -26 -175 26
rect -141 -26 -129 26
rect -187 -100 -129 -26
rect -29 26 29 100
rect -29 -26 -17 26
rect 17 -26 29 26
rect -29 -100 29 -26
rect 129 26 187 100
rect 129 -26 141 26
rect 175 -26 187 26
rect 129 -100 187 -26
rect 287 26 345 100
rect 287 -26 299 26
rect 333 -26 345 26
rect 287 -100 345 -26
rect -345 -268 -287 -194
rect -345 -320 -333 -268
rect -299 -320 -287 -268
rect -345 -394 -287 -320
rect -187 -268 -129 -194
rect -187 -320 -175 -268
rect -141 -320 -129 -268
rect -187 -394 -129 -320
rect -29 -268 29 -194
rect -29 -320 -17 -268
rect 17 -320 29 -268
rect -29 -394 29 -320
rect 129 -268 187 -194
rect 129 -320 141 -268
rect 175 -320 187 -268
rect 129 -394 187 -320
rect 287 -268 345 -194
rect 287 -320 299 -268
rect 333 -320 345 -268
rect 287 -394 345 -320
<< mvndiffc >>
rect -333 268 -299 320
rect -175 268 -141 320
rect -17 268 17 320
rect 141 268 175 320
rect 299 268 333 320
rect -333 -26 -299 26
rect -175 -26 -141 26
rect -17 -26 17 26
rect 141 -26 175 26
rect 299 -26 333 26
rect -333 -320 -299 -268
rect -175 -320 -141 -268
rect -17 -320 17 -268
rect 141 -320 175 -268
rect 299 -320 333 -268
<< poly >>
rect -287 394 -187 420
rect -129 394 -29 420
rect 29 394 129 420
rect 187 394 287 420
rect -287 168 -187 194
rect -129 168 -29 194
rect 29 168 129 194
rect 187 168 287 194
rect -287 100 -187 126
rect -129 100 -29 126
rect 29 100 129 126
rect 187 100 287 126
rect -287 -126 -187 -100
rect -129 -126 -29 -100
rect 29 -126 129 -100
rect 187 -126 287 -100
rect -287 -194 -187 -168
rect -129 -194 -29 -168
rect 29 -194 129 -168
rect 187 -194 287 -168
rect -287 -420 -187 -394
rect -129 -420 -29 -394
rect 29 -420 129 -394
rect 187 -420 287 -394
<< locali >>
rect -333 320 -299 336
rect -333 252 -299 268
rect -175 320 -141 336
rect -175 252 -141 268
rect -17 320 17 336
rect -17 252 17 268
rect 141 320 175 336
rect 141 252 175 268
rect 299 320 333 336
rect 299 252 333 268
rect -333 26 -299 42
rect -333 -42 -299 -26
rect -175 26 -141 42
rect -175 -42 -141 -26
rect -17 26 17 42
rect -17 -42 17 -26
rect 141 26 175 42
rect 141 -42 175 -26
rect 299 26 333 42
rect 299 -42 333 -26
rect -333 -268 -299 -252
rect -333 -336 -299 -320
rect -175 -268 -141 -252
rect -175 -336 -141 -320
rect -17 -268 17 -252
rect -17 -336 17 -320
rect 141 -268 175 -252
rect 141 -336 175 -320
rect 299 -268 333 -252
rect 299 -336 333 -320
<< viali >>
rect -333 268 -299 320
rect -175 268 -141 320
rect -17 268 17 320
rect 141 268 175 320
rect 299 268 333 320
rect -333 -26 -299 26
rect -175 -26 -141 26
rect -17 -26 17 26
rect 141 -26 175 26
rect 299 -26 333 26
rect -333 -320 -299 -268
rect -175 -320 -141 -268
rect -17 -320 17 -268
rect 141 -320 175 -268
rect 299 -320 333 -268
<< metal1 >>
rect -339 320 -293 332
rect -339 268 -333 320
rect -299 268 -293 320
rect -339 256 -293 268
rect -181 320 -135 332
rect -181 268 -175 320
rect -141 268 -135 320
rect -181 256 -135 268
rect -23 320 23 332
rect -23 268 -17 320
rect 17 268 23 320
rect -23 256 23 268
rect 135 320 181 332
rect 135 268 141 320
rect 175 268 181 320
rect 135 256 181 268
rect 293 320 339 332
rect 293 268 299 320
rect 333 268 339 320
rect 293 256 339 268
rect -339 26 -293 38
rect -339 -26 -333 26
rect -299 -26 -293 26
rect -339 -38 -293 -26
rect -181 26 -135 38
rect -181 -26 -175 26
rect -141 -26 -135 26
rect -181 -38 -135 -26
rect -23 26 23 38
rect -23 -26 -17 26
rect 17 -26 23 26
rect -23 -38 23 -26
rect 135 26 181 38
rect 135 -26 141 26
rect 175 -26 181 26
rect 135 -38 181 -26
rect 293 26 339 38
rect 293 -26 299 26
rect 333 -26 339 26
rect 293 -38 339 -26
rect -339 -268 -293 -256
rect -339 -320 -333 -268
rect -299 -320 -293 -268
rect -339 -332 -293 -320
rect -181 -268 -135 -256
rect -181 -320 -175 -268
rect -141 -320 -135 -268
rect -181 -332 -135 -320
rect -23 -268 23 -256
rect -23 -320 -17 -268
rect 17 -320 23 -268
rect -23 -332 23 -320
rect 135 -268 181 -256
rect 135 -320 141 -268
rect 175 -320 181 -268
rect 135 -332 181 -320
rect 293 -268 339 -256
rect 293 -320 299 -268
rect 333 -320 339 -268
rect 293 -332 339 -320
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string parameters w 1 l 0.5 m 3 nf 4 diffcov 30 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 30 viadrn 30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
