magic
tech sky130A
magscale 1 2
timestamp 1634046259
<< error_s >>
rect 4116 7552 4174 8308
rect 4110 7524 4176 7552
rect 4116 6308 4174 7524
rect 6174 6308 6232 8308
rect 4116 4214 4174 6214
rect 6174 4214 6232 6214
rect 4116 2120 4174 4120
rect 6174 2120 6232 4120
rect 4116 26 4174 2026
rect 6174 26 6232 2026
<< mvpsubdiff >>
rect -1062 7396 -492 7596
rect -1062 1444 -924 7396
rect -616 1444 -492 7396
rect -1062 874 -492 1444
<< mvpsubdiffcont >>
rect -924 1444 -616 7396
<< poly >>
rect 744 8326 4702 8380
rect 500 6228 1734 6288
rect 2546 6230 3780 6290
rect 4820 6230 6054 6290
rect 460 4138 1694 4198
rect 2628 4136 3862 4196
rect 4698 4138 5932 4198
rect 322 2044 1556 2104
rect 2624 2042 3858 2102
rect 4678 2044 5912 2104
<< locali >>
rect -4 8168 54 8202
rect 4110 8168 4176 8176
rect -4 8070 4176 8168
rect -4 8056 190 8070
rect -8 8000 190 8056
rect -1062 7396 -492 7596
rect -8 7404 58 8000
rect 4110 7524 4176 8070
rect -1062 1444 -924 7396
rect -616 1444 -492 7396
rect -1062 874 -492 1444
rect 0 1062 54 7404
rect 2062 1062 2116 7492
rect 4120 1088 4174 7518
rect 6178 1112 6232 7542
rect 2060 392 2106 926
rect 6178 392 6222 836
rect 2060 276 6230 392
rect 6178 268 6222 276
<< viali >>
rect -878 1736 -738 6980
<< metal1 >>
rect -1062 6980 -492 7596
rect -1062 1736 -878 6980
rect -738 1736 -492 6980
rect -1062 874 -492 1736
use sky130_fd_pr__nfet_g5v0d10v5_S5TLYR  sky130_fd_pr__nfet_g5v0d10v5_S5TLYR_0
timestamp 1634046259
transform 1 0 3116 0 1 4167
box -3116 -4167 3116 4167
<< end >>
