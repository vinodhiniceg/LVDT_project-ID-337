magic
tech sky130A
timestamp 1634049493
<< pwell >>
rect -89 10961 6980 11293
rect -89 10797 406 10961
rect 480 10887 6980 10961
rect 480 10797 6426 10887
rect -89 10707 6426 10797
rect 6540 10707 6980 10887
rect -89 -331 6980 10707
rect -89 -3599 3751 -331
rect 4059 -362 6980 -331
rect 4157 -3599 6980 -362
rect -89 -4250 6980 -3599
<< poly >>
rect 2983 11191 5183 11252
rect 2985 11068 3118 11191
rect 5047 11033 5180 11191
rect 961 5399 1143 5846
rect 1862 5400 2044 5847
rect 2900 5399 3082 5846
rect 4880 5427 4997 5827
rect 5472 5429 5589 5829
rect 1078 33 1263 180
rect 1942 31 2127 178
rect 2709 50 2894 176
rect 2709 29 2898 50
rect 2874 11 2898 29
rect 5038 -5 5155 194
rect 5541 -7 5658 192
<< locali >>
rect 406 10928 480 10961
rect 375 10827 562 10928
rect 2578 10843 5387 10913
rect 6368 10854 6646 10863
rect 6368 10834 6662 10854
rect 406 10797 480 10827
rect 6365 10744 6662 10834
rect 6365 10730 6646 10744
rect 6365 10620 6420 10730
rect 504 5107 604 6351
rect 6328 6026 6413 6076
rect 3589 5956 6413 6026
rect 2582 5154 5391 5224
rect 6328 4992 6413 5956
rect 504 -252 604 992
rect 3593 290 4484 417
rect 2559 -131 5383 -50
rect 2583 -439 2619 -306
rect 6324 -455 6405 471
rect 3574 -4011 6398 -3930
use nmos101024  nmos101024_0
timestamp 1634049309
transform 1 0 4283 0 1 -4177
box -582 -119 2337 4276
use nmos101025  nmos101025_1
timestamp 1634049374
transform 1 0 4299 0 1 178
box -505 -81 2337 5316
use nmos101025  nmos101025_0
timestamp 1634049374
transform 1 0 4314 0 1 5817
box -505 -81 2337 5316
use nmos101035  nmos101035_0 ~/layout test
timestamp 1634045183
transform 1 0 717 0 1 585
box -717 -585 3227 5050
use nmos101035  nmos101035_1
timestamp 1634045183
transform 1 0 715 0 1 6250
box -717 -585 3227 5050
use nmos101043  nmos101043_0 ~/layout test
timestamp 1634046259
transform 1 0 527 0 1 -4144
box -531 0 3116 4190
<< labels >>
flabel poly 4007 11205 4007 11205 0 FreeSans 800 0 0 0 g
flabel locali 421 10856 421 10856 0 FreeSans 800 0 0 0 d
flabel locali 6458 10789 6458 10789 0 FreeSans 800 0 0 0 s
<< end >>
