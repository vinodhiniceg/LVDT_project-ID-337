magic
tech sky130A
magscale 1 2
timestamp 1634272774
<< error_p >>
rect -1411 362 1411 366
rect -1411 -362 -1381 362
rect -1345 296 1345 300
rect -1345 -296 -1315 296
rect 1315 -296 1345 296
rect -1345 -300 1345 -296
rect 1381 -362 1411 362
rect -1411 -366 1411 -362
<< nwell >>
rect -1381 -362 1381 362
<< mvpmos >>
rect -1287 -300 -687 300
rect -629 -300 -29 300
rect 29 -300 629 300
rect 687 -300 1287 300
<< mvpdiff >>
rect -1345 86 -1287 300
rect -1345 -86 -1333 86
rect -1299 -86 -1287 86
rect -1345 -300 -1287 -86
rect -687 86 -629 300
rect -687 -86 -675 86
rect -641 -86 -629 86
rect -687 -300 -629 -86
rect -29 86 29 300
rect -29 -86 -17 86
rect 17 -86 29 86
rect -29 -300 29 -86
rect 629 86 687 300
rect 629 -86 641 86
rect 675 -86 687 86
rect 629 -300 687 -86
rect 1287 86 1345 300
rect 1287 -86 1299 86
rect 1333 -86 1345 86
rect 1287 -300 1345 -86
<< mvpdiffc >>
rect -1333 -86 -1299 86
rect -675 -86 -641 86
rect -17 -86 17 86
rect 641 -86 675 86
rect 1299 -86 1333 86
<< poly >>
rect -1287 300 -687 326
rect -629 300 -29 326
rect 29 300 629 326
rect 687 300 1287 326
rect -1287 -326 -687 -300
rect -629 -326 -29 -300
rect 29 -326 629 -300
rect 687 -326 1287 -300
<< locali >>
rect -1333 86 -1299 102
rect -1333 -102 -1299 -86
rect -675 86 -641 102
rect -675 -102 -641 -86
rect -17 86 17 102
rect -17 -102 17 -86
rect 641 86 675 102
rect 641 -102 675 -86
rect 1299 86 1333 102
rect 1299 -102 1333 -86
<< viali >>
rect -1333 -86 -1299 86
rect -675 -86 -641 86
rect -17 -86 17 86
rect 641 -86 675 86
rect 1299 -86 1333 86
<< metal1 >>
rect -1339 86 -1293 98
rect -1339 -86 -1333 86
rect -1299 -86 -1293 86
rect -1339 -98 -1293 -86
rect -681 86 -635 98
rect -681 -86 -675 86
rect -641 -86 -635 86
rect -681 -98 -635 -86
rect -23 86 23 98
rect -23 -86 -17 86
rect 17 -86 23 86
rect -23 -98 23 -86
rect 635 86 681 98
rect 635 -86 641 86
rect 675 -86 681 86
rect 635 -98 681 -86
rect 1293 86 1339 98
rect 1293 -86 1299 86
rect 1333 -86 1339 86
rect 1293 -98 1339 -86
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string parameters w 3 l 3 m 1 nf 4 diffcov 30 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 30 viadrn 30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
