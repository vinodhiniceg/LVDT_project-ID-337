magic
tech sky130A
magscale 1 2
timestamp 1634904592
<< nwell >>
rect -487 -914 487 914
<< mvpmos >>
rect -229 488 -29 688
rect 29 488 229 688
rect -229 194 -29 394
rect 29 194 229 394
rect -229 -100 -29 100
rect 29 -100 229 100
rect -229 -394 -29 -194
rect 29 -394 229 -194
rect -229 -688 -29 -488
rect 29 -688 229 -488
<< mvpdiff >>
rect -287 614 -229 688
rect -287 562 -275 614
rect -241 562 -229 614
rect -287 488 -229 562
rect -29 614 29 688
rect -29 562 -17 614
rect 17 562 29 614
rect -29 488 29 562
rect 229 614 287 688
rect 229 562 241 614
rect 275 562 287 614
rect 229 488 287 562
rect -287 320 -229 394
rect -287 268 -275 320
rect -241 268 -229 320
rect -287 194 -229 268
rect -29 320 29 394
rect -29 268 -17 320
rect 17 268 29 320
rect -29 194 29 268
rect 229 320 287 394
rect 229 268 241 320
rect 275 268 287 320
rect 229 194 287 268
rect -287 26 -229 100
rect -287 -26 -275 26
rect -241 -26 -229 26
rect -287 -100 -229 -26
rect -29 26 29 100
rect -29 -26 -17 26
rect 17 -26 29 26
rect -29 -100 29 -26
rect 229 26 287 100
rect 229 -26 241 26
rect 275 -26 287 26
rect 229 -100 287 -26
rect -287 -268 -229 -194
rect -287 -320 -275 -268
rect -241 -320 -229 -268
rect -287 -394 -229 -320
rect -29 -268 29 -194
rect -29 -320 -17 -268
rect 17 -320 29 -268
rect -29 -394 29 -320
rect 229 -268 287 -194
rect 229 -320 241 -268
rect 275 -320 287 -268
rect 229 -394 287 -320
rect -287 -562 -229 -488
rect -287 -614 -275 -562
rect -241 -614 -229 -562
rect -287 -688 -229 -614
rect -29 -562 29 -488
rect -29 -614 -17 -562
rect 17 -614 29 -562
rect -29 -688 29 -614
rect 229 -562 287 -488
rect 229 -614 241 -562
rect 275 -614 287 -562
rect 229 -688 287 -614
<< mvpdiffc >>
rect -275 562 -241 614
rect -17 562 17 614
rect 241 562 275 614
rect -275 268 -241 320
rect -17 268 17 320
rect 241 268 275 320
rect -275 -26 -241 26
rect -17 -26 17 26
rect 241 -26 275 26
rect -275 -320 -241 -268
rect -17 -320 17 -268
rect 241 -320 275 -268
rect -275 -614 -241 -562
rect -17 -614 17 -562
rect 241 -614 275 -562
<< mvnsubdiff >>
rect -421 790 421 848
rect -421 222 -363 790
rect -421 -222 -409 222
rect -375 -222 -363 222
rect 363 222 421 790
rect -421 -790 -363 -222
rect 363 -222 375 222
rect 409 -222 421 222
rect 363 -790 421 -222
rect -421 -848 421 -790
<< mvnsubdiffcont >>
rect -409 -222 -375 222
rect 375 -222 409 222
<< poly >>
rect -229 688 -29 714
rect 29 688 229 714
rect -229 462 -29 488
rect 29 462 229 488
rect -229 394 -29 420
rect 29 394 229 420
rect -229 168 -29 194
rect 29 168 229 194
rect -229 100 -29 126
rect 29 100 229 126
rect -229 -126 -29 -100
rect 29 -126 229 -100
rect -229 -194 -29 -168
rect 29 -194 229 -168
rect -229 -420 -29 -394
rect 29 -420 229 -394
rect -229 -488 -29 -462
rect 29 -488 229 -462
rect -229 -714 -29 -688
rect 29 -714 229 -688
<< locali >>
rect -275 614 -241 630
rect -275 546 -241 562
rect -17 614 17 630
rect -17 546 17 562
rect 241 614 275 630
rect 241 546 275 562
rect -275 320 -241 336
rect -275 252 -241 268
rect -17 320 17 336
rect -17 252 17 268
rect 241 320 275 336
rect 241 252 275 268
rect -409 222 -375 238
rect 375 222 409 238
rect -275 26 -241 42
rect -275 -42 -241 -26
rect -17 26 17 42
rect -17 -42 17 -26
rect 241 26 275 42
rect 241 -42 275 -26
rect -409 -238 -375 -222
rect 375 -238 409 -222
rect -275 -268 -241 -252
rect -275 -336 -241 -320
rect -17 -268 17 -252
rect -17 -336 17 -320
rect 241 -268 275 -252
rect 241 -336 275 -320
rect -275 -562 -241 -546
rect -275 -630 -241 -614
rect -17 -562 17 -546
rect -17 -630 17 -614
rect 241 -562 275 -546
rect 241 -630 275 -614
<< viali >>
rect -275 562 -241 614
rect -17 562 17 614
rect 241 562 275 614
rect -275 268 -241 320
rect -17 268 17 320
rect 241 268 275 320
rect -275 -26 -241 26
rect -17 -26 17 26
rect 241 -26 275 26
rect -275 -320 -241 -268
rect -17 -320 17 -268
rect 241 -320 275 -268
rect -275 -614 -241 -562
rect -17 -614 17 -562
rect 241 -614 275 -562
<< metal1 >>
rect -281 614 -235 626
rect -281 562 -275 614
rect -241 562 -235 614
rect -281 550 -235 562
rect -23 614 23 626
rect -23 562 -17 614
rect 17 562 23 614
rect -23 550 23 562
rect 235 614 281 626
rect 235 562 241 614
rect 275 562 281 614
rect 235 550 281 562
rect -281 320 -235 332
rect -281 268 -275 320
rect -241 268 -235 320
rect -281 256 -235 268
rect -23 320 23 332
rect -23 268 -17 320
rect 17 268 23 320
rect -23 256 23 268
rect 235 320 281 332
rect 235 268 241 320
rect 275 268 281 320
rect 235 256 281 268
rect -281 26 -235 38
rect -281 -26 -275 26
rect -241 -26 -235 26
rect -281 -38 -235 -26
rect -23 26 23 38
rect -23 -26 -17 26
rect 17 -26 23 26
rect -23 -38 23 -26
rect 235 26 281 38
rect 235 -26 241 26
rect 275 -26 281 26
rect 235 -38 281 -26
rect -281 -268 -235 -256
rect -281 -320 -275 -268
rect -241 -320 -235 -268
rect -281 -332 -235 -320
rect -23 -268 23 -256
rect -23 -320 -17 -268
rect 17 -320 23 -268
rect -23 -332 23 -320
rect 235 -268 281 -256
rect 235 -320 241 -268
rect 275 -320 281 -268
rect 235 -332 281 -320
rect -281 -562 -235 -550
rect -281 -614 -275 -562
rect -241 -614 -235 -562
rect -281 -626 -235 -614
rect -23 -562 23 -550
rect -23 -614 -17 -562
rect 17 -614 23 -562
rect -23 -626 23 -614
rect 235 -562 281 -550
rect 235 -614 241 -562
rect 275 -614 281 -562
rect 235 -626 281 -614
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string FIXED_BBOX -392 -819 392 819
string parameters w 1 l 1 m 5 nf 2 diffcov 30 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 30 rlcov 30 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 30 viadrn 30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
