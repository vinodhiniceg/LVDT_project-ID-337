magic
tech sky130A
magscale 1 2
timestamp 1634112475
<< mvnmos >>
rect -629 2823 -29 3423
rect 29 2823 629 3423
rect -629 2129 -29 2729
rect 29 2129 629 2729
rect -629 1435 -29 2035
rect 29 1435 629 2035
rect -629 741 -29 1341
rect 29 741 629 1341
rect -629 47 -29 647
rect 29 47 629 647
rect -629 -647 -29 -47
rect 29 -647 629 -47
rect -629 -1341 -29 -741
rect 29 -1341 629 -741
rect -629 -2035 -29 -1435
rect 29 -2035 629 -1435
rect -629 -2729 -29 -2129
rect 29 -2729 629 -2129
rect -629 -3423 -29 -2823
rect 29 -3423 629 -2823
<< mvndiff >>
rect -687 3209 -629 3423
rect -687 3037 -675 3209
rect -641 3037 -629 3209
rect -687 2823 -629 3037
rect -29 3209 29 3423
rect -29 3037 -17 3209
rect 17 3037 29 3209
rect -29 2823 29 3037
rect 629 3209 687 3423
rect 629 3037 641 3209
rect 675 3037 687 3209
rect 629 2823 687 3037
rect -687 2515 -629 2729
rect -687 2343 -675 2515
rect -641 2343 -629 2515
rect -687 2129 -629 2343
rect -29 2515 29 2729
rect -29 2343 -17 2515
rect 17 2343 29 2515
rect -29 2129 29 2343
rect 629 2515 687 2729
rect 629 2343 641 2515
rect 675 2343 687 2515
rect 629 2129 687 2343
rect -687 1821 -629 2035
rect -687 1649 -675 1821
rect -641 1649 -629 1821
rect -687 1435 -629 1649
rect -29 1821 29 2035
rect -29 1649 -17 1821
rect 17 1649 29 1821
rect -29 1435 29 1649
rect 629 1821 687 2035
rect 629 1649 641 1821
rect 675 1649 687 1821
rect 629 1435 687 1649
rect -687 1127 -629 1341
rect -687 955 -675 1127
rect -641 955 -629 1127
rect -687 741 -629 955
rect -29 1127 29 1341
rect -29 955 -17 1127
rect 17 955 29 1127
rect -29 741 29 955
rect 629 1127 687 1341
rect 629 955 641 1127
rect 675 955 687 1127
rect 629 741 687 955
rect -687 433 -629 647
rect -687 261 -675 433
rect -641 261 -629 433
rect -687 47 -629 261
rect -29 433 29 647
rect -29 261 -17 433
rect 17 261 29 433
rect -29 47 29 261
rect 629 433 687 647
rect 629 261 641 433
rect 675 261 687 433
rect 629 47 687 261
rect -687 -261 -629 -47
rect -687 -433 -675 -261
rect -641 -433 -629 -261
rect -687 -647 -629 -433
rect -29 -261 29 -47
rect -29 -433 -17 -261
rect 17 -433 29 -261
rect -29 -647 29 -433
rect 629 -261 687 -47
rect 629 -433 641 -261
rect 675 -433 687 -261
rect 629 -647 687 -433
rect -687 -955 -629 -741
rect -687 -1127 -675 -955
rect -641 -1127 -629 -955
rect -687 -1341 -629 -1127
rect -29 -955 29 -741
rect -29 -1127 -17 -955
rect 17 -1127 29 -955
rect -29 -1341 29 -1127
rect 629 -955 687 -741
rect 629 -1127 641 -955
rect 675 -1127 687 -955
rect 629 -1341 687 -1127
rect -687 -1649 -629 -1435
rect -687 -1821 -675 -1649
rect -641 -1821 -629 -1649
rect -687 -2035 -629 -1821
rect -29 -1649 29 -1435
rect -29 -1821 -17 -1649
rect 17 -1821 29 -1649
rect -29 -2035 29 -1821
rect 629 -1649 687 -1435
rect 629 -1821 641 -1649
rect 675 -1821 687 -1649
rect 629 -2035 687 -1821
rect -687 -2343 -629 -2129
rect -687 -2515 -675 -2343
rect -641 -2515 -629 -2343
rect -687 -2729 -629 -2515
rect -29 -2343 29 -2129
rect -29 -2515 -17 -2343
rect 17 -2515 29 -2343
rect -29 -2729 29 -2515
rect 629 -2343 687 -2129
rect 629 -2515 641 -2343
rect 675 -2515 687 -2343
rect 629 -2729 687 -2515
rect -687 -3037 -629 -2823
rect -687 -3209 -675 -3037
rect -641 -3209 -629 -3037
rect -687 -3423 -629 -3209
rect -29 -3037 29 -2823
rect -29 -3209 -17 -3037
rect 17 -3209 29 -3037
rect -29 -3423 29 -3209
rect 629 -3037 687 -2823
rect 629 -3209 641 -3037
rect 675 -3209 687 -3037
rect 629 -3423 687 -3209
<< mvndiffc >>
rect -675 3037 -641 3209
rect -17 3037 17 3209
rect 641 3037 675 3209
rect -675 2343 -641 2515
rect -17 2343 17 2515
rect 641 2343 675 2515
rect -675 1649 -641 1821
rect -17 1649 17 1821
rect 641 1649 675 1821
rect -675 955 -641 1127
rect -17 955 17 1127
rect 641 955 675 1127
rect -675 261 -641 433
rect -17 261 17 433
rect 641 261 675 433
rect -675 -433 -641 -261
rect -17 -433 17 -261
rect 641 -433 675 -261
rect -675 -1127 -641 -955
rect -17 -1127 17 -955
rect 641 -1127 675 -955
rect -675 -1821 -641 -1649
rect -17 -1821 17 -1649
rect 641 -1821 675 -1649
rect -675 -2515 -641 -2343
rect -17 -2515 17 -2343
rect 641 -2515 675 -2343
rect -675 -3209 -641 -3037
rect -17 -3209 17 -3037
rect 641 -3209 675 -3037
<< poly >>
rect -629 3423 -29 3449
rect 29 3423 629 3449
rect -629 2797 -29 2823
rect 29 2797 629 2823
rect -629 2729 -29 2755
rect 29 2729 629 2755
rect -629 2103 -29 2129
rect 29 2103 629 2129
rect -629 2035 -29 2061
rect 29 2035 629 2061
rect -629 1409 -29 1435
rect 29 1409 629 1435
rect -629 1341 -29 1367
rect 29 1341 629 1367
rect -629 715 -29 741
rect 29 715 629 741
rect -629 647 -29 673
rect 29 647 629 673
rect -629 21 -29 47
rect 29 21 629 47
rect -629 -47 -29 -21
rect 29 -47 629 -21
rect -629 -673 -29 -647
rect 29 -673 629 -647
rect -629 -741 -29 -715
rect 29 -741 629 -715
rect -629 -1367 -29 -1341
rect 29 -1367 629 -1341
rect -629 -1435 -29 -1409
rect 29 -1435 629 -1409
rect -629 -2061 -29 -2035
rect 29 -2061 629 -2035
rect -629 -2129 -29 -2103
rect 29 -2129 629 -2103
rect -629 -2755 -29 -2729
rect 29 -2755 629 -2729
rect -629 -2823 -29 -2797
rect 29 -2823 629 -2797
rect -629 -3449 -29 -3423
rect 29 -3449 629 -3423
<< locali >>
rect -675 3209 -641 3225
rect -675 3021 -641 3037
rect -17 3209 17 3225
rect -17 3021 17 3037
rect 641 3209 675 3225
rect 641 3021 675 3037
rect -675 2515 -641 2531
rect -675 2327 -641 2343
rect -17 2515 17 2531
rect -17 2327 17 2343
rect 641 2515 675 2531
rect 641 2327 675 2343
rect -675 1821 -641 1837
rect -675 1633 -641 1649
rect -17 1821 17 1837
rect -17 1633 17 1649
rect 641 1821 675 1837
rect 641 1633 675 1649
rect -675 1127 -641 1143
rect -675 939 -641 955
rect -17 1127 17 1143
rect -17 939 17 955
rect 641 1127 675 1143
rect 641 939 675 955
rect -675 433 -641 449
rect -675 245 -641 261
rect -17 433 17 449
rect -17 245 17 261
rect 641 433 675 449
rect 641 245 675 261
rect -675 -261 -641 -245
rect -675 -449 -641 -433
rect -17 -261 17 -245
rect -17 -449 17 -433
rect 641 -261 675 -245
rect 641 -449 675 -433
rect -675 -955 -641 -939
rect -675 -1143 -641 -1127
rect -17 -955 17 -939
rect -17 -1143 17 -1127
rect 641 -955 675 -939
rect 641 -1143 675 -1127
rect -675 -1649 -641 -1633
rect -675 -1837 -641 -1821
rect -17 -1649 17 -1633
rect -17 -1837 17 -1821
rect 641 -1649 675 -1633
rect 641 -1837 675 -1821
rect -675 -2343 -641 -2327
rect -675 -2531 -641 -2515
rect -17 -2343 17 -2327
rect -17 -2531 17 -2515
rect 641 -2343 675 -2327
rect 641 -2531 675 -2515
rect -675 -3037 -641 -3021
rect -675 -3225 -641 -3209
rect -17 -3037 17 -3021
rect -17 -3225 17 -3209
rect 641 -3037 675 -3021
rect 641 -3225 675 -3209
<< viali >>
rect -675 3037 -641 3209
rect -17 3037 17 3209
rect 641 3037 675 3209
rect -675 2343 -641 2515
rect -17 2343 17 2515
rect 641 2343 675 2515
rect -675 1649 -641 1821
rect -17 1649 17 1821
rect 641 1649 675 1821
rect -675 955 -641 1127
rect -17 955 17 1127
rect 641 955 675 1127
rect -675 261 -641 433
rect -17 261 17 433
rect 641 261 675 433
rect -675 -433 -641 -261
rect -17 -433 17 -261
rect 641 -433 675 -261
rect -675 -1127 -641 -955
rect -17 -1127 17 -955
rect 641 -1127 675 -955
rect -675 -1821 -641 -1649
rect -17 -1821 17 -1649
rect 641 -1821 675 -1649
rect -675 -2515 -641 -2343
rect -17 -2515 17 -2343
rect 641 -2515 675 -2343
rect -675 -3209 -641 -3037
rect -17 -3209 17 -3037
rect 641 -3209 675 -3037
<< metal1 >>
rect -681 3209 -635 3221
rect -681 3037 -675 3209
rect -641 3037 -635 3209
rect -681 3025 -635 3037
rect -23 3209 23 3221
rect -23 3037 -17 3209
rect 17 3037 23 3209
rect -23 3025 23 3037
rect 635 3209 681 3221
rect 635 3037 641 3209
rect 675 3037 681 3209
rect 635 3025 681 3037
rect -681 2515 -635 2527
rect -681 2343 -675 2515
rect -641 2343 -635 2515
rect -681 2331 -635 2343
rect -23 2515 23 2527
rect -23 2343 -17 2515
rect 17 2343 23 2515
rect -23 2331 23 2343
rect 635 2515 681 2527
rect 635 2343 641 2515
rect 675 2343 681 2515
rect 635 2331 681 2343
rect -681 1821 -635 1833
rect -681 1649 -675 1821
rect -641 1649 -635 1821
rect -681 1637 -635 1649
rect -23 1821 23 1833
rect -23 1649 -17 1821
rect 17 1649 23 1821
rect -23 1637 23 1649
rect 635 1821 681 1833
rect 635 1649 641 1821
rect 675 1649 681 1821
rect 635 1637 681 1649
rect -681 1127 -635 1139
rect -681 955 -675 1127
rect -641 955 -635 1127
rect -681 943 -635 955
rect -23 1127 23 1139
rect -23 955 -17 1127
rect 17 955 23 1127
rect -23 943 23 955
rect 635 1127 681 1139
rect 635 955 641 1127
rect 675 955 681 1127
rect 635 943 681 955
rect -681 433 -635 445
rect -681 261 -675 433
rect -641 261 -635 433
rect -681 249 -635 261
rect -23 433 23 445
rect -23 261 -17 433
rect 17 261 23 433
rect -23 249 23 261
rect 635 433 681 445
rect 635 261 641 433
rect 675 261 681 433
rect 635 249 681 261
rect -681 -261 -635 -249
rect -681 -433 -675 -261
rect -641 -433 -635 -261
rect -681 -445 -635 -433
rect -23 -261 23 -249
rect -23 -433 -17 -261
rect 17 -433 23 -261
rect -23 -445 23 -433
rect 635 -261 681 -249
rect 635 -433 641 -261
rect 675 -433 681 -261
rect 635 -445 681 -433
rect -681 -955 -635 -943
rect -681 -1127 -675 -955
rect -641 -1127 -635 -955
rect -681 -1139 -635 -1127
rect -23 -955 23 -943
rect -23 -1127 -17 -955
rect 17 -1127 23 -955
rect -23 -1139 23 -1127
rect 635 -955 681 -943
rect 635 -1127 641 -955
rect 675 -1127 681 -955
rect 635 -1139 681 -1127
rect -681 -1649 -635 -1637
rect -681 -1821 -675 -1649
rect -641 -1821 -635 -1649
rect -681 -1833 -635 -1821
rect -23 -1649 23 -1637
rect -23 -1821 -17 -1649
rect 17 -1821 23 -1649
rect -23 -1833 23 -1821
rect 635 -1649 681 -1637
rect 635 -1821 641 -1649
rect 675 -1821 681 -1649
rect 635 -1833 681 -1821
rect -681 -2343 -635 -2331
rect -681 -2515 -675 -2343
rect -641 -2515 -635 -2343
rect -681 -2527 -635 -2515
rect -23 -2343 23 -2331
rect -23 -2515 -17 -2343
rect 17 -2515 23 -2343
rect -23 -2527 23 -2515
rect 635 -2343 681 -2331
rect 635 -2515 641 -2343
rect 675 -2515 681 -2343
rect 635 -2527 681 -2515
rect -681 -3037 -635 -3025
rect -681 -3209 -675 -3037
rect -641 -3209 -635 -3037
rect -681 -3221 -635 -3209
rect -23 -3037 23 -3025
rect -23 -3209 -17 -3037
rect 17 -3209 23 -3037
rect -23 -3221 23 -3209
rect 635 -3037 681 -3025
rect 635 -3209 641 -3037
rect 675 -3209 681 -3037
rect 635 -3221 681 -3209
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string parameters w 3 l 3 m 10 nf 2 diffcov 30 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 30 viadrn 30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
