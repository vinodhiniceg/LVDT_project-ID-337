magic
tech sky130A
magscale 1 2
timestamp 1634564603
<< nwell >>
rect 70542 75224 82208 75552
rect 70542 75030 82222 75224
rect 70572 74254 82222 75030
rect 62 60088 21214 66356
rect 41674 65392 58346 74064
rect 70594 73624 82222 74254
rect 70594 73578 82226 73624
rect 34 59490 21214 60088
rect 41654 64462 58346 65392
rect 34 46856 21186 59490
rect 41654 56804 58326 64462
rect 41598 55790 58326 56804
rect 41598 47202 58270 55790
rect 70596 50894 82226 73578
rect 83206 53645 86410 54165
rect 70558 50824 82226 50894
rect 70558 49684 82222 50824
<< pwell >>
rect 30576 58170 30928 58184
rect 22890 51718 30928 58170
rect 22890 51704 30900 51718
rect 23066 51690 30900 51704
rect 83726 53485 85246 53551
rect 85895 53485 86340 53585
rect 83276 53311 86340 53485
rect 83246 53225 86370 53311
rect 0 45406 60208 45432
rect 0 44094 60238 45406
rect 48 8660 60238 44094
rect 61936 39382 74230 43948
rect 76540 40024 87260 40040
rect 76436 39788 87260 40024
rect 76436 39580 87274 39788
rect 62064 39342 73904 39382
rect 76460 34664 87274 39580
rect 60858 27536 61940 27564
rect 99996 27536 101526 27564
rect 60858 27000 101526 27536
rect 48 8546 21928 8660
rect 26402 8546 60238 8660
rect 48 1284 60238 8546
rect 60534 1904 101526 27000
rect 60908 1868 101526 1904
rect 60908 1844 101434 1868
rect 48 30 60292 1284
rect 59558 0 60238 30
<< mvnmos >>
rect 23420 56834 24020 57434
rect 24114 56834 24714 57434
rect 24808 56834 25408 57434
rect 25502 56834 26102 57434
rect 26196 56834 26796 57434
rect 26890 56834 27490 57434
rect 27584 56834 28184 57434
rect 28278 56834 28878 57434
rect 28972 56834 29572 57434
rect 29666 56834 30266 57434
rect 23420 56176 24020 56776
rect 24114 56176 24714 56776
rect 24808 56176 25408 56776
rect 25502 56176 26102 56776
rect 26196 56176 26796 56776
rect 26890 56176 27490 56776
rect 27584 56176 28184 56776
rect 28278 56176 28878 56776
rect 28972 56176 29572 56776
rect 29666 56176 30266 56776
rect 23426 54944 24026 55544
rect 24120 54944 24720 55544
rect 24814 54944 25414 55544
rect 25508 54944 26108 55544
rect 26202 54944 26802 55544
rect 26896 54944 27496 55544
rect 27590 54944 28190 55544
rect 28284 54944 28884 55544
rect 28978 54944 29578 55544
rect 29672 54944 30272 55544
rect 23426 54286 24026 54886
rect 24120 54286 24720 54886
rect 24814 54286 25414 54886
rect 25508 54286 26108 54886
rect 26202 54286 26802 54886
rect 26896 54286 27496 54886
rect 27590 54286 28190 54886
rect 28284 54286 28884 54886
rect 28978 54286 29578 54886
rect 29672 54286 30272 54886
rect 23442 53002 24042 53602
rect 24136 53002 24736 53602
rect 24830 53002 25430 53602
rect 25524 53002 26124 53602
rect 26218 53002 26818 53602
rect 26912 53002 27512 53602
rect 27606 53002 28206 53602
rect 28300 53002 28900 53602
rect 28994 53002 29594 53602
rect 29688 53002 30288 53602
rect 23442 52344 24042 52944
rect 24136 52344 24736 52944
rect 24830 52344 25430 52944
rect 25524 52344 26124 52944
rect 26218 52344 26818 52944
rect 26912 52344 27512 52944
rect 27606 52344 28206 52944
rect 28300 52344 28900 52944
rect 28994 52344 29594 52944
rect 29688 52344 30288 52944
rect 83359 53375 83459 53459
rect 83515 53375 83615 53459
rect 83809 53441 83909 53525
rect 83951 53441 84051 53525
rect 84107 53441 84207 53525
rect 84263 53441 84363 53525
rect 84405 53441 84505 53525
rect 84552 53441 84652 53525
rect 84905 53375 85005 53525
rect 85061 53375 85161 53525
rect 85978 53475 86078 53559
rect 85261 53375 85361 53459
rect 85403 53375 85503 53459
rect 85559 53375 85659 53459
rect 85701 53375 85801 53459
rect 86157 53409 86257 53559
rect 2004 42406 3004 43406
rect 3062 42406 4062 43406
rect 4120 42406 5120 43406
rect 5178 42406 6178 43406
rect 6236 42406 7236 43406
rect 8518 42414 9518 43414
rect 9576 42414 10576 43414
rect 10634 42414 11634 43414
rect 11692 42414 12692 43414
rect 12750 42414 13750 43414
rect 15024 42422 16024 43422
rect 16082 42422 17082 43422
rect 17140 42422 18140 43422
rect 18198 42422 19198 43422
rect 19256 42422 20256 43422
rect 21514 42406 22514 43406
rect 22572 42406 23572 43406
rect 23630 42406 24630 43406
rect 24688 42406 25688 43406
rect 25746 42406 26746 43406
rect 28036 42422 29036 43422
rect 29094 42422 30094 43422
rect 30152 42422 31152 43422
rect 31210 42422 32210 43422
rect 32268 42422 33268 43422
rect 34546 42428 35546 43428
rect 35604 42428 36604 43428
rect 36662 42428 37662 43428
rect 37720 42428 38720 43428
rect 38778 42428 39778 43428
rect 41036 42428 42036 43428
rect 42094 42428 43094 43428
rect 43152 42428 44152 43428
rect 44210 42428 45210 43428
rect 45268 42428 46268 43428
rect 47624 42450 48624 43450
rect 48682 42450 49682 43450
rect 49740 42450 50740 43450
rect 50798 42450 51798 43450
rect 51856 42450 52856 43450
rect 54138 42464 55138 43464
rect 55196 42464 56196 43464
rect 56254 42464 57254 43464
rect 57312 42464 58312 43464
rect 58370 42464 59370 43464
rect 2004 41312 3004 42312
rect 3062 41312 4062 42312
rect 4120 41312 5120 42312
rect 5178 41312 6178 42312
rect 6236 41312 7236 42312
rect 2004 40218 3004 41218
rect 3062 40218 4062 41218
rect 4120 40218 5120 41218
rect 5178 40218 6178 41218
rect 6236 40218 7236 41218
rect 8518 41320 9518 42320
rect 9576 41320 10576 42320
rect 10634 41320 11634 42320
rect 11692 41320 12692 42320
rect 12750 41320 13750 42320
rect 2004 39124 3004 40124
rect 3062 39124 4062 40124
rect 4120 39124 5120 40124
rect 5178 39124 6178 40124
rect 6236 39124 7236 40124
rect 8518 40226 9518 41226
rect 9576 40226 10576 41226
rect 10634 40226 11634 41226
rect 11692 40226 12692 41226
rect 12750 40226 13750 41226
rect 15024 41328 16024 42328
rect 16082 41328 17082 42328
rect 17140 41328 18140 42328
rect 18198 41328 19198 42328
rect 19256 41328 20256 42328
rect 8518 39132 9518 40132
rect 9576 39132 10576 40132
rect 10634 39132 11634 40132
rect 11692 39132 12692 40132
rect 12750 39132 13750 40132
rect 15024 40234 16024 41234
rect 16082 40234 17082 41234
rect 17140 40234 18140 41234
rect 18198 40234 19198 41234
rect 19256 40234 20256 41234
rect 21514 41312 22514 42312
rect 22572 41312 23572 42312
rect 23630 41312 24630 42312
rect 24688 41312 25688 42312
rect 25746 41312 26746 42312
rect 15024 39140 16024 40140
rect 16082 39140 17082 40140
rect 17140 39140 18140 40140
rect 18198 39140 19198 40140
rect 19256 39140 20256 40140
rect 21514 40218 22514 41218
rect 22572 40218 23572 41218
rect 23630 40218 24630 41218
rect 24688 40218 25688 41218
rect 25746 40218 26746 41218
rect 28036 41328 29036 42328
rect 29094 41328 30094 42328
rect 30152 41328 31152 42328
rect 31210 41328 32210 42328
rect 32268 41328 33268 42328
rect 21514 39124 22514 40124
rect 22572 39124 23572 40124
rect 23630 39124 24630 40124
rect 24688 39124 25688 40124
rect 25746 39124 26746 40124
rect 28036 40234 29036 41234
rect 29094 40234 30094 41234
rect 30152 40234 31152 41234
rect 31210 40234 32210 41234
rect 32268 40234 33268 41234
rect 34546 41334 35546 42334
rect 35604 41334 36604 42334
rect 36662 41334 37662 42334
rect 37720 41334 38720 42334
rect 38778 41334 39778 42334
rect 28036 39140 29036 40140
rect 29094 39140 30094 40140
rect 30152 39140 31152 40140
rect 31210 39140 32210 40140
rect 32268 39140 33268 40140
rect 34546 40240 35546 41240
rect 35604 40240 36604 41240
rect 36662 40240 37662 41240
rect 37720 40240 38720 41240
rect 38778 40240 39778 41240
rect 41036 41334 42036 42334
rect 42094 41334 43094 42334
rect 43152 41334 44152 42334
rect 44210 41334 45210 42334
rect 45268 41334 46268 42334
rect 34546 39146 35546 40146
rect 35604 39146 36604 40146
rect 36662 39146 37662 40146
rect 37720 39146 38720 40146
rect 38778 39146 39778 40146
rect 41036 40240 42036 41240
rect 42094 40240 43094 41240
rect 43152 40240 44152 41240
rect 44210 40240 45210 41240
rect 45268 40240 46268 41240
rect 47624 41356 48624 42356
rect 48682 41356 49682 42356
rect 49740 41356 50740 42356
rect 50798 41356 51798 42356
rect 51856 41356 52856 42356
rect 41036 39146 42036 40146
rect 42094 39146 43094 40146
rect 43152 39146 44152 40146
rect 44210 39146 45210 40146
rect 45268 39146 46268 40146
rect 47624 40262 48624 41262
rect 48682 40262 49682 41262
rect 49740 40262 50740 41262
rect 50798 40262 51798 41262
rect 51856 40262 52856 41262
rect 54138 41370 55138 42370
rect 55196 41370 56196 42370
rect 56254 41370 57254 42370
rect 57312 41370 58312 42370
rect 58370 41370 59370 42370
rect 47624 39168 48624 40168
rect 48682 39168 49682 40168
rect 49740 39168 50740 40168
rect 50798 39168 51798 40168
rect 51856 39168 52856 40168
rect 54138 40276 55138 41276
rect 55196 40276 56196 41276
rect 56254 40276 57254 41276
rect 57312 40276 58312 41276
rect 58370 40276 59370 41276
rect 54138 39182 55138 40182
rect 55196 39182 56196 40182
rect 56254 39182 57254 40182
rect 57312 39182 58312 40182
rect 58370 39182 59370 40182
rect 2004 38030 3004 39030
rect 3062 38030 4062 39030
rect 4120 38030 5120 39030
rect 5178 38030 6178 39030
rect 6236 38030 7236 39030
rect 8518 38038 9518 39038
rect 9576 38038 10576 39038
rect 10634 38038 11634 39038
rect 11692 38038 12692 39038
rect 12750 38038 13750 39038
rect 15024 38046 16024 39046
rect 16082 38046 17082 39046
rect 17140 38046 18140 39046
rect 18198 38046 19198 39046
rect 19256 38046 20256 39046
rect 21514 38030 22514 39030
rect 22572 38030 23572 39030
rect 23630 38030 24630 39030
rect 24688 38030 25688 39030
rect 25746 38030 26746 39030
rect 28036 38046 29036 39046
rect 29094 38046 30094 39046
rect 30152 38046 31152 39046
rect 31210 38046 32210 39046
rect 32268 38046 33268 39046
rect 34546 38052 35546 39052
rect 35604 38052 36604 39052
rect 36662 38052 37662 39052
rect 37720 38052 38720 39052
rect 38778 38052 39778 39052
rect 41036 38052 42036 39052
rect 42094 38052 43094 39052
rect 43152 38052 44152 39052
rect 44210 38052 45210 39052
rect 45268 38052 46268 39052
rect 47624 38074 48624 39074
rect 48682 38074 49682 39074
rect 49740 38074 50740 39074
rect 50798 38074 51798 39074
rect 51856 38074 52856 39074
rect 54138 38088 55138 39088
rect 55196 38088 56196 39088
rect 56254 38088 57254 39088
rect 57312 38088 58312 39088
rect 58370 38088 59370 39088
rect 2004 36590 3004 37590
rect 3062 36590 4062 37590
rect 4120 36590 5120 37590
rect 5178 36590 6178 37590
rect 6236 36590 7236 37590
rect 8518 36598 9518 37598
rect 9576 36598 10576 37598
rect 10634 36598 11634 37598
rect 11692 36598 12692 37598
rect 12750 36598 13750 37598
rect 15024 36606 16024 37606
rect 16082 36606 17082 37606
rect 17140 36606 18140 37606
rect 18198 36606 19198 37606
rect 19256 36606 20256 37606
rect 21514 36590 22514 37590
rect 22572 36590 23572 37590
rect 23630 36590 24630 37590
rect 24688 36590 25688 37590
rect 25746 36590 26746 37590
rect 28036 36606 29036 37606
rect 29094 36606 30094 37606
rect 30152 36606 31152 37606
rect 31210 36606 32210 37606
rect 32268 36606 33268 37606
rect 34546 36612 35546 37612
rect 35604 36612 36604 37612
rect 36662 36612 37662 37612
rect 37720 36612 38720 37612
rect 38778 36612 39778 37612
rect 41036 36612 42036 37612
rect 42094 36612 43094 37612
rect 43152 36612 44152 37612
rect 44210 36612 45210 37612
rect 45268 36612 46268 37612
rect 47624 36634 48624 37634
rect 48682 36634 49682 37634
rect 49740 36634 50740 37634
rect 50798 36634 51798 37634
rect 51856 36634 52856 37634
rect 54138 36648 55138 37648
rect 55196 36648 56196 37648
rect 56254 36648 57254 37648
rect 57312 36648 58312 37648
rect 58370 36648 59370 37648
rect 2004 35496 3004 36496
rect 3062 35496 4062 36496
rect 4120 35496 5120 36496
rect 5178 35496 6178 36496
rect 6236 35496 7236 36496
rect 2004 34402 3004 35402
rect 3062 34402 4062 35402
rect 4120 34402 5120 35402
rect 5178 34402 6178 35402
rect 6236 34402 7236 35402
rect 8518 35504 9518 36504
rect 9576 35504 10576 36504
rect 10634 35504 11634 36504
rect 11692 35504 12692 36504
rect 12750 35504 13750 36504
rect 2004 33308 3004 34308
rect 3062 33308 4062 34308
rect 4120 33308 5120 34308
rect 5178 33308 6178 34308
rect 6236 33308 7236 34308
rect 8518 34410 9518 35410
rect 9576 34410 10576 35410
rect 10634 34410 11634 35410
rect 11692 34410 12692 35410
rect 12750 34410 13750 35410
rect 15024 35512 16024 36512
rect 16082 35512 17082 36512
rect 17140 35512 18140 36512
rect 18198 35512 19198 36512
rect 19256 35512 20256 36512
rect 8518 33316 9518 34316
rect 9576 33316 10576 34316
rect 10634 33316 11634 34316
rect 11692 33316 12692 34316
rect 12750 33316 13750 34316
rect 15024 34418 16024 35418
rect 16082 34418 17082 35418
rect 17140 34418 18140 35418
rect 18198 34418 19198 35418
rect 19256 34418 20256 35418
rect 21514 35496 22514 36496
rect 22572 35496 23572 36496
rect 23630 35496 24630 36496
rect 24688 35496 25688 36496
rect 25746 35496 26746 36496
rect 15024 33324 16024 34324
rect 16082 33324 17082 34324
rect 17140 33324 18140 34324
rect 18198 33324 19198 34324
rect 19256 33324 20256 34324
rect 21514 34402 22514 35402
rect 22572 34402 23572 35402
rect 23630 34402 24630 35402
rect 24688 34402 25688 35402
rect 25746 34402 26746 35402
rect 28036 35512 29036 36512
rect 29094 35512 30094 36512
rect 30152 35512 31152 36512
rect 31210 35512 32210 36512
rect 32268 35512 33268 36512
rect 21514 33308 22514 34308
rect 22572 33308 23572 34308
rect 23630 33308 24630 34308
rect 24688 33308 25688 34308
rect 25746 33308 26746 34308
rect 28036 34418 29036 35418
rect 29094 34418 30094 35418
rect 30152 34418 31152 35418
rect 31210 34418 32210 35418
rect 32268 34418 33268 35418
rect 34546 35518 35546 36518
rect 35604 35518 36604 36518
rect 36662 35518 37662 36518
rect 37720 35518 38720 36518
rect 38778 35518 39778 36518
rect 28036 33324 29036 34324
rect 29094 33324 30094 34324
rect 30152 33324 31152 34324
rect 31210 33324 32210 34324
rect 32268 33324 33268 34324
rect 34546 34424 35546 35424
rect 35604 34424 36604 35424
rect 36662 34424 37662 35424
rect 37720 34424 38720 35424
rect 38778 34424 39778 35424
rect 41036 35518 42036 36518
rect 42094 35518 43094 36518
rect 43152 35518 44152 36518
rect 44210 35518 45210 36518
rect 45268 35518 46268 36518
rect 34546 33330 35546 34330
rect 35604 33330 36604 34330
rect 36662 33330 37662 34330
rect 37720 33330 38720 34330
rect 38778 33330 39778 34330
rect 41036 34424 42036 35424
rect 42094 34424 43094 35424
rect 43152 34424 44152 35424
rect 44210 34424 45210 35424
rect 45268 34424 46268 35424
rect 47624 35540 48624 36540
rect 48682 35540 49682 36540
rect 49740 35540 50740 36540
rect 50798 35540 51798 36540
rect 51856 35540 52856 36540
rect 41036 33330 42036 34330
rect 42094 33330 43094 34330
rect 43152 33330 44152 34330
rect 44210 33330 45210 34330
rect 45268 33330 46268 34330
rect 47624 34446 48624 35446
rect 48682 34446 49682 35446
rect 49740 34446 50740 35446
rect 50798 34446 51798 35446
rect 51856 34446 52856 35446
rect 54138 35554 55138 36554
rect 55196 35554 56196 36554
rect 56254 35554 57254 36554
rect 57312 35554 58312 36554
rect 58370 35554 59370 36554
rect 62554 42722 63154 43322
rect 63212 42722 63812 43322
rect 63870 42722 64470 43322
rect 64528 42722 65128 43322
rect 65186 42722 65786 43322
rect 66348 42724 66948 43324
rect 67006 42724 67606 43324
rect 67664 42724 68264 43324
rect 68322 42724 68922 43324
rect 68980 42724 69580 43324
rect 70156 42738 70756 43338
rect 70814 42738 71414 43338
rect 71472 42738 72072 43338
rect 72130 42738 72730 43338
rect 72788 42738 73388 43338
rect 62554 42028 63154 42628
rect 63212 42028 63812 42628
rect 63870 42028 64470 42628
rect 64528 42028 65128 42628
rect 65186 42028 65786 42628
rect 62554 41334 63154 41934
rect 63212 41334 63812 41934
rect 63870 41334 64470 41934
rect 64528 41334 65128 41934
rect 65186 41334 65786 41934
rect 62554 40640 63154 41240
rect 63212 40640 63812 41240
rect 63870 40640 64470 41240
rect 64528 40640 65128 41240
rect 65186 40640 65786 41240
rect 66348 42030 66948 42630
rect 67006 42030 67606 42630
rect 67664 42030 68264 42630
rect 68322 42030 68922 42630
rect 68980 42030 69580 42630
rect 66348 41336 66948 41936
rect 67006 41336 67606 41936
rect 67664 41336 68264 41936
rect 68322 41336 68922 41936
rect 68980 41336 69580 41936
rect 66348 40642 66948 41242
rect 67006 40642 67606 41242
rect 67664 40642 68264 41242
rect 68322 40642 68922 41242
rect 68980 40642 69580 41242
rect 70156 42044 70756 42644
rect 70814 42044 71414 42644
rect 71472 42044 72072 42644
rect 72130 42044 72730 42644
rect 72788 42044 73388 42644
rect 70156 41350 70756 41950
rect 70814 41350 71414 41950
rect 71472 41350 72072 41950
rect 72130 41350 72730 41950
rect 72788 41350 73388 41950
rect 70156 40656 70756 41256
rect 70814 40656 71414 41256
rect 71472 40656 72072 41256
rect 72130 40656 72730 41256
rect 72788 40656 73388 41256
rect 62554 39946 63154 40546
rect 63212 39946 63812 40546
rect 63870 39946 64470 40546
rect 64528 39946 65128 40546
rect 65186 39946 65786 40546
rect 66348 39948 66948 40548
rect 67006 39948 67606 40548
rect 67664 39948 68264 40548
rect 68322 39948 68922 40548
rect 68980 39948 69580 40548
rect 70156 39962 70756 40562
rect 70814 39962 71414 40562
rect 71472 39962 72072 40562
rect 72130 39962 72730 40562
rect 72788 39962 73388 40562
rect 47624 33352 48624 34352
rect 48682 33352 49682 34352
rect 49740 33352 50740 34352
rect 50798 33352 51798 34352
rect 51856 33352 52856 34352
rect 54138 34460 55138 35460
rect 55196 34460 56196 35460
rect 56254 34460 57254 35460
rect 57312 34460 58312 35460
rect 58370 34460 59370 35460
rect 77216 38708 77816 39308
rect 77874 38708 78474 39308
rect 78532 38708 79132 39308
rect 79190 38708 79790 39308
rect 77216 38014 77816 38614
rect 77874 38014 78474 38614
rect 78532 38014 79132 38614
rect 79190 38014 79790 38614
rect 77216 37320 77816 37920
rect 77874 37320 78474 37920
rect 78532 37320 79132 37920
rect 79190 37320 79790 37920
rect 77216 36626 77816 37226
rect 77874 36626 78474 37226
rect 78532 36626 79132 37226
rect 79190 36626 79790 37226
rect 77216 35932 77816 36532
rect 77874 35932 78474 36532
rect 78532 35932 79132 36532
rect 79190 35932 79790 36532
rect 77216 35238 77816 35838
rect 77874 35238 78474 35838
rect 78532 35238 79132 35838
rect 79190 35238 79790 35838
rect 80542 38702 81142 39302
rect 81200 38702 81800 39302
rect 81858 38702 82458 39302
rect 82516 38702 83116 39302
rect 80542 38008 81142 38608
rect 81200 38008 81800 38608
rect 81858 38008 82458 38608
rect 82516 38008 83116 38608
rect 80542 37314 81142 37914
rect 81200 37314 81800 37914
rect 81858 37314 82458 37914
rect 82516 37314 83116 37914
rect 80542 36620 81142 37220
rect 81200 36620 81800 37220
rect 81858 36620 82458 37220
rect 82516 36620 83116 37220
rect 80542 35926 81142 36526
rect 81200 35926 81800 36526
rect 81858 35926 82458 36526
rect 82516 35926 83116 36526
rect 80542 35232 81142 35832
rect 81200 35232 81800 35832
rect 81858 35232 82458 35832
rect 82516 35232 83116 35832
rect 83852 38702 84452 39302
rect 84510 38702 85110 39302
rect 85168 38702 85768 39302
rect 85826 38702 86426 39302
rect 83852 38008 84452 38608
rect 84510 38008 85110 38608
rect 85168 38008 85768 38608
rect 85826 38008 86426 38608
rect 83852 37314 84452 37914
rect 84510 37314 85110 37914
rect 85168 37314 85768 37914
rect 85826 37314 86426 37914
rect 83852 36620 84452 37220
rect 84510 36620 85110 37220
rect 85168 36620 85768 37220
rect 85826 36620 86426 37220
rect 83852 35926 84452 36526
rect 84510 35926 85110 36526
rect 85168 35926 85768 36526
rect 85826 35926 86426 36526
rect 83852 35232 84452 35832
rect 84510 35232 85110 35832
rect 85168 35232 85768 35832
rect 85826 35232 86426 35832
rect 54138 33366 55138 34366
rect 55196 33366 56196 34366
rect 56254 33366 57254 34366
rect 57312 33366 58312 34366
rect 58370 33366 59370 34366
rect 2004 32214 3004 33214
rect 3062 32214 4062 33214
rect 4120 32214 5120 33214
rect 5178 32214 6178 33214
rect 6236 32214 7236 33214
rect 8518 32222 9518 33222
rect 9576 32222 10576 33222
rect 10634 32222 11634 33222
rect 11692 32222 12692 33222
rect 12750 32222 13750 33222
rect 15024 32230 16024 33230
rect 16082 32230 17082 33230
rect 17140 32230 18140 33230
rect 18198 32230 19198 33230
rect 19256 32230 20256 33230
rect 21514 32214 22514 33214
rect 22572 32214 23572 33214
rect 23630 32214 24630 33214
rect 24688 32214 25688 33214
rect 25746 32214 26746 33214
rect 28036 32230 29036 33230
rect 29094 32230 30094 33230
rect 30152 32230 31152 33230
rect 31210 32230 32210 33230
rect 32268 32230 33268 33230
rect 34546 32236 35546 33236
rect 35604 32236 36604 33236
rect 36662 32236 37662 33236
rect 37720 32236 38720 33236
rect 38778 32236 39778 33236
rect 41036 32236 42036 33236
rect 42094 32236 43094 33236
rect 43152 32236 44152 33236
rect 44210 32236 45210 33236
rect 45268 32236 46268 33236
rect 47624 32258 48624 33258
rect 48682 32258 49682 33258
rect 49740 32258 50740 33258
rect 50798 32258 51798 33258
rect 51856 32258 52856 33258
rect 54138 32272 55138 33272
rect 55196 32272 56196 33272
rect 56254 32272 57254 33272
rect 57312 32272 58312 33272
rect 58370 32272 59370 33272
rect 2004 30756 3004 31756
rect 3062 30756 4062 31756
rect 4120 30756 5120 31756
rect 5178 30756 6178 31756
rect 6236 30756 7236 31756
rect 8518 30764 9518 31764
rect 9576 30764 10576 31764
rect 10634 30764 11634 31764
rect 11692 30764 12692 31764
rect 12750 30764 13750 31764
rect 15024 30772 16024 31772
rect 16082 30772 17082 31772
rect 17140 30772 18140 31772
rect 18198 30772 19198 31772
rect 19256 30772 20256 31772
rect 21514 30756 22514 31756
rect 22572 30756 23572 31756
rect 23630 30756 24630 31756
rect 24688 30756 25688 31756
rect 25746 30756 26746 31756
rect 28036 30772 29036 31772
rect 29094 30772 30094 31772
rect 30152 30772 31152 31772
rect 31210 30772 32210 31772
rect 32268 30772 33268 31772
rect 34546 30778 35546 31778
rect 35604 30778 36604 31778
rect 36662 30778 37662 31778
rect 37720 30778 38720 31778
rect 38778 30778 39778 31778
rect 41036 30778 42036 31778
rect 42094 30778 43094 31778
rect 43152 30778 44152 31778
rect 44210 30778 45210 31778
rect 45268 30778 46268 31778
rect 47624 30800 48624 31800
rect 48682 30800 49682 31800
rect 49740 30800 50740 31800
rect 50798 30800 51798 31800
rect 51856 30800 52856 31800
rect 54138 30814 55138 31814
rect 55196 30814 56196 31814
rect 56254 30814 57254 31814
rect 57312 30814 58312 31814
rect 58370 30814 59370 31814
rect 2004 29662 3004 30662
rect 3062 29662 4062 30662
rect 4120 29662 5120 30662
rect 5178 29662 6178 30662
rect 6236 29662 7236 30662
rect 2004 28568 3004 29568
rect 3062 28568 4062 29568
rect 4120 28568 5120 29568
rect 5178 28568 6178 29568
rect 6236 28568 7236 29568
rect 8518 29670 9518 30670
rect 9576 29670 10576 30670
rect 10634 29670 11634 30670
rect 11692 29670 12692 30670
rect 12750 29670 13750 30670
rect 2004 27474 3004 28474
rect 3062 27474 4062 28474
rect 4120 27474 5120 28474
rect 5178 27474 6178 28474
rect 6236 27474 7236 28474
rect 8518 28576 9518 29576
rect 9576 28576 10576 29576
rect 10634 28576 11634 29576
rect 11692 28576 12692 29576
rect 12750 28576 13750 29576
rect 15024 29678 16024 30678
rect 16082 29678 17082 30678
rect 17140 29678 18140 30678
rect 18198 29678 19198 30678
rect 19256 29678 20256 30678
rect 8518 27482 9518 28482
rect 9576 27482 10576 28482
rect 10634 27482 11634 28482
rect 11692 27482 12692 28482
rect 12750 27482 13750 28482
rect 15024 28584 16024 29584
rect 16082 28584 17082 29584
rect 17140 28584 18140 29584
rect 18198 28584 19198 29584
rect 19256 28584 20256 29584
rect 21514 29662 22514 30662
rect 22572 29662 23572 30662
rect 23630 29662 24630 30662
rect 24688 29662 25688 30662
rect 25746 29662 26746 30662
rect 15024 27490 16024 28490
rect 16082 27490 17082 28490
rect 17140 27490 18140 28490
rect 18198 27490 19198 28490
rect 19256 27490 20256 28490
rect 21514 28568 22514 29568
rect 22572 28568 23572 29568
rect 23630 28568 24630 29568
rect 24688 28568 25688 29568
rect 25746 28568 26746 29568
rect 28036 29678 29036 30678
rect 29094 29678 30094 30678
rect 30152 29678 31152 30678
rect 31210 29678 32210 30678
rect 32268 29678 33268 30678
rect 21514 27474 22514 28474
rect 22572 27474 23572 28474
rect 23630 27474 24630 28474
rect 24688 27474 25688 28474
rect 25746 27474 26746 28474
rect 28036 28584 29036 29584
rect 29094 28584 30094 29584
rect 30152 28584 31152 29584
rect 31210 28584 32210 29584
rect 32268 28584 33268 29584
rect 34546 29684 35546 30684
rect 35604 29684 36604 30684
rect 36662 29684 37662 30684
rect 37720 29684 38720 30684
rect 38778 29684 39778 30684
rect 28036 27490 29036 28490
rect 29094 27490 30094 28490
rect 30152 27490 31152 28490
rect 31210 27490 32210 28490
rect 32268 27490 33268 28490
rect 34546 28590 35546 29590
rect 35604 28590 36604 29590
rect 36662 28590 37662 29590
rect 37720 28590 38720 29590
rect 38778 28590 39778 29590
rect 41036 29684 42036 30684
rect 42094 29684 43094 30684
rect 43152 29684 44152 30684
rect 44210 29684 45210 30684
rect 45268 29684 46268 30684
rect 34546 27496 35546 28496
rect 35604 27496 36604 28496
rect 36662 27496 37662 28496
rect 37720 27496 38720 28496
rect 38778 27496 39778 28496
rect 41036 28590 42036 29590
rect 42094 28590 43094 29590
rect 43152 28590 44152 29590
rect 44210 28590 45210 29590
rect 45268 28590 46268 29590
rect 47624 29706 48624 30706
rect 48682 29706 49682 30706
rect 49740 29706 50740 30706
rect 50798 29706 51798 30706
rect 51856 29706 52856 30706
rect 41036 27496 42036 28496
rect 42094 27496 43094 28496
rect 43152 27496 44152 28496
rect 44210 27496 45210 28496
rect 45268 27496 46268 28496
rect 47624 28612 48624 29612
rect 48682 28612 49682 29612
rect 49740 28612 50740 29612
rect 50798 28612 51798 29612
rect 51856 28612 52856 29612
rect 54138 29720 55138 30720
rect 55196 29720 56196 30720
rect 56254 29720 57254 30720
rect 57312 29720 58312 30720
rect 58370 29720 59370 30720
rect 47624 27518 48624 28518
rect 48682 27518 49682 28518
rect 49740 27518 50740 28518
rect 50798 27518 51798 28518
rect 51856 27518 52856 28518
rect 54138 28626 55138 29626
rect 55196 28626 56196 29626
rect 56254 28626 57254 29626
rect 57312 28626 58312 29626
rect 58370 28626 59370 29626
rect 54138 27532 55138 28532
rect 55196 27532 56196 28532
rect 56254 27532 57254 28532
rect 57312 27532 58312 28532
rect 58370 27532 59370 28532
rect 2004 26380 3004 27380
rect 3062 26380 4062 27380
rect 4120 26380 5120 27380
rect 5178 26380 6178 27380
rect 6236 26380 7236 27380
rect 8518 26388 9518 27388
rect 9576 26388 10576 27388
rect 10634 26388 11634 27388
rect 11692 26388 12692 27388
rect 12750 26388 13750 27388
rect 15024 26396 16024 27396
rect 16082 26396 17082 27396
rect 17140 26396 18140 27396
rect 18198 26396 19198 27396
rect 19256 26396 20256 27396
rect 21514 26380 22514 27380
rect 22572 26380 23572 27380
rect 23630 26380 24630 27380
rect 24688 26380 25688 27380
rect 25746 26380 26746 27380
rect 28036 26396 29036 27396
rect 29094 26396 30094 27396
rect 30152 26396 31152 27396
rect 31210 26396 32210 27396
rect 32268 26396 33268 27396
rect 34546 26402 35546 27402
rect 35604 26402 36604 27402
rect 36662 26402 37662 27402
rect 37720 26402 38720 27402
rect 38778 26402 39778 27402
rect 41036 26402 42036 27402
rect 42094 26402 43094 27402
rect 43152 26402 44152 27402
rect 44210 26402 45210 27402
rect 45268 26402 46268 27402
rect 47624 26424 48624 27424
rect 48682 26424 49682 27424
rect 49740 26424 50740 27424
rect 50798 26424 51798 27424
rect 51856 26424 52856 27424
rect 54138 26438 55138 27438
rect 55196 26438 56196 27438
rect 56254 26438 57254 27438
rect 57312 26438 58312 27438
rect 58370 26438 59370 27438
rect 2004 24920 3004 25920
rect 3062 24920 4062 25920
rect 4120 24920 5120 25920
rect 5178 24920 6178 25920
rect 6236 24920 7236 25920
rect 8518 24928 9518 25928
rect 9576 24928 10576 25928
rect 10634 24928 11634 25928
rect 11692 24928 12692 25928
rect 12750 24928 13750 25928
rect 15024 24936 16024 25936
rect 16082 24936 17082 25936
rect 17140 24936 18140 25936
rect 18198 24936 19198 25936
rect 19256 24936 20256 25936
rect 21514 24920 22514 25920
rect 22572 24920 23572 25920
rect 23630 24920 24630 25920
rect 24688 24920 25688 25920
rect 25746 24920 26746 25920
rect 28036 24936 29036 25936
rect 29094 24936 30094 25936
rect 30152 24936 31152 25936
rect 31210 24936 32210 25936
rect 32268 24936 33268 25936
rect 34546 24942 35546 25942
rect 35604 24942 36604 25942
rect 36662 24942 37662 25942
rect 37720 24942 38720 25942
rect 38778 24942 39778 25942
rect 41036 24942 42036 25942
rect 42094 24942 43094 25942
rect 43152 24942 44152 25942
rect 44210 24942 45210 25942
rect 45268 24942 46268 25942
rect 47624 24964 48624 25964
rect 48682 24964 49682 25964
rect 49740 24964 50740 25964
rect 50798 24964 51798 25964
rect 51856 24964 52856 25964
rect 54138 24978 55138 25978
rect 55196 24978 56196 25978
rect 56254 24978 57254 25978
rect 57312 24978 58312 25978
rect 58370 24978 59370 25978
rect 2004 23826 3004 24826
rect 3062 23826 4062 24826
rect 4120 23826 5120 24826
rect 5178 23826 6178 24826
rect 6236 23826 7236 24826
rect 2004 22732 3004 23732
rect 3062 22732 4062 23732
rect 4120 22732 5120 23732
rect 5178 22732 6178 23732
rect 6236 22732 7236 23732
rect 8518 23834 9518 24834
rect 9576 23834 10576 24834
rect 10634 23834 11634 24834
rect 11692 23834 12692 24834
rect 12750 23834 13750 24834
rect 2004 21638 3004 22638
rect 3062 21638 4062 22638
rect 4120 21638 5120 22638
rect 5178 21638 6178 22638
rect 6236 21638 7236 22638
rect 8518 22740 9518 23740
rect 9576 22740 10576 23740
rect 10634 22740 11634 23740
rect 11692 22740 12692 23740
rect 12750 22740 13750 23740
rect 15024 23842 16024 24842
rect 16082 23842 17082 24842
rect 17140 23842 18140 24842
rect 18198 23842 19198 24842
rect 19256 23842 20256 24842
rect 8518 21646 9518 22646
rect 9576 21646 10576 22646
rect 10634 21646 11634 22646
rect 11692 21646 12692 22646
rect 12750 21646 13750 22646
rect 15024 22748 16024 23748
rect 16082 22748 17082 23748
rect 17140 22748 18140 23748
rect 18198 22748 19198 23748
rect 19256 22748 20256 23748
rect 21514 23826 22514 24826
rect 22572 23826 23572 24826
rect 23630 23826 24630 24826
rect 24688 23826 25688 24826
rect 25746 23826 26746 24826
rect 15024 21654 16024 22654
rect 16082 21654 17082 22654
rect 17140 21654 18140 22654
rect 18198 21654 19198 22654
rect 19256 21654 20256 22654
rect 21514 22732 22514 23732
rect 22572 22732 23572 23732
rect 23630 22732 24630 23732
rect 24688 22732 25688 23732
rect 25746 22732 26746 23732
rect 28036 23842 29036 24842
rect 29094 23842 30094 24842
rect 30152 23842 31152 24842
rect 31210 23842 32210 24842
rect 32268 23842 33268 24842
rect 21514 21638 22514 22638
rect 22572 21638 23572 22638
rect 23630 21638 24630 22638
rect 24688 21638 25688 22638
rect 25746 21638 26746 22638
rect 28036 22748 29036 23748
rect 29094 22748 30094 23748
rect 30152 22748 31152 23748
rect 31210 22748 32210 23748
rect 32268 22748 33268 23748
rect 34546 23848 35546 24848
rect 35604 23848 36604 24848
rect 36662 23848 37662 24848
rect 37720 23848 38720 24848
rect 38778 23848 39778 24848
rect 28036 21654 29036 22654
rect 29094 21654 30094 22654
rect 30152 21654 31152 22654
rect 31210 21654 32210 22654
rect 32268 21654 33268 22654
rect 34546 22754 35546 23754
rect 35604 22754 36604 23754
rect 36662 22754 37662 23754
rect 37720 22754 38720 23754
rect 38778 22754 39778 23754
rect 41036 23848 42036 24848
rect 42094 23848 43094 24848
rect 43152 23848 44152 24848
rect 44210 23848 45210 24848
rect 45268 23848 46268 24848
rect 34546 21660 35546 22660
rect 35604 21660 36604 22660
rect 36662 21660 37662 22660
rect 37720 21660 38720 22660
rect 38778 21660 39778 22660
rect 41036 22754 42036 23754
rect 42094 22754 43094 23754
rect 43152 22754 44152 23754
rect 44210 22754 45210 23754
rect 45268 22754 46268 23754
rect 47624 23870 48624 24870
rect 48682 23870 49682 24870
rect 49740 23870 50740 24870
rect 50798 23870 51798 24870
rect 51856 23870 52856 24870
rect 41036 21660 42036 22660
rect 42094 21660 43094 22660
rect 43152 21660 44152 22660
rect 44210 21660 45210 22660
rect 45268 21660 46268 22660
rect 47624 22776 48624 23776
rect 48682 22776 49682 23776
rect 49740 22776 50740 23776
rect 50798 22776 51798 23776
rect 51856 22776 52856 23776
rect 54138 23884 55138 24884
rect 55196 23884 56196 24884
rect 56254 23884 57254 24884
rect 57312 23884 58312 24884
rect 58370 23884 59370 24884
rect 47624 21682 48624 22682
rect 48682 21682 49682 22682
rect 49740 21682 50740 22682
rect 50798 21682 51798 22682
rect 51856 21682 52856 22682
rect 54138 22790 55138 23790
rect 55196 22790 56196 23790
rect 56254 22790 57254 23790
rect 57312 22790 58312 23790
rect 58370 22790 59370 23790
rect 54138 21696 55138 22696
rect 55196 21696 56196 22696
rect 56254 21696 57254 22696
rect 57312 21696 58312 22696
rect 58370 21696 59370 22696
rect 2004 20544 3004 21544
rect 3062 20544 4062 21544
rect 4120 20544 5120 21544
rect 5178 20544 6178 21544
rect 6236 20544 7236 21544
rect 8518 20552 9518 21552
rect 9576 20552 10576 21552
rect 10634 20552 11634 21552
rect 11692 20552 12692 21552
rect 12750 20552 13750 21552
rect 15024 20560 16024 21560
rect 16082 20560 17082 21560
rect 17140 20560 18140 21560
rect 18198 20560 19198 21560
rect 19256 20560 20256 21560
rect 21514 20544 22514 21544
rect 22572 20544 23572 21544
rect 23630 20544 24630 21544
rect 24688 20544 25688 21544
rect 25746 20544 26746 21544
rect 28036 20560 29036 21560
rect 29094 20560 30094 21560
rect 30152 20560 31152 21560
rect 31210 20560 32210 21560
rect 32268 20560 33268 21560
rect 34546 20566 35546 21566
rect 35604 20566 36604 21566
rect 36662 20566 37662 21566
rect 37720 20566 38720 21566
rect 38778 20566 39778 21566
rect 41036 20566 42036 21566
rect 42094 20566 43094 21566
rect 43152 20566 44152 21566
rect 44210 20566 45210 21566
rect 45268 20566 46268 21566
rect 47624 20588 48624 21588
rect 48682 20588 49682 21588
rect 49740 20588 50740 21588
rect 50798 20588 51798 21588
rect 51856 20588 52856 21588
rect 54138 20602 55138 21602
rect 55196 20602 56196 21602
rect 56254 20602 57254 21602
rect 57312 20602 58312 21602
rect 58370 20602 59370 21602
rect 2004 19056 3004 20056
rect 3062 19056 4062 20056
rect 4120 19056 5120 20056
rect 5178 19056 6178 20056
rect 6236 19056 7236 20056
rect 8518 19064 9518 20064
rect 9576 19064 10576 20064
rect 10634 19064 11634 20064
rect 11692 19064 12692 20064
rect 12750 19064 13750 20064
rect 15024 19072 16024 20072
rect 16082 19072 17082 20072
rect 17140 19072 18140 20072
rect 18198 19072 19198 20072
rect 19256 19072 20256 20072
rect 21514 19056 22514 20056
rect 22572 19056 23572 20056
rect 23630 19056 24630 20056
rect 24688 19056 25688 20056
rect 25746 19056 26746 20056
rect 28036 19072 29036 20072
rect 29094 19072 30094 20072
rect 30152 19072 31152 20072
rect 31210 19072 32210 20072
rect 32268 19072 33268 20072
rect 34546 19078 35546 20078
rect 35604 19078 36604 20078
rect 36662 19078 37662 20078
rect 37720 19078 38720 20078
rect 38778 19078 39778 20078
rect 41036 19078 42036 20078
rect 42094 19078 43094 20078
rect 43152 19078 44152 20078
rect 44210 19078 45210 20078
rect 45268 19078 46268 20078
rect 47624 19100 48624 20100
rect 48682 19100 49682 20100
rect 49740 19100 50740 20100
rect 50798 19100 51798 20100
rect 51856 19100 52856 20100
rect 54138 19114 55138 20114
rect 55196 19114 56196 20114
rect 56254 19114 57254 20114
rect 57312 19114 58312 20114
rect 58370 19114 59370 20114
rect 2004 17962 3004 18962
rect 3062 17962 4062 18962
rect 4120 17962 5120 18962
rect 5178 17962 6178 18962
rect 6236 17962 7236 18962
rect 2004 16868 3004 17868
rect 3062 16868 4062 17868
rect 4120 16868 5120 17868
rect 5178 16868 6178 17868
rect 6236 16868 7236 17868
rect 8518 17970 9518 18970
rect 9576 17970 10576 18970
rect 10634 17970 11634 18970
rect 11692 17970 12692 18970
rect 12750 17970 13750 18970
rect 2004 15774 3004 16774
rect 3062 15774 4062 16774
rect 4120 15774 5120 16774
rect 5178 15774 6178 16774
rect 6236 15774 7236 16774
rect 8518 16876 9518 17876
rect 9576 16876 10576 17876
rect 10634 16876 11634 17876
rect 11692 16876 12692 17876
rect 12750 16876 13750 17876
rect 15024 17978 16024 18978
rect 16082 17978 17082 18978
rect 17140 17978 18140 18978
rect 18198 17978 19198 18978
rect 19256 17978 20256 18978
rect 8518 15782 9518 16782
rect 9576 15782 10576 16782
rect 10634 15782 11634 16782
rect 11692 15782 12692 16782
rect 12750 15782 13750 16782
rect 15024 16884 16024 17884
rect 16082 16884 17082 17884
rect 17140 16884 18140 17884
rect 18198 16884 19198 17884
rect 19256 16884 20256 17884
rect 21514 17962 22514 18962
rect 22572 17962 23572 18962
rect 23630 17962 24630 18962
rect 24688 17962 25688 18962
rect 25746 17962 26746 18962
rect 15024 15790 16024 16790
rect 16082 15790 17082 16790
rect 17140 15790 18140 16790
rect 18198 15790 19198 16790
rect 19256 15790 20256 16790
rect 21514 16868 22514 17868
rect 22572 16868 23572 17868
rect 23630 16868 24630 17868
rect 24688 16868 25688 17868
rect 25746 16868 26746 17868
rect 28036 17978 29036 18978
rect 29094 17978 30094 18978
rect 30152 17978 31152 18978
rect 31210 17978 32210 18978
rect 32268 17978 33268 18978
rect 21514 15774 22514 16774
rect 22572 15774 23572 16774
rect 23630 15774 24630 16774
rect 24688 15774 25688 16774
rect 25746 15774 26746 16774
rect 28036 16884 29036 17884
rect 29094 16884 30094 17884
rect 30152 16884 31152 17884
rect 31210 16884 32210 17884
rect 32268 16884 33268 17884
rect 34546 17984 35546 18984
rect 35604 17984 36604 18984
rect 36662 17984 37662 18984
rect 37720 17984 38720 18984
rect 38778 17984 39778 18984
rect 28036 15790 29036 16790
rect 29094 15790 30094 16790
rect 30152 15790 31152 16790
rect 31210 15790 32210 16790
rect 32268 15790 33268 16790
rect 34546 16890 35546 17890
rect 35604 16890 36604 17890
rect 36662 16890 37662 17890
rect 37720 16890 38720 17890
rect 38778 16890 39778 17890
rect 41036 17984 42036 18984
rect 42094 17984 43094 18984
rect 43152 17984 44152 18984
rect 44210 17984 45210 18984
rect 45268 17984 46268 18984
rect 34546 15796 35546 16796
rect 35604 15796 36604 16796
rect 36662 15796 37662 16796
rect 37720 15796 38720 16796
rect 38778 15796 39778 16796
rect 41036 16890 42036 17890
rect 42094 16890 43094 17890
rect 43152 16890 44152 17890
rect 44210 16890 45210 17890
rect 45268 16890 46268 17890
rect 47624 18006 48624 19006
rect 48682 18006 49682 19006
rect 49740 18006 50740 19006
rect 50798 18006 51798 19006
rect 51856 18006 52856 19006
rect 41036 15796 42036 16796
rect 42094 15796 43094 16796
rect 43152 15796 44152 16796
rect 44210 15796 45210 16796
rect 45268 15796 46268 16796
rect 47624 16912 48624 17912
rect 48682 16912 49682 17912
rect 49740 16912 50740 17912
rect 50798 16912 51798 17912
rect 51856 16912 52856 17912
rect 54138 18020 55138 19020
rect 55196 18020 56196 19020
rect 56254 18020 57254 19020
rect 57312 18020 58312 19020
rect 58370 18020 59370 19020
rect 47624 15818 48624 16818
rect 48682 15818 49682 16818
rect 49740 15818 50740 16818
rect 50798 15818 51798 16818
rect 51856 15818 52856 16818
rect 54138 16926 55138 17926
rect 55196 16926 56196 17926
rect 56254 16926 57254 17926
rect 57312 16926 58312 17926
rect 58370 16926 59370 17926
rect 54138 15832 55138 16832
rect 55196 15832 56196 16832
rect 56254 15832 57254 16832
rect 57312 15832 58312 16832
rect 58370 15832 59370 16832
rect 2004 14680 3004 15680
rect 3062 14680 4062 15680
rect 4120 14680 5120 15680
rect 5178 14680 6178 15680
rect 6236 14680 7236 15680
rect 8518 14688 9518 15688
rect 9576 14688 10576 15688
rect 10634 14688 11634 15688
rect 11692 14688 12692 15688
rect 12750 14688 13750 15688
rect 15024 14696 16024 15696
rect 16082 14696 17082 15696
rect 17140 14696 18140 15696
rect 18198 14696 19198 15696
rect 19256 14696 20256 15696
rect 21514 14680 22514 15680
rect 22572 14680 23572 15680
rect 23630 14680 24630 15680
rect 24688 14680 25688 15680
rect 25746 14680 26746 15680
rect 28036 14696 29036 15696
rect 29094 14696 30094 15696
rect 30152 14696 31152 15696
rect 31210 14696 32210 15696
rect 32268 14696 33268 15696
rect 34546 14702 35546 15702
rect 35604 14702 36604 15702
rect 36662 14702 37662 15702
rect 37720 14702 38720 15702
rect 38778 14702 39778 15702
rect 41036 14702 42036 15702
rect 42094 14702 43094 15702
rect 43152 14702 44152 15702
rect 44210 14702 45210 15702
rect 45268 14702 46268 15702
rect 47624 14724 48624 15724
rect 48682 14724 49682 15724
rect 49740 14724 50740 15724
rect 50798 14724 51798 15724
rect 51856 14724 52856 15724
rect 54138 14738 55138 15738
rect 55196 14738 56196 15738
rect 56254 14738 57254 15738
rect 57312 14738 58312 15738
rect 58370 14738 59370 15738
rect 2014 13200 3014 14200
rect 3072 13200 4072 14200
rect 4130 13200 5130 14200
rect 5188 13200 6188 14200
rect 6246 13200 7246 14200
rect 8528 13208 9528 14208
rect 9586 13208 10586 14208
rect 10644 13208 11644 14208
rect 11702 13208 12702 14208
rect 12760 13208 13760 14208
rect 15034 13216 16034 14216
rect 16092 13216 17092 14216
rect 17150 13216 18150 14216
rect 18208 13216 19208 14216
rect 19266 13216 20266 14216
rect 21524 13200 22524 14200
rect 22582 13200 23582 14200
rect 23640 13200 24640 14200
rect 24698 13200 25698 14200
rect 25756 13200 26756 14200
rect 28046 13216 29046 14216
rect 29104 13216 30104 14216
rect 30162 13216 31162 14216
rect 31220 13216 32220 14216
rect 32278 13216 33278 14216
rect 34556 13222 35556 14222
rect 35614 13222 36614 14222
rect 36672 13222 37672 14222
rect 37730 13222 38730 14222
rect 38788 13222 39788 14222
rect 41046 13222 42046 14222
rect 42104 13222 43104 14222
rect 43162 13222 44162 14222
rect 44220 13222 45220 14222
rect 45278 13222 46278 14222
rect 47634 13244 48634 14244
rect 48692 13244 49692 14244
rect 49750 13244 50750 14244
rect 50808 13244 51808 14244
rect 51866 13244 52866 14244
rect 54148 13258 55148 14258
rect 55206 13258 56206 14258
rect 56264 13258 57264 14258
rect 57322 13258 58322 14258
rect 58380 13258 59380 14258
rect 2014 12106 3014 13106
rect 3072 12106 4072 13106
rect 4130 12106 5130 13106
rect 5188 12106 6188 13106
rect 6246 12106 7246 13106
rect 2014 11012 3014 12012
rect 3072 11012 4072 12012
rect 4130 11012 5130 12012
rect 5188 11012 6188 12012
rect 6246 11012 7246 12012
rect 8528 12114 9528 13114
rect 9586 12114 10586 13114
rect 10644 12114 11644 13114
rect 11702 12114 12702 13114
rect 12760 12114 13760 13114
rect 2014 9918 3014 10918
rect 3072 9918 4072 10918
rect 4130 9918 5130 10918
rect 5188 9918 6188 10918
rect 6246 9918 7246 10918
rect 8528 11020 9528 12020
rect 9586 11020 10586 12020
rect 10644 11020 11644 12020
rect 11702 11020 12702 12020
rect 12760 11020 13760 12020
rect 15034 12122 16034 13122
rect 16092 12122 17092 13122
rect 17150 12122 18150 13122
rect 18208 12122 19208 13122
rect 19266 12122 20266 13122
rect 8528 9926 9528 10926
rect 9586 9926 10586 10926
rect 10644 9926 11644 10926
rect 11702 9926 12702 10926
rect 12760 9926 13760 10926
rect 15034 11028 16034 12028
rect 16092 11028 17092 12028
rect 17150 11028 18150 12028
rect 18208 11028 19208 12028
rect 19266 11028 20266 12028
rect 21524 12106 22524 13106
rect 22582 12106 23582 13106
rect 23640 12106 24640 13106
rect 24698 12106 25698 13106
rect 25756 12106 26756 13106
rect 15034 9934 16034 10934
rect 16092 9934 17092 10934
rect 17150 9934 18150 10934
rect 18208 9934 19208 10934
rect 19266 9934 20266 10934
rect 21524 11012 22524 12012
rect 22582 11012 23582 12012
rect 23640 11012 24640 12012
rect 24698 11012 25698 12012
rect 25756 11012 26756 12012
rect 28046 12122 29046 13122
rect 29104 12122 30104 13122
rect 30162 12122 31162 13122
rect 31220 12122 32220 13122
rect 32278 12122 33278 13122
rect 21524 9918 22524 10918
rect 22582 9918 23582 10918
rect 23640 9918 24640 10918
rect 24698 9918 25698 10918
rect 25756 9918 26756 10918
rect 28046 11028 29046 12028
rect 29104 11028 30104 12028
rect 30162 11028 31162 12028
rect 31220 11028 32220 12028
rect 32278 11028 33278 12028
rect 34556 12128 35556 13128
rect 35614 12128 36614 13128
rect 36672 12128 37672 13128
rect 37730 12128 38730 13128
rect 38788 12128 39788 13128
rect 28046 9934 29046 10934
rect 29104 9934 30104 10934
rect 30162 9934 31162 10934
rect 31220 9934 32220 10934
rect 32278 9934 33278 10934
rect 34556 11034 35556 12034
rect 35614 11034 36614 12034
rect 36672 11034 37672 12034
rect 37730 11034 38730 12034
rect 38788 11034 39788 12034
rect 41046 12128 42046 13128
rect 42104 12128 43104 13128
rect 43162 12128 44162 13128
rect 44220 12128 45220 13128
rect 45278 12128 46278 13128
rect 34556 9940 35556 10940
rect 35614 9940 36614 10940
rect 36672 9940 37672 10940
rect 37730 9940 38730 10940
rect 38788 9940 39788 10940
rect 41046 11034 42046 12034
rect 42104 11034 43104 12034
rect 43162 11034 44162 12034
rect 44220 11034 45220 12034
rect 45278 11034 46278 12034
rect 47634 12150 48634 13150
rect 48692 12150 49692 13150
rect 49750 12150 50750 13150
rect 50808 12150 51808 13150
rect 51866 12150 52866 13150
rect 41046 9940 42046 10940
rect 42104 9940 43104 10940
rect 43162 9940 44162 10940
rect 44220 9940 45220 10940
rect 45278 9940 46278 10940
rect 47634 11056 48634 12056
rect 48692 11056 49692 12056
rect 49750 11056 50750 12056
rect 50808 11056 51808 12056
rect 51866 11056 52866 12056
rect 54148 12164 55148 13164
rect 55206 12164 56206 13164
rect 56264 12164 57264 13164
rect 57322 12164 58322 13164
rect 58380 12164 59380 13164
rect 47634 9962 48634 10962
rect 48692 9962 49692 10962
rect 49750 9962 50750 10962
rect 50808 9962 51808 10962
rect 51866 9962 52866 10962
rect 54148 11070 55148 12070
rect 55206 11070 56206 12070
rect 56264 11070 57264 12070
rect 57322 11070 58322 12070
rect 58380 11070 59380 12070
rect 54148 9976 55148 10976
rect 55206 9976 56206 10976
rect 56264 9976 57264 10976
rect 57322 9976 58322 10976
rect 58380 9976 59380 10976
rect 2014 8824 3014 9824
rect 3072 8824 4072 9824
rect 4130 8824 5130 9824
rect 5188 8824 6188 9824
rect 6246 8824 7246 9824
rect 8528 8832 9528 9832
rect 9586 8832 10586 9832
rect 10644 8832 11644 9832
rect 11702 8832 12702 9832
rect 12760 8832 13760 9832
rect 15034 8840 16034 9840
rect 16092 8840 17092 9840
rect 17150 8840 18150 9840
rect 18208 8840 19208 9840
rect 19266 8840 20266 9840
rect 21524 8824 22524 9824
rect 22582 8824 23582 9824
rect 23640 8824 24640 9824
rect 24698 8824 25698 9824
rect 25756 8824 26756 9824
rect 28046 8840 29046 9840
rect 29104 8840 30104 9840
rect 30162 8840 31162 9840
rect 31220 8840 32220 9840
rect 32278 8840 33278 9840
rect 34556 8846 35556 9846
rect 35614 8846 36614 9846
rect 36672 8846 37672 9846
rect 37730 8846 38730 9846
rect 38788 8846 39788 9846
rect 41046 8846 42046 9846
rect 42104 8846 43104 9846
rect 43162 8846 44162 9846
rect 44220 8846 45220 9846
rect 45278 8846 46278 9846
rect 47634 8868 48634 9868
rect 48692 8868 49692 9868
rect 49750 8868 50750 9868
rect 50808 8868 51808 9868
rect 51866 8868 52866 9868
rect 54148 8882 55148 9882
rect 55206 8882 56206 9882
rect 56264 8882 57264 9882
rect 57322 8882 58322 9882
rect 58380 8882 59380 9882
rect 2032 7292 3032 8292
rect 3090 7292 4090 8292
rect 4148 7292 5148 8292
rect 5206 7292 6206 8292
rect 6264 7292 7264 8292
rect 8546 7300 9546 8300
rect 9604 7300 10604 8300
rect 10662 7300 11662 8300
rect 11720 7300 12720 8300
rect 12778 7300 13778 8300
rect 15052 7308 16052 8308
rect 16110 7308 17110 8308
rect 17168 7308 18168 8308
rect 18226 7308 19226 8308
rect 19284 7308 20284 8308
rect 21542 7292 22542 8292
rect 22600 7292 23600 8292
rect 23658 7292 24658 8292
rect 24716 7292 25716 8292
rect 25774 7292 26774 8292
rect 28064 7308 29064 8308
rect 29122 7308 30122 8308
rect 30180 7308 31180 8308
rect 31238 7308 32238 8308
rect 32296 7308 33296 8308
rect 34574 7314 35574 8314
rect 35632 7314 36632 8314
rect 36690 7314 37690 8314
rect 37748 7314 38748 8314
rect 38806 7314 39806 8314
rect 41064 7314 42064 8314
rect 42122 7314 43122 8314
rect 43180 7314 44180 8314
rect 44238 7314 45238 8314
rect 45296 7314 46296 8314
rect 47652 7336 48652 8336
rect 48710 7336 49710 8336
rect 49768 7336 50768 8336
rect 50826 7336 51826 8336
rect 51884 7336 52884 8336
rect 54166 7350 55166 8350
rect 55224 7350 56224 8350
rect 56282 7350 57282 8350
rect 57340 7350 58340 8350
rect 58398 7350 59398 8350
rect 2032 6198 3032 7198
rect 3090 6198 4090 7198
rect 4148 6198 5148 7198
rect 5206 6198 6206 7198
rect 6264 6198 7264 7198
rect 2032 5104 3032 6104
rect 3090 5104 4090 6104
rect 4148 5104 5148 6104
rect 5206 5104 6206 6104
rect 6264 5104 7264 6104
rect 8546 6206 9546 7206
rect 9604 6206 10604 7206
rect 10662 6206 11662 7206
rect 11720 6206 12720 7206
rect 12778 6206 13778 7206
rect 2032 4010 3032 5010
rect 3090 4010 4090 5010
rect 4148 4010 5148 5010
rect 5206 4010 6206 5010
rect 6264 4010 7264 5010
rect 8546 5112 9546 6112
rect 9604 5112 10604 6112
rect 10662 5112 11662 6112
rect 11720 5112 12720 6112
rect 12778 5112 13778 6112
rect 15052 6214 16052 7214
rect 16110 6214 17110 7214
rect 17168 6214 18168 7214
rect 18226 6214 19226 7214
rect 19284 6214 20284 7214
rect 8546 4018 9546 5018
rect 9604 4018 10604 5018
rect 10662 4018 11662 5018
rect 11720 4018 12720 5018
rect 12778 4018 13778 5018
rect 15052 5120 16052 6120
rect 16110 5120 17110 6120
rect 17168 5120 18168 6120
rect 18226 5120 19226 6120
rect 19284 5120 20284 6120
rect 21542 6198 22542 7198
rect 22600 6198 23600 7198
rect 23658 6198 24658 7198
rect 24716 6198 25716 7198
rect 25774 6198 26774 7198
rect 15052 4026 16052 5026
rect 16110 4026 17110 5026
rect 17168 4026 18168 5026
rect 18226 4026 19226 5026
rect 19284 4026 20284 5026
rect 21542 5104 22542 6104
rect 22600 5104 23600 6104
rect 23658 5104 24658 6104
rect 24716 5104 25716 6104
rect 25774 5104 26774 6104
rect 28064 6214 29064 7214
rect 29122 6214 30122 7214
rect 30180 6214 31180 7214
rect 31238 6214 32238 7214
rect 32296 6214 33296 7214
rect 21542 4010 22542 5010
rect 22600 4010 23600 5010
rect 23658 4010 24658 5010
rect 24716 4010 25716 5010
rect 25774 4010 26774 5010
rect 28064 5120 29064 6120
rect 29122 5120 30122 6120
rect 30180 5120 31180 6120
rect 31238 5120 32238 6120
rect 32296 5120 33296 6120
rect 34574 6220 35574 7220
rect 35632 6220 36632 7220
rect 36690 6220 37690 7220
rect 37748 6220 38748 7220
rect 38806 6220 39806 7220
rect 28064 4026 29064 5026
rect 29122 4026 30122 5026
rect 30180 4026 31180 5026
rect 31238 4026 32238 5026
rect 32296 4026 33296 5026
rect 34574 5126 35574 6126
rect 35632 5126 36632 6126
rect 36690 5126 37690 6126
rect 37748 5126 38748 6126
rect 38806 5126 39806 6126
rect 41064 6220 42064 7220
rect 42122 6220 43122 7220
rect 43180 6220 44180 7220
rect 44238 6220 45238 7220
rect 45296 6220 46296 7220
rect 34574 4032 35574 5032
rect 35632 4032 36632 5032
rect 36690 4032 37690 5032
rect 37748 4032 38748 5032
rect 38806 4032 39806 5032
rect 41064 5126 42064 6126
rect 42122 5126 43122 6126
rect 43180 5126 44180 6126
rect 44238 5126 45238 6126
rect 45296 5126 46296 6126
rect 47652 6242 48652 7242
rect 48710 6242 49710 7242
rect 49768 6242 50768 7242
rect 50826 6242 51826 7242
rect 51884 6242 52884 7242
rect 41064 4032 42064 5032
rect 42122 4032 43122 5032
rect 43180 4032 44180 5032
rect 44238 4032 45238 5032
rect 45296 4032 46296 5032
rect 47652 5148 48652 6148
rect 48710 5148 49710 6148
rect 49768 5148 50768 6148
rect 50826 5148 51826 6148
rect 51884 5148 52884 6148
rect 54166 6256 55166 7256
rect 55224 6256 56224 7256
rect 56282 6256 57282 7256
rect 57340 6256 58340 7256
rect 58398 6256 59398 7256
rect 47652 4054 48652 5054
rect 48710 4054 49710 5054
rect 49768 4054 50768 5054
rect 50826 4054 51826 5054
rect 51884 4054 52884 5054
rect 54166 5162 55166 6162
rect 55224 5162 56224 6162
rect 56282 5162 57282 6162
rect 57340 5162 58340 6162
rect 58398 5162 59398 6162
rect 54166 4068 55166 5068
rect 55224 4068 56224 5068
rect 56282 4068 57282 5068
rect 57340 4068 58340 5068
rect 58398 4068 59398 5068
rect 2032 2916 3032 3916
rect 3090 2916 4090 3916
rect 4148 2916 5148 3916
rect 5206 2916 6206 3916
rect 6264 2916 7264 3916
rect 8546 2924 9546 3924
rect 9604 2924 10604 3924
rect 10662 2924 11662 3924
rect 11720 2924 12720 3924
rect 12778 2924 13778 3924
rect 15052 2932 16052 3932
rect 16110 2932 17110 3932
rect 17168 2932 18168 3932
rect 18226 2932 19226 3932
rect 19284 2932 20284 3932
rect 21542 2916 22542 3916
rect 22600 2916 23600 3916
rect 23658 2916 24658 3916
rect 24716 2916 25716 3916
rect 25774 2916 26774 3916
rect 28064 2932 29064 3932
rect 29122 2932 30122 3932
rect 30180 2932 31180 3932
rect 31238 2932 32238 3932
rect 32296 2932 33296 3932
rect 34574 2938 35574 3938
rect 35632 2938 36632 3938
rect 36690 2938 37690 3938
rect 37748 2938 38748 3938
rect 38806 2938 39806 3938
rect 41064 2938 42064 3938
rect 42122 2938 43122 3938
rect 43180 2938 44180 3938
rect 44238 2938 45238 3938
rect 45296 2938 46296 3938
rect 47652 2960 48652 3960
rect 48710 2960 49710 3960
rect 49768 2960 50768 3960
rect 50826 2960 51826 3960
rect 51884 2960 52884 3960
rect 54166 2974 55166 3974
rect 55224 2974 56224 3974
rect 56282 2974 57282 3974
rect 57340 2974 58340 3974
rect 58398 2974 59398 3974
rect 62158 24922 63158 25922
rect 63216 24922 64216 25922
rect 64274 24922 65274 25922
rect 65332 24922 66332 25922
rect 66390 24922 67390 25922
rect 68620 24920 69620 25920
rect 69678 24920 70678 25920
rect 70736 24920 71736 25920
rect 71794 24920 72794 25920
rect 72852 24920 73852 25920
rect 75314 24894 76314 25894
rect 76372 24894 77372 25894
rect 77430 24894 78430 25894
rect 78488 24894 79488 25894
rect 79546 24894 80546 25894
rect 81776 24892 82776 25892
rect 82834 24892 83834 25892
rect 83892 24892 84892 25892
rect 84950 24892 85950 25892
rect 86008 24892 87008 25892
rect 62158 23828 63158 24828
rect 63216 23828 64216 24828
rect 64274 23828 65274 24828
rect 65332 23828 66332 24828
rect 66390 23828 67390 24828
rect 88548 24886 89548 25886
rect 89606 24886 90606 25886
rect 90664 24886 91664 25886
rect 91722 24886 92722 25886
rect 92780 24886 93780 25886
rect 62158 22734 63158 23734
rect 63216 22734 64216 23734
rect 64274 22734 65274 23734
rect 65332 22734 66332 23734
rect 66390 22734 67390 23734
rect 68620 23826 69620 24826
rect 69678 23826 70678 24826
rect 70736 23826 71736 24826
rect 71794 23826 72794 24826
rect 72852 23826 73852 24826
rect 95010 24884 96010 25884
rect 96068 24884 97068 25884
rect 97126 24884 98126 25884
rect 98184 24884 99184 25884
rect 99242 24884 100242 25884
rect 62158 21640 63158 22640
rect 63216 21640 64216 22640
rect 64274 21640 65274 22640
rect 65332 21640 66332 22640
rect 66390 21640 67390 22640
rect 68620 22732 69620 23732
rect 69678 22732 70678 23732
rect 70736 22732 71736 23732
rect 71794 22732 72794 23732
rect 72852 22732 73852 23732
rect 75314 23800 76314 24800
rect 76372 23800 77372 24800
rect 77430 23800 78430 24800
rect 78488 23800 79488 24800
rect 79546 23800 80546 24800
rect 68620 21638 69620 22638
rect 69678 21638 70678 22638
rect 70736 21638 71736 22638
rect 71794 21638 72794 22638
rect 72852 21638 73852 22638
rect 75314 22706 76314 23706
rect 76372 22706 77372 23706
rect 77430 22706 78430 23706
rect 78488 22706 79488 23706
rect 79546 22706 80546 23706
rect 81776 23798 82776 24798
rect 82834 23798 83834 24798
rect 83892 23798 84892 24798
rect 84950 23798 85950 24798
rect 86008 23798 87008 24798
rect 75314 21612 76314 22612
rect 76372 21612 77372 22612
rect 77430 21612 78430 22612
rect 78488 21612 79488 22612
rect 79546 21612 80546 22612
rect 81776 22704 82776 23704
rect 82834 22704 83834 23704
rect 83892 22704 84892 23704
rect 84950 22704 85950 23704
rect 86008 22704 87008 23704
rect 88548 23792 89548 24792
rect 89606 23792 90606 24792
rect 90664 23792 91664 24792
rect 91722 23792 92722 24792
rect 92780 23792 93780 24792
rect 81776 21610 82776 22610
rect 82834 21610 83834 22610
rect 83892 21610 84892 22610
rect 84950 21610 85950 22610
rect 86008 21610 87008 22610
rect 88548 22698 89548 23698
rect 89606 22698 90606 23698
rect 90664 22698 91664 23698
rect 91722 22698 92722 23698
rect 92780 22698 93780 23698
rect 95010 23790 96010 24790
rect 96068 23790 97068 24790
rect 97126 23790 98126 24790
rect 98184 23790 99184 24790
rect 99242 23790 100242 24790
rect 62158 20546 63158 21546
rect 63216 20546 64216 21546
rect 64274 20546 65274 21546
rect 65332 20546 66332 21546
rect 66390 20546 67390 21546
rect 88548 21604 89548 22604
rect 89606 21604 90606 22604
rect 90664 21604 91664 22604
rect 91722 21604 92722 22604
rect 92780 21604 93780 22604
rect 95010 22696 96010 23696
rect 96068 22696 97068 23696
rect 97126 22696 98126 23696
rect 98184 22696 99184 23696
rect 99242 22696 100242 23696
rect 68620 20544 69620 21544
rect 69678 20544 70678 21544
rect 70736 20544 71736 21544
rect 71794 20544 72794 21544
rect 72852 20544 73852 21544
rect 95010 21602 96010 22602
rect 96068 21602 97068 22602
rect 97126 21602 98126 22602
rect 98184 21602 99184 22602
rect 99242 21602 100242 22602
rect 75314 20518 76314 21518
rect 76372 20518 77372 21518
rect 77430 20518 78430 21518
rect 78488 20518 79488 21518
rect 79546 20518 80546 21518
rect 81776 20516 82776 21516
rect 82834 20516 83834 21516
rect 83892 20516 84892 21516
rect 84950 20516 85950 21516
rect 86008 20516 87008 21516
rect 88548 20510 89548 21510
rect 89606 20510 90606 21510
rect 90664 20510 91664 21510
rect 91722 20510 92722 21510
rect 92780 20510 93780 21510
rect 95010 20508 96010 21508
rect 96068 20508 97068 21508
rect 97126 20508 98126 21508
rect 98184 20508 99184 21508
rect 99242 20508 100242 21508
rect 62164 19084 63164 20084
rect 63222 19084 64222 20084
rect 64280 19084 65280 20084
rect 65338 19084 66338 20084
rect 66396 19084 67396 20084
rect 68628 19096 69628 20096
rect 69686 19096 70686 20096
rect 70744 19096 71744 20096
rect 71802 19096 72802 20096
rect 72860 19096 73860 20096
rect 75320 19056 76320 20056
rect 76378 19056 77378 20056
rect 77436 19056 78436 20056
rect 78494 19056 79494 20056
rect 79552 19056 80552 20056
rect 81784 19068 82784 20068
rect 82842 19068 83842 20068
rect 83900 19068 84900 20068
rect 84958 19068 85958 20068
rect 86016 19068 87016 20068
rect 88554 19048 89554 20048
rect 89612 19048 90612 20048
rect 90670 19048 91670 20048
rect 91728 19048 92728 20048
rect 92786 19048 93786 20048
rect 95018 19060 96018 20060
rect 96076 19060 97076 20060
rect 97134 19060 98134 20060
rect 98192 19060 99192 20060
rect 99250 19060 100250 20060
rect 62164 17990 63164 18990
rect 63222 17990 64222 18990
rect 64280 17990 65280 18990
rect 65338 17990 66338 18990
rect 66396 17990 67396 18990
rect 62164 16896 63164 17896
rect 63222 16896 64222 17896
rect 64280 16896 65280 17896
rect 65338 16896 66338 17896
rect 66396 16896 67396 17896
rect 68628 18002 69628 19002
rect 69686 18002 70686 19002
rect 70744 18002 71744 19002
rect 71802 18002 72802 19002
rect 72860 18002 73860 19002
rect 62164 15802 63164 16802
rect 63222 15802 64222 16802
rect 64280 15802 65280 16802
rect 65338 15802 66338 16802
rect 66396 15802 67396 16802
rect 68628 16908 69628 17908
rect 69686 16908 70686 17908
rect 70744 16908 71744 17908
rect 71802 16908 72802 17908
rect 72860 16908 73860 17908
rect 75320 17962 76320 18962
rect 76378 17962 77378 18962
rect 77436 17962 78436 18962
rect 78494 17962 79494 18962
rect 79552 17962 80552 18962
rect 68628 15814 69628 16814
rect 69686 15814 70686 16814
rect 70744 15814 71744 16814
rect 71802 15814 72802 16814
rect 72860 15814 73860 16814
rect 75320 16868 76320 17868
rect 76378 16868 77378 17868
rect 77436 16868 78436 17868
rect 78494 16868 79494 17868
rect 79552 16868 80552 17868
rect 81784 17974 82784 18974
rect 82842 17974 83842 18974
rect 83900 17974 84900 18974
rect 84958 17974 85958 18974
rect 86016 17974 87016 18974
rect 75320 15774 76320 16774
rect 76378 15774 77378 16774
rect 77436 15774 78436 16774
rect 78494 15774 79494 16774
rect 79552 15774 80552 16774
rect 81784 16880 82784 17880
rect 82842 16880 83842 17880
rect 83900 16880 84900 17880
rect 84958 16880 85958 17880
rect 86016 16880 87016 17880
rect 88554 17954 89554 18954
rect 89612 17954 90612 18954
rect 90670 17954 91670 18954
rect 91728 17954 92728 18954
rect 92786 17954 93786 18954
rect 81784 15786 82784 16786
rect 82842 15786 83842 16786
rect 83900 15786 84900 16786
rect 84958 15786 85958 16786
rect 86016 15786 87016 16786
rect 88554 16860 89554 17860
rect 89612 16860 90612 17860
rect 90670 16860 91670 17860
rect 91728 16860 92728 17860
rect 92786 16860 93786 17860
rect 95018 17966 96018 18966
rect 96076 17966 97076 18966
rect 97134 17966 98134 18966
rect 98192 17966 99192 18966
rect 99250 17966 100250 18966
rect 88554 15766 89554 16766
rect 89612 15766 90612 16766
rect 90670 15766 91670 16766
rect 91728 15766 92728 16766
rect 92786 15766 93786 16766
rect 95018 16872 96018 17872
rect 96076 16872 97076 17872
rect 97134 16872 98134 17872
rect 98192 16872 99192 17872
rect 99250 16872 100250 17872
rect 95018 15778 96018 16778
rect 96076 15778 97076 16778
rect 97134 15778 98134 16778
rect 98192 15778 99192 16778
rect 99250 15778 100250 16778
rect 62164 14708 63164 15708
rect 63222 14708 64222 15708
rect 64280 14708 65280 15708
rect 65338 14708 66338 15708
rect 66396 14708 67396 15708
rect 68628 14720 69628 15720
rect 69686 14720 70686 15720
rect 70744 14720 71744 15720
rect 71802 14720 72802 15720
rect 72860 14720 73860 15720
rect 75320 14680 76320 15680
rect 76378 14680 77378 15680
rect 77436 14680 78436 15680
rect 78494 14680 79494 15680
rect 79552 14680 80552 15680
rect 81784 14692 82784 15692
rect 82842 14692 83842 15692
rect 83900 14692 84900 15692
rect 84958 14692 85958 15692
rect 86016 14692 87016 15692
rect 88554 14672 89554 15672
rect 89612 14672 90612 15672
rect 90670 14672 91670 15672
rect 91728 14672 92728 15672
rect 92786 14672 93786 15672
rect 95018 14684 96018 15684
rect 96076 14684 97076 15684
rect 97134 14684 98134 15684
rect 98192 14684 99192 15684
rect 99250 14684 100250 15684
rect 62164 13226 63164 14226
rect 63222 13226 64222 14226
rect 64280 13226 65280 14226
rect 65338 13226 66338 14226
rect 66396 13226 67396 14226
rect 68632 13224 69632 14224
rect 69690 13224 70690 14224
rect 70748 13224 71748 14224
rect 71806 13224 72806 14224
rect 72864 13224 73864 14224
rect 75320 13198 76320 14198
rect 76378 13198 77378 14198
rect 77436 13198 78436 14198
rect 78494 13198 79494 14198
rect 79552 13198 80552 14198
rect 81788 13196 82788 14196
rect 82846 13196 83846 14196
rect 83904 13196 84904 14196
rect 84962 13196 85962 14196
rect 86020 13196 87020 14196
rect 62164 12132 63164 13132
rect 63222 12132 64222 13132
rect 64280 12132 65280 13132
rect 65338 12132 66338 13132
rect 66396 12132 67396 13132
rect 88554 13190 89554 14190
rect 89612 13190 90612 14190
rect 90670 13190 91670 14190
rect 91728 13190 92728 14190
rect 92786 13190 93786 14190
rect 62164 11038 63164 12038
rect 63222 11038 64222 12038
rect 64280 11038 65280 12038
rect 65338 11038 66338 12038
rect 66396 11038 67396 12038
rect 68632 12130 69632 13130
rect 69690 12130 70690 13130
rect 70748 12130 71748 13130
rect 71806 12130 72806 13130
rect 72864 12130 73864 13130
rect 95022 13188 96022 14188
rect 96080 13188 97080 14188
rect 97138 13188 98138 14188
rect 98196 13188 99196 14188
rect 99254 13188 100254 14188
rect 62164 9944 63164 10944
rect 63222 9944 64222 10944
rect 64280 9944 65280 10944
rect 65338 9944 66338 10944
rect 66396 9944 67396 10944
rect 68632 11036 69632 12036
rect 69690 11036 70690 12036
rect 70748 11036 71748 12036
rect 71806 11036 72806 12036
rect 72864 11036 73864 12036
rect 75320 12104 76320 13104
rect 76378 12104 77378 13104
rect 77436 12104 78436 13104
rect 78494 12104 79494 13104
rect 79552 12104 80552 13104
rect 68632 9942 69632 10942
rect 69690 9942 70690 10942
rect 70748 9942 71748 10942
rect 71806 9942 72806 10942
rect 72864 9942 73864 10942
rect 75320 11010 76320 12010
rect 76378 11010 77378 12010
rect 77436 11010 78436 12010
rect 78494 11010 79494 12010
rect 79552 11010 80552 12010
rect 81788 12102 82788 13102
rect 82846 12102 83846 13102
rect 83904 12102 84904 13102
rect 84962 12102 85962 13102
rect 86020 12102 87020 13102
rect 75320 9916 76320 10916
rect 76378 9916 77378 10916
rect 77436 9916 78436 10916
rect 78494 9916 79494 10916
rect 79552 9916 80552 10916
rect 81788 11008 82788 12008
rect 82846 11008 83846 12008
rect 83904 11008 84904 12008
rect 84962 11008 85962 12008
rect 86020 11008 87020 12008
rect 88554 12096 89554 13096
rect 89612 12096 90612 13096
rect 90670 12096 91670 13096
rect 91728 12096 92728 13096
rect 92786 12096 93786 13096
rect 81788 9914 82788 10914
rect 82846 9914 83846 10914
rect 83904 9914 84904 10914
rect 84962 9914 85962 10914
rect 86020 9914 87020 10914
rect 88554 11002 89554 12002
rect 89612 11002 90612 12002
rect 90670 11002 91670 12002
rect 91728 11002 92728 12002
rect 92786 11002 93786 12002
rect 95022 12094 96022 13094
rect 96080 12094 97080 13094
rect 97138 12094 98138 13094
rect 98196 12094 99196 13094
rect 99254 12094 100254 13094
rect 62164 8850 63164 9850
rect 63222 8850 64222 9850
rect 64280 8850 65280 9850
rect 65338 8850 66338 9850
rect 66396 8850 67396 9850
rect 88554 9908 89554 10908
rect 89612 9908 90612 10908
rect 90670 9908 91670 10908
rect 91728 9908 92728 10908
rect 92786 9908 93786 10908
rect 95022 11000 96022 12000
rect 96080 11000 97080 12000
rect 97138 11000 98138 12000
rect 98196 11000 99196 12000
rect 99254 11000 100254 12000
rect 68632 8848 69632 9848
rect 69690 8848 70690 9848
rect 70748 8848 71748 9848
rect 71806 8848 72806 9848
rect 72864 8848 73864 9848
rect 95022 9906 96022 10906
rect 96080 9906 97080 10906
rect 97138 9906 98138 10906
rect 98196 9906 99196 10906
rect 99254 9906 100254 10906
rect 75320 8822 76320 9822
rect 76378 8822 77378 9822
rect 77436 8822 78436 9822
rect 78494 8822 79494 9822
rect 79552 8822 80552 9822
rect 81788 8820 82788 9820
rect 82846 8820 83846 9820
rect 83904 8820 84904 9820
rect 84962 8820 85962 9820
rect 86020 8820 87020 9820
rect 88554 8814 89554 9814
rect 89612 8814 90612 9814
rect 90670 8814 91670 9814
rect 91728 8814 92728 9814
rect 92786 8814 93786 9814
rect 62164 7368 63164 8368
rect 63222 7368 64222 8368
rect 64280 7368 65280 8368
rect 65338 7368 66338 8368
rect 66396 7368 67396 8368
rect 95022 8812 96022 9812
rect 96080 8812 97080 9812
rect 97138 8812 98138 9812
rect 98196 8812 99196 9812
rect 99254 8812 100254 9812
rect 68636 7366 69636 8366
rect 69694 7366 70694 8366
rect 70752 7366 71752 8366
rect 71810 7366 72810 8366
rect 72868 7366 73868 8366
rect 75320 7340 76320 8340
rect 76378 7340 77378 8340
rect 77436 7340 78436 8340
rect 78494 7340 79494 8340
rect 79552 7340 80552 8340
rect 81792 7338 82792 8338
rect 82850 7338 83850 8338
rect 83908 7338 84908 8338
rect 84966 7338 85966 8338
rect 86024 7338 87024 8338
rect 62164 6274 63164 7274
rect 63222 6274 64222 7274
rect 64280 6274 65280 7274
rect 65338 6274 66338 7274
rect 66396 6274 67396 7274
rect 88554 7332 89554 8332
rect 89612 7332 90612 8332
rect 90670 7332 91670 8332
rect 91728 7332 92728 8332
rect 92786 7332 93786 8332
rect 62164 5180 63164 6180
rect 63222 5180 64222 6180
rect 64280 5180 65280 6180
rect 65338 5180 66338 6180
rect 66396 5180 67396 6180
rect 68636 6272 69636 7272
rect 69694 6272 70694 7272
rect 70752 6272 71752 7272
rect 71810 6272 72810 7272
rect 72868 6272 73868 7272
rect 95026 7330 96026 8330
rect 96084 7330 97084 8330
rect 97142 7330 98142 8330
rect 98200 7330 99200 8330
rect 99258 7330 100258 8330
rect 62164 4086 63164 5086
rect 63222 4086 64222 5086
rect 64280 4086 65280 5086
rect 65338 4086 66338 5086
rect 66396 4086 67396 5086
rect 68636 5178 69636 6178
rect 69694 5178 70694 6178
rect 70752 5178 71752 6178
rect 71810 5178 72810 6178
rect 72868 5178 73868 6178
rect 75320 6246 76320 7246
rect 76378 6246 77378 7246
rect 77436 6246 78436 7246
rect 78494 6246 79494 7246
rect 79552 6246 80552 7246
rect 68636 4084 69636 5084
rect 69694 4084 70694 5084
rect 70752 4084 71752 5084
rect 71810 4084 72810 5084
rect 72868 4084 73868 5084
rect 75320 5152 76320 6152
rect 76378 5152 77378 6152
rect 77436 5152 78436 6152
rect 78494 5152 79494 6152
rect 79552 5152 80552 6152
rect 81792 6244 82792 7244
rect 82850 6244 83850 7244
rect 83908 6244 84908 7244
rect 84966 6244 85966 7244
rect 86024 6244 87024 7244
rect 75320 4058 76320 5058
rect 76378 4058 77378 5058
rect 77436 4058 78436 5058
rect 78494 4058 79494 5058
rect 79552 4058 80552 5058
rect 81792 5150 82792 6150
rect 82850 5150 83850 6150
rect 83908 5150 84908 6150
rect 84966 5150 85966 6150
rect 86024 5150 87024 6150
rect 88554 6238 89554 7238
rect 89612 6238 90612 7238
rect 90670 6238 91670 7238
rect 91728 6238 92728 7238
rect 92786 6238 93786 7238
rect 81792 4056 82792 5056
rect 82850 4056 83850 5056
rect 83908 4056 84908 5056
rect 84966 4056 85966 5056
rect 86024 4056 87024 5056
rect 88554 5144 89554 6144
rect 89612 5144 90612 6144
rect 90670 5144 91670 6144
rect 91728 5144 92728 6144
rect 92786 5144 93786 6144
rect 95026 6236 96026 7236
rect 96084 6236 97084 7236
rect 97142 6236 98142 7236
rect 98200 6236 99200 7236
rect 99258 6236 100258 7236
rect 62164 2992 63164 3992
rect 63222 2992 64222 3992
rect 64280 2992 65280 3992
rect 65338 2992 66338 3992
rect 66396 2992 67396 3992
rect 88554 4050 89554 5050
rect 89612 4050 90612 5050
rect 90670 4050 91670 5050
rect 91728 4050 92728 5050
rect 92786 4050 93786 5050
rect 95026 5142 96026 6142
rect 96084 5142 97084 6142
rect 97142 5142 98142 6142
rect 98200 5142 99200 6142
rect 99258 5142 100258 6142
rect 68636 2990 69636 3990
rect 69694 2990 70694 3990
rect 70752 2990 71752 3990
rect 71810 2990 72810 3990
rect 72868 2990 73868 3990
rect 95026 4048 96026 5048
rect 96084 4048 97084 5048
rect 97142 4048 98142 5048
rect 98200 4048 99200 5048
rect 99258 4048 100258 5048
rect 75320 2964 76320 3964
rect 76378 2964 77378 3964
rect 77436 2964 78436 3964
rect 78494 2964 79494 3964
rect 79552 2964 80552 3964
rect 81792 2962 82792 3962
rect 82850 2962 83850 3962
rect 83908 2962 84908 3962
rect 84966 2962 85966 3962
rect 86024 2962 87024 3962
rect 88554 2956 89554 3956
rect 89612 2956 90612 3956
rect 90670 2956 91670 3956
rect 91728 2956 92728 3956
rect 92786 2956 93786 3956
rect 95026 2954 96026 3954
rect 96084 2954 97084 3954
rect 97142 2954 98142 3954
rect 98200 2954 99200 3954
rect 99258 2954 100258 3954
<< mvpmos >>
rect 42196 72582 42796 73182
rect 42890 72582 43490 73182
rect 43584 72582 44184 73182
rect 44278 72582 44878 73182
rect 44972 72582 45572 73182
rect 46204 72580 46804 73180
rect 46898 72580 47498 73180
rect 47592 72580 48192 73180
rect 48286 72580 48886 73180
rect 48980 72580 49580 73180
rect 50216 72580 50816 73180
rect 50910 72580 51510 73180
rect 51604 72580 52204 73180
rect 52298 72580 52898 73180
rect 52992 72580 53592 73180
rect 54226 72580 54826 73180
rect 54920 72580 55520 73180
rect 55614 72580 56214 73180
rect 56308 72580 56908 73180
rect 57002 72580 57602 73180
rect 71384 73654 71984 74254
rect 72042 73654 72642 74254
rect 72700 73654 73300 74254
rect 73358 73654 73958 74254
rect 75248 73634 75848 74234
rect 75906 73634 76506 74234
rect 76564 73634 77164 74234
rect 77222 73634 77822 74234
rect 79098 73648 79698 74248
rect 79756 73648 80356 74248
rect 80414 73648 81014 74248
rect 81072 73648 81672 74248
rect 42196 71924 42796 72524
rect 42890 71924 43490 72524
rect 43584 71924 44184 72524
rect 44278 71924 44878 72524
rect 44972 71924 45572 72524
rect 46204 71922 46804 72522
rect 46898 71922 47498 72522
rect 47592 71922 48192 72522
rect 48286 71922 48886 72522
rect 48980 71922 49580 72522
rect 50216 71922 50816 72522
rect 50910 71922 51510 72522
rect 51604 71922 52204 72522
rect 52298 71922 52898 72522
rect 52992 71922 53592 72522
rect 54226 71922 54826 72522
rect 54920 71922 55520 72522
rect 55614 71922 56214 72522
rect 56308 71922 56908 72522
rect 57002 71922 57602 72522
rect 42196 71266 42796 71866
rect 42890 71266 43490 71866
rect 43584 71266 44184 71866
rect 44278 71266 44878 71866
rect 44972 71266 45572 71866
rect 46204 71264 46804 71864
rect 46898 71264 47498 71864
rect 47592 71264 48192 71864
rect 48286 71264 48886 71864
rect 48980 71264 49580 71864
rect 50216 71264 50816 71864
rect 50910 71264 51510 71864
rect 51604 71264 52204 71864
rect 52298 71264 52898 71864
rect 52992 71264 53592 71864
rect 54226 71264 54826 71864
rect 54920 71264 55520 71864
rect 55614 71264 56214 71864
rect 56308 71264 56908 71864
rect 57002 71264 57602 71864
rect 42196 70608 42796 71208
rect 42890 70608 43490 71208
rect 43584 70608 44184 71208
rect 44278 70608 44878 71208
rect 44972 70608 45572 71208
rect 46204 70606 46804 71206
rect 46898 70606 47498 71206
rect 47592 70606 48192 71206
rect 48286 70606 48886 71206
rect 48980 70606 49580 71206
rect 50216 70606 50816 71206
rect 50910 70606 51510 71206
rect 51604 70606 52204 71206
rect 52298 70606 52898 71206
rect 52992 70606 53592 71206
rect 54226 70606 54826 71206
rect 54920 70606 55520 71206
rect 55614 70606 56214 71206
rect 56308 70606 56908 71206
rect 57002 70606 57602 71206
rect 42196 69950 42796 70550
rect 42890 69950 43490 70550
rect 43584 69950 44184 70550
rect 44278 69950 44878 70550
rect 44972 69950 45572 70550
rect 46204 69948 46804 70548
rect 46898 69948 47498 70548
rect 47592 69948 48192 70548
rect 48286 69948 48886 70548
rect 48980 69948 49580 70548
rect 50216 69948 50816 70548
rect 50910 69948 51510 70548
rect 51604 69948 52204 70548
rect 52298 69948 52898 70548
rect 52992 69948 53592 70548
rect 54226 69948 54826 70548
rect 54920 69948 55520 70548
rect 55614 69948 56214 70548
rect 56308 69948 56908 70548
rect 57002 69948 57602 70548
rect 42188 68384 42788 68984
rect 42882 68384 43482 68984
rect 43576 68384 44176 68984
rect 44270 68384 44870 68984
rect 44964 68384 45564 68984
rect 46182 68384 46782 68984
rect 46876 68384 47476 68984
rect 47570 68384 48170 68984
rect 48264 68384 48864 68984
rect 48958 68384 49558 68984
rect 50204 68384 50804 68984
rect 50898 68384 51498 68984
rect 51592 68384 52192 68984
rect 52286 68384 52886 68984
rect 52980 68384 53580 68984
rect 54226 68384 54826 68984
rect 54920 68384 55520 68984
rect 55614 68384 56214 68984
rect 56308 68384 56908 68984
rect 57002 68384 57602 68984
rect 71356 72740 71956 73340
rect 72014 72740 72614 73340
rect 72672 72740 73272 73340
rect 73330 72740 73930 73340
rect 71356 72046 71956 72646
rect 72014 72046 72614 72646
rect 72672 72046 73272 72646
rect 73330 72046 73930 72646
rect 71356 71352 71956 71952
rect 72014 71352 72614 71952
rect 72672 71352 73272 71952
rect 73330 71352 73930 71952
rect 71356 70658 71956 71258
rect 72014 70658 72614 71258
rect 72672 70658 73272 71258
rect 73330 70658 73930 71258
rect 71356 69964 71956 70564
rect 72014 69964 72614 70564
rect 72672 69964 73272 70564
rect 73330 69964 73930 70564
rect 75220 72720 75820 73320
rect 75878 72720 76478 73320
rect 76536 72720 77136 73320
rect 77194 72720 77794 73320
rect 75220 72026 75820 72626
rect 75878 72026 76478 72626
rect 76536 72026 77136 72626
rect 77194 72026 77794 72626
rect 75220 71332 75820 71932
rect 75878 71332 76478 71932
rect 76536 71332 77136 71932
rect 77194 71332 77794 71932
rect 75220 70638 75820 71238
rect 75878 70638 76478 71238
rect 76536 70638 77136 71238
rect 77194 70638 77794 71238
rect 75220 69944 75820 70544
rect 75878 69944 76478 70544
rect 76536 69944 77136 70544
rect 77194 69944 77794 70544
rect 79070 72734 79670 73334
rect 79728 72734 80328 73334
rect 80386 72734 80986 73334
rect 81044 72734 81644 73334
rect 79070 72040 79670 72640
rect 79728 72040 80328 72640
rect 80386 72040 80986 72640
rect 81044 72040 81644 72640
rect 79070 71346 79670 71946
rect 79728 71346 80328 71946
rect 80386 71346 80986 71946
rect 81044 71346 81644 71946
rect 79070 70652 79670 71252
rect 79728 70652 80328 71252
rect 80386 70652 80986 71252
rect 81044 70652 81644 71252
rect 79070 69958 79670 70558
rect 79728 69958 80328 70558
rect 80386 69958 80986 70558
rect 81044 69958 81644 70558
rect 42188 67726 42788 68326
rect 42882 67726 43482 68326
rect 43576 67726 44176 68326
rect 44270 67726 44870 68326
rect 44964 67726 45564 68326
rect 46182 67726 46782 68326
rect 46876 67726 47476 68326
rect 47570 67726 48170 68326
rect 48264 67726 48864 68326
rect 48958 67726 49558 68326
rect 50204 67726 50804 68326
rect 50898 67726 51498 68326
rect 51592 67726 52192 68326
rect 52286 67726 52886 68326
rect 52980 67726 53580 68326
rect 54226 67726 54826 68326
rect 54920 67726 55520 68326
rect 55614 67726 56214 68326
rect 56308 67726 56908 68326
rect 57002 67726 57602 68326
rect 42188 67068 42788 67668
rect 42882 67068 43482 67668
rect 43576 67068 44176 67668
rect 44270 67068 44870 67668
rect 44964 67068 45564 67668
rect 46182 67068 46782 67668
rect 46876 67068 47476 67668
rect 47570 67068 48170 67668
rect 48264 67068 48864 67668
rect 48958 67068 49558 67668
rect 50204 67068 50804 67668
rect 50898 67068 51498 67668
rect 51592 67068 52192 67668
rect 52286 67068 52886 67668
rect 52980 67068 53580 67668
rect 54226 67068 54826 67668
rect 54920 67068 55520 67668
rect 55614 67068 56214 67668
rect 56308 67068 56908 67668
rect 57002 67068 57602 67668
rect 42188 66410 42788 67010
rect 42882 66410 43482 67010
rect 43576 66410 44176 67010
rect 44270 66410 44870 67010
rect 44964 66410 45564 67010
rect 46182 66410 46782 67010
rect 46876 66410 47476 67010
rect 47570 66410 48170 67010
rect 48264 66410 48864 67010
rect 48958 66410 49558 67010
rect 50204 66410 50804 67010
rect 50898 66410 51498 67010
rect 51592 66410 52192 67010
rect 52286 66410 52886 67010
rect 52980 66410 53580 67010
rect 54226 66410 54826 67010
rect 54920 66410 55520 67010
rect 55614 66410 56214 67010
rect 56308 66410 56908 67010
rect 57002 66410 57602 67010
rect 42188 65752 42788 66352
rect 42882 65752 43482 66352
rect 43576 65752 44176 66352
rect 44270 65752 44870 66352
rect 44964 65752 45564 66352
rect 46182 65752 46782 66352
rect 46876 65752 47476 66352
rect 47570 65752 48170 66352
rect 48264 65752 48864 66352
rect 48958 65752 49558 66352
rect 50204 65752 50804 66352
rect 50898 65752 51498 66352
rect 51592 65752 52192 66352
rect 52286 65752 52886 66352
rect 52980 65752 53580 66352
rect 54226 65752 54826 66352
rect 54920 65752 55520 66352
rect 55614 65752 56214 66352
rect 56308 65752 56908 66352
rect 57002 65752 57602 66352
rect 71352 68964 71952 69564
rect 72010 68964 72610 69564
rect 72668 68964 73268 69564
rect 73326 68964 73926 69564
rect 71352 68270 71952 68870
rect 72010 68270 72610 68870
rect 72668 68270 73268 68870
rect 73326 68270 73926 68870
rect 71352 67576 71952 68176
rect 72010 67576 72610 68176
rect 72668 67576 73268 68176
rect 73326 67576 73926 68176
rect 71352 66882 71952 67482
rect 72010 66882 72610 67482
rect 72668 66882 73268 67482
rect 73326 66882 73926 67482
rect 752 64924 1352 65524
rect 1446 64924 2046 65524
rect 2140 64924 2740 65524
rect 3420 64920 4020 65520
rect 4114 64920 4714 65520
rect 4808 64920 5408 65520
rect 6094 64926 6694 65526
rect 6788 64926 7388 65526
rect 7482 64926 8082 65526
rect 8740 64926 9340 65526
rect 9434 64926 10034 65526
rect 10128 64926 10728 65526
rect 752 64266 1352 64866
rect 1446 64266 2046 64866
rect 2140 64266 2740 64866
rect 11394 64920 11994 65520
rect 12088 64920 12688 65520
rect 12782 64920 13382 65520
rect 14048 64926 14648 65526
rect 14742 64926 15342 65526
rect 15436 64926 16036 65526
rect 16674 64930 17274 65530
rect 17368 64930 17968 65530
rect 18062 64930 18662 65530
rect 19358 64974 19958 65574
rect 20052 64974 20652 65574
rect 3420 64262 4020 64862
rect 4114 64262 4714 64862
rect 4808 64262 5408 64862
rect 6094 64268 6694 64868
rect 6788 64268 7388 64868
rect 7482 64268 8082 64868
rect 8740 64268 9340 64868
rect 9434 64268 10034 64868
rect 10128 64268 10728 64868
rect 752 63608 1352 64208
rect 1446 63608 2046 64208
rect 2140 63608 2740 64208
rect 11394 64262 11994 64862
rect 12088 64262 12688 64862
rect 12782 64262 13382 64862
rect 14048 64268 14648 64868
rect 14742 64268 15342 64868
rect 15436 64268 16036 64868
rect 16674 64272 17274 64872
rect 17368 64272 17968 64872
rect 18062 64272 18662 64872
rect 19358 64316 19958 64916
rect 20052 64316 20652 64916
rect 3420 63604 4020 64204
rect 4114 63604 4714 64204
rect 4808 63604 5408 64204
rect 6094 63610 6694 64210
rect 6788 63610 7388 64210
rect 7482 63610 8082 64210
rect 8740 63610 9340 64210
rect 9434 63610 10034 64210
rect 10128 63610 10728 64210
rect 752 62950 1352 63550
rect 1446 62950 2046 63550
rect 2140 62950 2740 63550
rect 11394 63604 11994 64204
rect 12088 63604 12688 64204
rect 12782 63604 13382 64204
rect 14048 63610 14648 64210
rect 14742 63610 15342 64210
rect 15436 63610 16036 64210
rect 16674 63614 17274 64214
rect 17368 63614 17968 64214
rect 18062 63614 18662 64214
rect 19358 63658 19958 64258
rect 20052 63658 20652 64258
rect 3420 62946 4020 63546
rect 4114 62946 4714 63546
rect 4808 62946 5408 63546
rect 6094 62952 6694 63552
rect 6788 62952 7388 63552
rect 7482 62952 8082 63552
rect 8740 62952 9340 63552
rect 9434 62952 10034 63552
rect 10128 62952 10728 63552
rect 752 62292 1352 62892
rect 1446 62292 2046 62892
rect 2140 62292 2740 62892
rect 11394 62946 11994 63546
rect 12088 62946 12688 63546
rect 12782 62946 13382 63546
rect 14048 62952 14648 63552
rect 14742 62952 15342 63552
rect 15436 62952 16036 63552
rect 16674 62956 17274 63556
rect 17368 62956 17968 63556
rect 18062 62956 18662 63556
rect 19358 63000 19958 63600
rect 20052 63000 20652 63600
rect 3420 62288 4020 62888
rect 4114 62288 4714 62888
rect 4808 62288 5408 62888
rect 6094 62294 6694 62894
rect 6788 62294 7388 62894
rect 7482 62294 8082 62894
rect 8740 62294 9340 62894
rect 9434 62294 10034 62894
rect 10128 62294 10728 62894
rect 752 61634 1352 62234
rect 1446 61634 2046 62234
rect 2140 61634 2740 62234
rect 11394 62288 11994 62888
rect 12088 62288 12688 62888
rect 12782 62288 13382 62888
rect 14048 62294 14648 62894
rect 14742 62294 15342 62894
rect 15436 62294 16036 62894
rect 16674 62298 17274 62898
rect 17368 62298 17968 62898
rect 18062 62298 18662 62898
rect 19358 62342 19958 62942
rect 20052 62342 20652 62942
rect 3420 61630 4020 62230
rect 4114 61630 4714 62230
rect 4808 61630 5408 62230
rect 6094 61636 6694 62236
rect 6788 61636 7388 62236
rect 7482 61636 8082 62236
rect 8740 61636 9340 62236
rect 9434 61636 10034 62236
rect 10128 61636 10728 62236
rect 752 60976 1352 61576
rect 1446 60976 2046 61576
rect 2140 60976 2740 61576
rect 11394 61630 11994 62230
rect 12088 61630 12688 62230
rect 12782 61630 13382 62230
rect 14048 61636 14648 62236
rect 14742 61636 15342 62236
rect 15436 61636 16036 62236
rect 16674 61640 17274 62240
rect 17368 61640 17968 62240
rect 18062 61640 18662 62240
rect 19358 61684 19958 62284
rect 20052 61684 20652 62284
rect 3420 60972 4020 61572
rect 4114 60972 4714 61572
rect 4808 60972 5408 61572
rect 6094 60978 6694 61578
rect 6788 60978 7388 61578
rect 7482 60978 8082 61578
rect 8740 60978 9340 61578
rect 9434 60978 10034 61578
rect 10128 60978 10728 61578
rect 752 60318 1352 60918
rect 1446 60318 2046 60918
rect 2140 60318 2740 60918
rect 11394 60972 11994 61572
rect 12088 60972 12688 61572
rect 12782 60972 13382 61572
rect 14048 60978 14648 61578
rect 14742 60978 15342 61578
rect 15436 60978 16036 61578
rect 16674 60982 17274 61582
rect 17368 60982 17968 61582
rect 18062 60982 18662 61582
rect 19358 61026 19958 61626
rect 20052 61026 20652 61626
rect 3420 60314 4020 60914
rect 4114 60314 4714 60914
rect 4808 60314 5408 60914
rect 6094 60320 6694 60920
rect 6788 60320 7388 60920
rect 7482 60320 8082 60920
rect 8740 60320 9340 60920
rect 9434 60320 10034 60920
rect 10128 60320 10728 60920
rect 11394 60314 11994 60914
rect 12088 60314 12688 60914
rect 12782 60314 13382 60914
rect 14048 60320 14648 60920
rect 14742 60320 15342 60920
rect 15436 60320 16036 60920
rect 16674 60324 17274 60924
rect 17368 60324 17968 60924
rect 18062 60324 18662 60924
rect 19358 60368 19958 60968
rect 20052 60368 20652 60968
rect 724 58656 1324 59256
rect 1418 58656 2018 59256
rect 2112 58656 2712 59256
rect 3392 58652 3992 59252
rect 4086 58652 4686 59252
rect 4780 58652 5380 59252
rect 6066 58658 6666 59258
rect 6760 58658 7360 59258
rect 7454 58658 8054 59258
rect 8712 58658 9312 59258
rect 9406 58658 10006 59258
rect 10100 58658 10700 59258
rect 724 57998 1324 58598
rect 1418 57998 2018 58598
rect 2112 57998 2712 58598
rect 11366 58652 11966 59252
rect 12060 58652 12660 59252
rect 12754 58652 13354 59252
rect 14020 58658 14620 59258
rect 14714 58658 15314 59258
rect 15408 58658 16008 59258
rect 16646 58662 17246 59262
rect 17340 58662 17940 59262
rect 18034 58662 18634 59262
rect 19330 58706 19930 59306
rect 20024 58706 20624 59306
rect 3392 57994 3992 58594
rect 4086 57994 4686 58594
rect 4780 57994 5380 58594
rect 6066 58000 6666 58600
rect 6760 58000 7360 58600
rect 7454 58000 8054 58600
rect 8712 58000 9312 58600
rect 9406 58000 10006 58600
rect 10100 58000 10700 58600
rect 724 57340 1324 57940
rect 1418 57340 2018 57940
rect 2112 57340 2712 57940
rect 11366 57994 11966 58594
rect 12060 57994 12660 58594
rect 12754 57994 13354 58594
rect 14020 58000 14620 58600
rect 14714 58000 15314 58600
rect 15408 58000 16008 58600
rect 16646 58004 17246 58604
rect 17340 58004 17940 58604
rect 18034 58004 18634 58604
rect 19330 58048 19930 58648
rect 20024 58048 20624 58648
rect 3392 57336 3992 57936
rect 4086 57336 4686 57936
rect 4780 57336 5380 57936
rect 6066 57342 6666 57942
rect 6760 57342 7360 57942
rect 7454 57342 8054 57942
rect 8712 57342 9312 57942
rect 9406 57342 10006 57942
rect 10100 57342 10700 57942
rect 724 56682 1324 57282
rect 1418 56682 2018 57282
rect 2112 56682 2712 57282
rect 11366 57336 11966 57936
rect 12060 57336 12660 57936
rect 12754 57336 13354 57936
rect 14020 57342 14620 57942
rect 14714 57342 15314 57942
rect 15408 57342 16008 57942
rect 16646 57346 17246 57946
rect 17340 57346 17940 57946
rect 18034 57346 18634 57946
rect 19330 57390 19930 57990
rect 20024 57390 20624 57990
rect 3392 56678 3992 57278
rect 4086 56678 4686 57278
rect 4780 56678 5380 57278
rect 6066 56684 6666 57284
rect 6760 56684 7360 57284
rect 7454 56684 8054 57284
rect 8712 56684 9312 57284
rect 9406 56684 10006 57284
rect 10100 56684 10700 57284
rect 724 56024 1324 56624
rect 1418 56024 2018 56624
rect 2112 56024 2712 56624
rect 11366 56678 11966 57278
rect 12060 56678 12660 57278
rect 12754 56678 13354 57278
rect 14020 56684 14620 57284
rect 14714 56684 15314 57284
rect 15408 56684 16008 57284
rect 16646 56688 17246 57288
rect 17340 56688 17940 57288
rect 18034 56688 18634 57288
rect 19330 56732 19930 57332
rect 20024 56732 20624 57332
rect 3392 56020 3992 56620
rect 4086 56020 4686 56620
rect 4780 56020 5380 56620
rect 6066 56026 6666 56626
rect 6760 56026 7360 56626
rect 7454 56026 8054 56626
rect 8712 56026 9312 56626
rect 9406 56026 10006 56626
rect 10100 56026 10700 56626
rect 724 55366 1324 55966
rect 1418 55366 2018 55966
rect 2112 55366 2712 55966
rect 11366 56020 11966 56620
rect 12060 56020 12660 56620
rect 12754 56020 13354 56620
rect 14020 56026 14620 56626
rect 14714 56026 15314 56626
rect 15408 56026 16008 56626
rect 16646 56030 17246 56630
rect 17340 56030 17940 56630
rect 18034 56030 18634 56630
rect 19330 56074 19930 56674
rect 20024 56074 20624 56674
rect 3392 55362 3992 55962
rect 4086 55362 4686 55962
rect 4780 55362 5380 55962
rect 6066 55368 6666 55968
rect 6760 55368 7360 55968
rect 7454 55368 8054 55968
rect 8712 55368 9312 55968
rect 9406 55368 10006 55968
rect 10100 55368 10700 55968
rect 724 54708 1324 55308
rect 1418 54708 2018 55308
rect 2112 54708 2712 55308
rect 11366 55362 11966 55962
rect 12060 55362 12660 55962
rect 12754 55362 13354 55962
rect 14020 55368 14620 55968
rect 14714 55368 15314 55968
rect 15408 55368 16008 55968
rect 16646 55372 17246 55972
rect 17340 55372 17940 55972
rect 18034 55372 18634 55972
rect 19330 55416 19930 56016
rect 20024 55416 20624 56016
rect 3392 54704 3992 55304
rect 4086 54704 4686 55304
rect 4780 54704 5380 55304
rect 6066 54710 6666 55310
rect 6760 54710 7360 55310
rect 7454 54710 8054 55310
rect 8712 54710 9312 55310
rect 9406 54710 10006 55310
rect 10100 54710 10700 55310
rect 724 54050 1324 54650
rect 1418 54050 2018 54650
rect 2112 54050 2712 54650
rect 11366 54704 11966 55304
rect 12060 54704 12660 55304
rect 12754 54704 13354 55304
rect 14020 54710 14620 55310
rect 14714 54710 15314 55310
rect 15408 54710 16008 55310
rect 16646 54714 17246 55314
rect 17340 54714 17940 55314
rect 18034 54714 18634 55314
rect 19330 54758 19930 55358
rect 20024 54758 20624 55358
rect 3392 54046 3992 54646
rect 4086 54046 4686 54646
rect 4780 54046 5380 54646
rect 6066 54052 6666 54652
rect 6760 54052 7360 54652
rect 7454 54052 8054 54652
rect 8712 54052 9312 54652
rect 9406 54052 10006 54652
rect 10100 54052 10700 54652
rect 11366 54046 11966 54646
rect 12060 54046 12660 54646
rect 12754 54046 13354 54646
rect 14020 54052 14620 54652
rect 14714 54052 15314 54652
rect 15408 54052 16008 54652
rect 16646 54056 17246 54656
rect 17340 54056 17940 54656
rect 18034 54056 18634 54656
rect 19330 54100 19930 54700
rect 20024 54100 20624 54700
rect 724 52290 1324 52890
rect 1418 52290 2018 52890
rect 2112 52290 2712 52890
rect 3392 52286 3992 52886
rect 4086 52286 4686 52886
rect 4780 52286 5380 52886
rect 6066 52292 6666 52892
rect 6760 52292 7360 52892
rect 7454 52292 8054 52892
rect 8712 52292 9312 52892
rect 9406 52292 10006 52892
rect 10100 52292 10700 52892
rect 724 51632 1324 52232
rect 1418 51632 2018 52232
rect 2112 51632 2712 52232
rect 11366 52286 11966 52886
rect 12060 52286 12660 52886
rect 12754 52286 13354 52886
rect 14020 52292 14620 52892
rect 14714 52292 15314 52892
rect 15408 52292 16008 52892
rect 16646 52296 17246 52896
rect 17340 52296 17940 52896
rect 18034 52296 18634 52896
rect 19330 52340 19930 52940
rect 20024 52340 20624 52940
rect 3392 51628 3992 52228
rect 4086 51628 4686 52228
rect 4780 51628 5380 52228
rect 6066 51634 6666 52234
rect 6760 51634 7360 52234
rect 7454 51634 8054 52234
rect 8712 51634 9312 52234
rect 9406 51634 10006 52234
rect 10100 51634 10700 52234
rect 724 50974 1324 51574
rect 1418 50974 2018 51574
rect 2112 50974 2712 51574
rect 11366 51628 11966 52228
rect 12060 51628 12660 52228
rect 12754 51628 13354 52228
rect 14020 51634 14620 52234
rect 14714 51634 15314 52234
rect 15408 51634 16008 52234
rect 16646 51638 17246 52238
rect 17340 51638 17940 52238
rect 18034 51638 18634 52238
rect 19330 51682 19930 52282
rect 20024 51682 20624 52282
rect 3392 50970 3992 51570
rect 4086 50970 4686 51570
rect 4780 50970 5380 51570
rect 6066 50976 6666 51576
rect 6760 50976 7360 51576
rect 7454 50976 8054 51576
rect 8712 50976 9312 51576
rect 9406 50976 10006 51576
rect 10100 50976 10700 51576
rect 724 50316 1324 50916
rect 1418 50316 2018 50916
rect 2112 50316 2712 50916
rect 11366 50970 11966 51570
rect 12060 50970 12660 51570
rect 12754 50970 13354 51570
rect 14020 50976 14620 51576
rect 14714 50976 15314 51576
rect 15408 50976 16008 51576
rect 16646 50980 17246 51580
rect 17340 50980 17940 51580
rect 18034 50980 18634 51580
rect 19330 51024 19930 51624
rect 20024 51024 20624 51624
rect 3392 50312 3992 50912
rect 4086 50312 4686 50912
rect 4780 50312 5380 50912
rect 6066 50318 6666 50918
rect 6760 50318 7360 50918
rect 7454 50318 8054 50918
rect 8712 50318 9312 50918
rect 9406 50318 10006 50918
rect 10100 50318 10700 50918
rect 724 49658 1324 50258
rect 1418 49658 2018 50258
rect 2112 49658 2712 50258
rect 11366 50312 11966 50912
rect 12060 50312 12660 50912
rect 12754 50312 13354 50912
rect 14020 50318 14620 50918
rect 14714 50318 15314 50918
rect 15408 50318 16008 50918
rect 16646 50322 17246 50922
rect 17340 50322 17940 50922
rect 18034 50322 18634 50922
rect 19330 50366 19930 50966
rect 20024 50366 20624 50966
rect 3392 49654 3992 50254
rect 4086 49654 4686 50254
rect 4780 49654 5380 50254
rect 6066 49660 6666 50260
rect 6760 49660 7360 50260
rect 7454 49660 8054 50260
rect 8712 49660 9312 50260
rect 9406 49660 10006 50260
rect 10100 49660 10700 50260
rect 724 49000 1324 49600
rect 1418 49000 2018 49600
rect 2112 49000 2712 49600
rect 11366 49654 11966 50254
rect 12060 49654 12660 50254
rect 12754 49654 13354 50254
rect 14020 49660 14620 50260
rect 14714 49660 15314 50260
rect 15408 49660 16008 50260
rect 16646 49664 17246 50264
rect 17340 49664 17940 50264
rect 18034 49664 18634 50264
rect 19330 49708 19930 50308
rect 20024 49708 20624 50308
rect 3392 48996 3992 49596
rect 4086 48996 4686 49596
rect 4780 48996 5380 49596
rect 6066 49002 6666 49602
rect 6760 49002 7360 49602
rect 7454 49002 8054 49602
rect 8712 49002 9312 49602
rect 9406 49002 10006 49602
rect 10100 49002 10700 49602
rect 724 48342 1324 48942
rect 1418 48342 2018 48942
rect 2112 48342 2712 48942
rect 11366 48996 11966 49596
rect 12060 48996 12660 49596
rect 12754 48996 13354 49596
rect 14020 49002 14620 49602
rect 14714 49002 15314 49602
rect 15408 49002 16008 49602
rect 16646 49006 17246 49606
rect 17340 49006 17940 49606
rect 18034 49006 18634 49606
rect 19330 49050 19930 49650
rect 20024 49050 20624 49650
rect 3392 48338 3992 48938
rect 4086 48338 4686 48938
rect 4780 48338 5380 48938
rect 6066 48344 6666 48944
rect 6760 48344 7360 48944
rect 7454 48344 8054 48944
rect 8712 48344 9312 48944
rect 9406 48344 10006 48944
rect 10100 48344 10700 48944
rect 724 47684 1324 48284
rect 1418 47684 2018 48284
rect 2112 47684 2712 48284
rect 11366 48338 11966 48938
rect 12060 48338 12660 48938
rect 12754 48338 13354 48938
rect 14020 48344 14620 48944
rect 14714 48344 15314 48944
rect 15408 48344 16008 48944
rect 16646 48348 17246 48948
rect 17340 48348 17940 48948
rect 18034 48348 18634 48948
rect 19330 48392 19930 48992
rect 20024 48392 20624 48992
rect 3392 47680 3992 48280
rect 4086 47680 4686 48280
rect 4780 47680 5380 48280
rect 6066 47686 6666 48286
rect 6760 47686 7360 48286
rect 7454 47686 8054 48286
rect 8712 47686 9312 48286
rect 9406 47686 10006 48286
rect 10100 47686 10700 48286
rect 11366 47680 11966 48280
rect 12060 47680 12660 48280
rect 12754 47680 13354 48280
rect 14020 47686 14620 48286
rect 14714 47686 15314 48286
rect 15408 47686 16008 48286
rect 16646 47690 17246 48290
rect 17340 47690 17940 48290
rect 18034 47690 18634 48290
rect 19330 47734 19930 48334
rect 20024 47734 20624 48334
rect 71352 66188 71952 66788
rect 72010 66188 72610 66788
rect 72668 66188 73268 66788
rect 73326 66188 73926 66788
rect 75216 68944 75816 69544
rect 75874 68944 76474 69544
rect 76532 68944 77132 69544
rect 77190 68944 77790 69544
rect 75216 68250 75816 68850
rect 75874 68250 76474 68850
rect 76532 68250 77132 68850
rect 77190 68250 77790 68850
rect 75216 67556 75816 68156
rect 75874 67556 76474 68156
rect 76532 67556 77132 68156
rect 77190 67556 77790 68156
rect 75216 66862 75816 67462
rect 75874 66862 76474 67462
rect 76532 66862 77132 67462
rect 77190 66862 77790 67462
rect 75216 66168 75816 66768
rect 75874 66168 76474 66768
rect 76532 66168 77132 66768
rect 77190 66168 77790 66768
rect 79066 68958 79666 69558
rect 79724 68958 80324 69558
rect 80382 68958 80982 69558
rect 81040 68958 81640 69558
rect 79066 68264 79666 68864
rect 79724 68264 80324 68864
rect 80382 68264 80982 68864
rect 81040 68264 81640 68864
rect 79066 67570 79666 68170
rect 79724 67570 80324 68170
rect 80382 67570 80982 68170
rect 81040 67570 81640 68170
rect 79066 66876 79666 67476
rect 79724 66876 80324 67476
rect 80382 66876 80982 67476
rect 81040 66876 81640 67476
rect 79066 66182 79666 66782
rect 79724 66182 80324 66782
rect 80382 66182 80982 66782
rect 81040 66182 81640 66782
rect 42176 63910 42776 64510
rect 42870 63910 43470 64510
rect 43564 63910 44164 64510
rect 44258 63910 44858 64510
rect 44952 63910 45552 64510
rect 46184 63908 46784 64508
rect 46878 63908 47478 64508
rect 47572 63908 48172 64508
rect 48266 63908 48866 64508
rect 48960 63908 49560 64508
rect 50196 63908 50796 64508
rect 50890 63908 51490 64508
rect 51584 63908 52184 64508
rect 52278 63908 52878 64508
rect 52972 63908 53572 64508
rect 54206 63908 54806 64508
rect 54900 63908 55500 64508
rect 55594 63908 56194 64508
rect 56288 63908 56888 64508
rect 56982 63908 57582 64508
rect 42176 63252 42776 63852
rect 42870 63252 43470 63852
rect 43564 63252 44164 63852
rect 44258 63252 44858 63852
rect 44952 63252 45552 63852
rect 46184 63250 46784 63850
rect 46878 63250 47478 63850
rect 47572 63250 48172 63850
rect 48266 63250 48866 63850
rect 48960 63250 49560 63850
rect 50196 63250 50796 63850
rect 50890 63250 51490 63850
rect 51584 63250 52184 63850
rect 52278 63250 52878 63850
rect 52972 63250 53572 63850
rect 54206 63250 54806 63850
rect 54900 63250 55500 63850
rect 55594 63250 56194 63850
rect 56288 63250 56888 63850
rect 56982 63250 57582 63850
rect 42176 62594 42776 63194
rect 42870 62594 43470 63194
rect 43564 62594 44164 63194
rect 44258 62594 44858 63194
rect 44952 62594 45552 63194
rect 46184 62592 46784 63192
rect 46878 62592 47478 63192
rect 47572 62592 48172 63192
rect 48266 62592 48866 63192
rect 48960 62592 49560 63192
rect 50196 62592 50796 63192
rect 50890 62592 51490 63192
rect 51584 62592 52184 63192
rect 52278 62592 52878 63192
rect 52972 62592 53572 63192
rect 54206 62592 54806 63192
rect 54900 62592 55500 63192
rect 55594 62592 56194 63192
rect 56288 62592 56888 63192
rect 56982 62592 57582 63192
rect 42176 61936 42776 62536
rect 42870 61936 43470 62536
rect 43564 61936 44164 62536
rect 44258 61936 44858 62536
rect 44952 61936 45552 62536
rect 46184 61934 46784 62534
rect 46878 61934 47478 62534
rect 47572 61934 48172 62534
rect 48266 61934 48866 62534
rect 48960 61934 49560 62534
rect 50196 61934 50796 62534
rect 50890 61934 51490 62534
rect 51584 61934 52184 62534
rect 52278 61934 52878 62534
rect 52972 61934 53572 62534
rect 54206 61934 54806 62534
rect 54900 61934 55500 62534
rect 55594 61934 56194 62534
rect 56288 61934 56888 62534
rect 56982 61934 57582 62534
rect 71352 65194 71952 65794
rect 72010 65194 72610 65794
rect 72668 65194 73268 65794
rect 73326 65194 73926 65794
rect 71352 64500 71952 65100
rect 72010 64500 72610 65100
rect 72668 64500 73268 65100
rect 73326 64500 73926 65100
rect 71352 63806 71952 64406
rect 72010 63806 72610 64406
rect 72668 63806 73268 64406
rect 73326 63806 73926 64406
rect 71352 63112 71952 63712
rect 72010 63112 72610 63712
rect 72668 63112 73268 63712
rect 73326 63112 73926 63712
rect 42176 61278 42776 61878
rect 42870 61278 43470 61878
rect 43564 61278 44164 61878
rect 44258 61278 44858 61878
rect 44952 61278 45552 61878
rect 46184 61276 46784 61876
rect 46878 61276 47478 61876
rect 47572 61276 48172 61876
rect 48266 61276 48866 61876
rect 48960 61276 49560 61876
rect 50196 61276 50796 61876
rect 50890 61276 51490 61876
rect 51584 61276 52184 61876
rect 52278 61276 52878 61876
rect 52972 61276 53572 61876
rect 54206 61276 54806 61876
rect 54900 61276 55500 61876
rect 55594 61276 56194 61876
rect 56288 61276 56888 61876
rect 56982 61276 57582 61876
rect 71352 62418 71952 63018
rect 72010 62418 72610 63018
rect 72668 62418 73268 63018
rect 73326 62418 73926 63018
rect 75216 65174 75816 65774
rect 75874 65174 76474 65774
rect 76532 65174 77132 65774
rect 77190 65174 77790 65774
rect 75216 64480 75816 65080
rect 75874 64480 76474 65080
rect 76532 64480 77132 65080
rect 77190 64480 77790 65080
rect 75216 63786 75816 64386
rect 75874 63786 76474 64386
rect 76532 63786 77132 64386
rect 77190 63786 77790 64386
rect 75216 63092 75816 63692
rect 75874 63092 76474 63692
rect 76532 63092 77132 63692
rect 77190 63092 77790 63692
rect 75216 62398 75816 62998
rect 75874 62398 76474 62998
rect 76532 62398 77132 62998
rect 77190 62398 77790 62998
rect 79066 65188 79666 65788
rect 79724 65188 80324 65788
rect 80382 65188 80982 65788
rect 81040 65188 81640 65788
rect 79066 64494 79666 65094
rect 79724 64494 80324 65094
rect 80382 64494 80982 65094
rect 81040 64494 81640 65094
rect 79066 63800 79666 64400
rect 79724 63800 80324 64400
rect 80382 63800 80982 64400
rect 81040 63800 81640 64400
rect 79066 63106 79666 63706
rect 79724 63106 80324 63706
rect 80382 63106 80982 63706
rect 81040 63106 81640 63706
rect 79066 62412 79666 63012
rect 79724 62412 80324 63012
rect 80382 62412 80982 63012
rect 81040 62412 81640 63012
rect 42168 59712 42768 60312
rect 42862 59712 43462 60312
rect 43556 59712 44156 60312
rect 44250 59712 44850 60312
rect 44944 59712 45544 60312
rect 46162 59712 46762 60312
rect 46856 59712 47456 60312
rect 47550 59712 48150 60312
rect 48244 59712 48844 60312
rect 48938 59712 49538 60312
rect 50184 59712 50784 60312
rect 50878 59712 51478 60312
rect 51572 59712 52172 60312
rect 52266 59712 52866 60312
rect 52960 59712 53560 60312
rect 54206 59712 54806 60312
rect 54900 59712 55500 60312
rect 55594 59712 56194 60312
rect 56288 59712 56888 60312
rect 56982 59712 57582 60312
rect 42168 59054 42768 59654
rect 42862 59054 43462 59654
rect 43556 59054 44156 59654
rect 44250 59054 44850 59654
rect 44944 59054 45544 59654
rect 46162 59054 46762 59654
rect 46856 59054 47456 59654
rect 47550 59054 48150 59654
rect 48244 59054 48844 59654
rect 48938 59054 49538 59654
rect 50184 59054 50784 59654
rect 50878 59054 51478 59654
rect 51572 59054 52172 59654
rect 52266 59054 52866 59654
rect 52960 59054 53560 59654
rect 54206 59054 54806 59654
rect 54900 59054 55500 59654
rect 55594 59054 56194 59654
rect 56288 59054 56888 59654
rect 56982 59054 57582 59654
rect 42168 58396 42768 58996
rect 42862 58396 43462 58996
rect 43556 58396 44156 58996
rect 44250 58396 44850 58996
rect 44944 58396 45544 58996
rect 46162 58396 46762 58996
rect 46856 58396 47456 58996
rect 47550 58396 48150 58996
rect 48244 58396 48844 58996
rect 48938 58396 49538 58996
rect 50184 58396 50784 58996
rect 50878 58396 51478 58996
rect 51572 58396 52172 58996
rect 52266 58396 52866 58996
rect 52960 58396 53560 58996
rect 54206 58396 54806 58996
rect 54900 58396 55500 58996
rect 55594 58396 56194 58996
rect 56288 58396 56888 58996
rect 56982 58396 57582 58996
rect 42168 57738 42768 58338
rect 42862 57738 43462 58338
rect 43556 57738 44156 58338
rect 44250 57738 44850 58338
rect 44944 57738 45544 58338
rect 46162 57738 46762 58338
rect 46856 57738 47456 58338
rect 47550 57738 48150 58338
rect 48244 57738 48844 58338
rect 48938 57738 49538 58338
rect 50184 57738 50784 58338
rect 50878 57738 51478 58338
rect 51572 57738 52172 58338
rect 52266 57738 52866 58338
rect 52960 57738 53560 58338
rect 54206 57738 54806 58338
rect 54900 57738 55500 58338
rect 55594 57738 56194 58338
rect 56288 57738 56888 58338
rect 56982 57738 57582 58338
rect 42168 57080 42768 57680
rect 42862 57080 43462 57680
rect 43556 57080 44156 57680
rect 44250 57080 44850 57680
rect 44944 57080 45544 57680
rect 46162 57080 46762 57680
rect 46856 57080 47456 57680
rect 47550 57080 48150 57680
rect 48244 57080 48844 57680
rect 48938 57080 49538 57680
rect 50184 57080 50784 57680
rect 50878 57080 51478 57680
rect 51572 57080 52172 57680
rect 52266 57080 52866 57680
rect 52960 57080 53560 57680
rect 54206 57080 54806 57680
rect 54900 57080 55500 57680
rect 55594 57080 56194 57680
rect 56288 57080 56888 57680
rect 56982 57080 57582 57680
rect 71352 61430 71952 62030
rect 72010 61430 72610 62030
rect 72668 61430 73268 62030
rect 73326 61430 73926 62030
rect 71352 60736 71952 61336
rect 72010 60736 72610 61336
rect 72668 60736 73268 61336
rect 73326 60736 73926 61336
rect 71352 60042 71952 60642
rect 72010 60042 72610 60642
rect 72668 60042 73268 60642
rect 73326 60042 73926 60642
rect 71352 59348 71952 59948
rect 72010 59348 72610 59948
rect 72668 59348 73268 59948
rect 73326 59348 73926 59948
rect 71352 58654 71952 59254
rect 72010 58654 72610 59254
rect 72668 58654 73268 59254
rect 73326 58654 73926 59254
rect 75216 61410 75816 62010
rect 75874 61410 76474 62010
rect 76532 61410 77132 62010
rect 77190 61410 77790 62010
rect 75216 60716 75816 61316
rect 75874 60716 76474 61316
rect 76532 60716 77132 61316
rect 77190 60716 77790 61316
rect 75216 60022 75816 60622
rect 75874 60022 76474 60622
rect 76532 60022 77132 60622
rect 77190 60022 77790 60622
rect 75216 59328 75816 59928
rect 75874 59328 76474 59928
rect 76532 59328 77132 59928
rect 77190 59328 77790 59928
rect 75216 58634 75816 59234
rect 75874 58634 76474 59234
rect 76532 58634 77132 59234
rect 77190 58634 77790 59234
rect 79066 61424 79666 62024
rect 79724 61424 80324 62024
rect 80382 61424 80982 62024
rect 81040 61424 81640 62024
rect 79066 60730 79666 61330
rect 79724 60730 80324 61330
rect 80382 60730 80982 61330
rect 81040 60730 81640 61330
rect 79066 60036 79666 60636
rect 79724 60036 80324 60636
rect 80382 60036 80982 60636
rect 81040 60036 81640 60636
rect 79066 59342 79666 59942
rect 79724 59342 80324 59942
rect 80382 59342 80982 59942
rect 81040 59342 81640 59942
rect 79066 58648 79666 59248
rect 79724 58648 80324 59248
rect 80382 58648 80982 59248
rect 81040 58648 81640 59248
rect 42120 55322 42720 55922
rect 42814 55322 43414 55922
rect 43508 55322 44108 55922
rect 44202 55322 44802 55922
rect 44896 55322 45496 55922
rect 46128 55320 46728 55920
rect 46822 55320 47422 55920
rect 47516 55320 48116 55920
rect 48210 55320 48810 55920
rect 48904 55320 49504 55920
rect 50140 55320 50740 55920
rect 50834 55320 51434 55920
rect 51528 55320 52128 55920
rect 52222 55320 52822 55920
rect 52916 55320 53516 55920
rect 54150 55320 54750 55920
rect 54844 55320 55444 55920
rect 55538 55320 56138 55920
rect 56232 55320 56832 55920
rect 56926 55320 57526 55920
rect 42120 54664 42720 55264
rect 42814 54664 43414 55264
rect 43508 54664 44108 55264
rect 44202 54664 44802 55264
rect 44896 54664 45496 55264
rect 46128 54662 46728 55262
rect 46822 54662 47422 55262
rect 47516 54662 48116 55262
rect 48210 54662 48810 55262
rect 48904 54662 49504 55262
rect 50140 54662 50740 55262
rect 50834 54662 51434 55262
rect 51528 54662 52128 55262
rect 52222 54662 52822 55262
rect 52916 54662 53516 55262
rect 54150 54662 54750 55262
rect 54844 54662 55444 55262
rect 55538 54662 56138 55262
rect 56232 54662 56832 55262
rect 56926 54662 57526 55262
rect 42120 54006 42720 54606
rect 42814 54006 43414 54606
rect 43508 54006 44108 54606
rect 44202 54006 44802 54606
rect 44896 54006 45496 54606
rect 46128 54004 46728 54604
rect 46822 54004 47422 54604
rect 47516 54004 48116 54604
rect 48210 54004 48810 54604
rect 48904 54004 49504 54604
rect 50140 54004 50740 54604
rect 50834 54004 51434 54604
rect 51528 54004 52128 54604
rect 52222 54004 52822 54604
rect 52916 54004 53516 54604
rect 54150 54004 54750 54604
rect 54844 54004 55444 54604
rect 55538 54004 56138 54604
rect 56232 54004 56832 54604
rect 56926 54004 57526 54604
rect 42120 53348 42720 53948
rect 42814 53348 43414 53948
rect 43508 53348 44108 53948
rect 44202 53348 44802 53948
rect 44896 53348 45496 53948
rect 46128 53346 46728 53946
rect 46822 53346 47422 53946
rect 47516 53346 48116 53946
rect 48210 53346 48810 53946
rect 48904 53346 49504 53946
rect 50140 53346 50740 53946
rect 50834 53346 51434 53946
rect 51528 53346 52128 53946
rect 52222 53346 52822 53946
rect 52916 53346 53516 53946
rect 54150 53346 54750 53946
rect 54844 53346 55444 53946
rect 55538 53346 56138 53946
rect 56232 53346 56832 53946
rect 56926 53346 57526 53946
rect 71352 57654 71952 58254
rect 72010 57654 72610 58254
rect 72668 57654 73268 58254
rect 73326 57654 73926 58254
rect 71352 56960 71952 57560
rect 72010 56960 72610 57560
rect 72668 56960 73268 57560
rect 73326 56960 73926 57560
rect 71352 56266 71952 56866
rect 72010 56266 72610 56866
rect 72668 56266 73268 56866
rect 73326 56266 73926 56866
rect 71352 55572 71952 56172
rect 72010 55572 72610 56172
rect 72668 55572 73268 56172
rect 73326 55572 73926 56172
rect 71352 54878 71952 55478
rect 72010 54878 72610 55478
rect 72668 54878 73268 55478
rect 73326 54878 73926 55478
rect 75216 57634 75816 58234
rect 75874 57634 76474 58234
rect 76532 57634 77132 58234
rect 77190 57634 77790 58234
rect 75216 56940 75816 57540
rect 75874 56940 76474 57540
rect 76532 56940 77132 57540
rect 77190 56940 77790 57540
rect 75216 56246 75816 56846
rect 75874 56246 76474 56846
rect 76532 56246 77132 56846
rect 77190 56246 77790 56846
rect 75216 55552 75816 56152
rect 75874 55552 76474 56152
rect 76532 55552 77132 56152
rect 77190 55552 77790 56152
rect 75216 54858 75816 55458
rect 75874 54858 76474 55458
rect 76532 54858 77132 55458
rect 77190 54858 77790 55458
rect 79066 57648 79666 58248
rect 79724 57648 80324 58248
rect 80382 57648 80982 58248
rect 81040 57648 81640 58248
rect 79066 56954 79666 57554
rect 79724 56954 80324 57554
rect 80382 56954 80982 57554
rect 81040 56954 81640 57554
rect 79066 56260 79666 56860
rect 79724 56260 80324 56860
rect 80382 56260 80982 56860
rect 81040 56260 81640 56860
rect 79066 55566 79666 56166
rect 79724 55566 80324 56166
rect 80382 55566 80982 56166
rect 81040 55566 81640 56166
rect 79066 54872 79666 55472
rect 79724 54872 80324 55472
rect 80382 54872 80982 55472
rect 81040 54872 81640 55472
rect 42120 52690 42720 53290
rect 42814 52690 43414 53290
rect 43508 52690 44108 53290
rect 44202 52690 44802 53290
rect 44896 52690 45496 53290
rect 46128 52688 46728 53288
rect 46822 52688 47422 53288
rect 47516 52688 48116 53288
rect 48210 52688 48810 53288
rect 48904 52688 49504 53288
rect 50140 52688 50740 53288
rect 50834 52688 51434 53288
rect 51528 52688 52128 53288
rect 52222 52688 52822 53288
rect 52916 52688 53516 53288
rect 54150 52688 54750 53288
rect 54844 52688 55444 53288
rect 55538 52688 56138 53288
rect 56232 52688 56832 53288
rect 56926 52688 57526 53288
rect 42112 51124 42712 51724
rect 42806 51124 43406 51724
rect 43500 51124 44100 51724
rect 44194 51124 44794 51724
rect 44888 51124 45488 51724
rect 46106 51124 46706 51724
rect 46800 51124 47400 51724
rect 47494 51124 48094 51724
rect 48188 51124 48788 51724
rect 48882 51124 49482 51724
rect 50128 51124 50728 51724
rect 50822 51124 51422 51724
rect 51516 51124 52116 51724
rect 52210 51124 52810 51724
rect 52904 51124 53504 51724
rect 54150 51124 54750 51724
rect 54844 51124 55444 51724
rect 55538 51124 56138 51724
rect 56232 51124 56832 51724
rect 56926 51124 57526 51724
rect 71356 53882 71956 54482
rect 72014 53882 72614 54482
rect 72672 53882 73272 54482
rect 73330 53882 73930 54482
rect 71356 53188 71956 53788
rect 72014 53188 72614 53788
rect 72672 53188 73272 53788
rect 73330 53188 73930 53788
rect 71356 52494 71956 53094
rect 72014 52494 72614 53094
rect 72672 52494 73272 53094
rect 73330 52494 73930 53094
rect 71356 51800 71956 52400
rect 72014 51800 72614 52400
rect 72672 51800 73272 52400
rect 73330 51800 73930 52400
rect 42112 50466 42712 51066
rect 42806 50466 43406 51066
rect 43500 50466 44100 51066
rect 44194 50466 44794 51066
rect 44888 50466 45488 51066
rect 46106 50466 46706 51066
rect 46800 50466 47400 51066
rect 47494 50466 48094 51066
rect 48188 50466 48788 51066
rect 48882 50466 49482 51066
rect 50128 50466 50728 51066
rect 50822 50466 51422 51066
rect 51516 50466 52116 51066
rect 52210 50466 52810 51066
rect 52904 50466 53504 51066
rect 54150 50466 54750 51066
rect 54844 50466 55444 51066
rect 55538 50466 56138 51066
rect 56232 50466 56832 51066
rect 56926 50466 57526 51066
rect 71356 51106 71956 51706
rect 72014 51106 72614 51706
rect 72672 51106 73272 51706
rect 73330 51106 73930 51706
rect 75220 53862 75820 54462
rect 75878 53862 76478 54462
rect 76536 53862 77136 54462
rect 77194 53862 77794 54462
rect 75220 53168 75820 53768
rect 75878 53168 76478 53768
rect 76536 53168 77136 53768
rect 77194 53168 77794 53768
rect 75220 52474 75820 53074
rect 75878 52474 76478 53074
rect 76536 52474 77136 53074
rect 77194 52474 77794 53074
rect 75220 51780 75820 52380
rect 75878 51780 76478 52380
rect 76536 51780 77136 52380
rect 77194 51780 77794 52380
rect 75220 51086 75820 51686
rect 75878 51086 76478 51686
rect 76536 51086 77136 51686
rect 77194 51086 77794 51686
rect 79070 53876 79670 54476
rect 79728 53876 80328 54476
rect 80386 53876 80986 54476
rect 81044 53876 81644 54476
rect 79070 53182 79670 53782
rect 79728 53182 80328 53782
rect 80386 53182 80986 53782
rect 81044 53182 81644 53782
rect 79070 52488 79670 53088
rect 79728 52488 80328 53088
rect 80386 52488 80986 53088
rect 81044 52488 81644 53088
rect 79070 51794 79670 52394
rect 79728 51794 80328 52394
rect 80386 51794 80986 52394
rect 81044 51794 81644 52394
rect 79070 51100 79670 51700
rect 79728 51100 80328 51700
rect 80386 51100 80986 51700
rect 81044 51100 81644 51700
rect 83355 53805 83455 53955
rect 83511 53805 83611 53955
rect 83781 53900 83881 53984
rect 83937 53900 84037 53984
rect 84093 53900 84193 53984
rect 84249 53900 84349 53984
rect 84391 53900 84491 53984
rect 84563 53900 84663 53984
rect 84891 53811 84991 54011
rect 85047 53811 85147 54011
rect 85226 53811 85326 53895
rect 85368 53811 85468 53895
rect 85545 53811 85645 53895
rect 85701 53811 85801 53895
rect 85986 53711 86086 53861
rect 86161 53711 86261 54011
rect 42112 49808 42712 50408
rect 42806 49808 43406 50408
rect 43500 49808 44100 50408
rect 44194 49808 44794 50408
rect 44888 49808 45488 50408
rect 46106 49808 46706 50408
rect 46800 49808 47400 50408
rect 47494 49808 48094 50408
rect 48188 49808 48788 50408
rect 48882 49808 49482 50408
rect 50128 49808 50728 50408
rect 50822 49808 51422 50408
rect 51516 49808 52116 50408
rect 52210 49808 52810 50408
rect 52904 49808 53504 50408
rect 54150 49808 54750 50408
rect 54844 49808 55444 50408
rect 55538 49808 56138 50408
rect 56232 49808 56832 50408
rect 56926 49808 57526 50408
rect 42112 49150 42712 49750
rect 42806 49150 43406 49750
rect 43500 49150 44100 49750
rect 44194 49150 44794 49750
rect 44888 49150 45488 49750
rect 46106 49150 46706 49750
rect 46800 49150 47400 49750
rect 47494 49150 48094 49750
rect 48188 49150 48788 49750
rect 48882 49150 49482 49750
rect 50128 49150 50728 49750
rect 50822 49150 51422 49750
rect 51516 49150 52116 49750
rect 52210 49150 52810 49750
rect 52904 49150 53504 49750
rect 54150 49150 54750 49750
rect 54844 49150 55444 49750
rect 55538 49150 56138 49750
rect 56232 49150 56832 49750
rect 56926 49150 57526 49750
rect 42112 48492 42712 49092
rect 42806 48492 43406 49092
rect 43500 48492 44100 49092
rect 44194 48492 44794 49092
rect 44888 48492 45488 49092
rect 46106 48492 46706 49092
rect 46800 48492 47400 49092
rect 47494 48492 48094 49092
rect 48188 48492 48788 49092
rect 48882 48492 49482 49092
rect 50128 48492 50728 49092
rect 50822 48492 51422 49092
rect 51516 48492 52116 49092
rect 52210 48492 52810 49092
rect 52904 48492 53504 49092
rect 54150 48492 54750 49092
rect 54844 48492 55444 49092
rect 55538 48492 56138 49092
rect 56232 48492 56832 49092
rect 56926 48492 57526 49092
<< mvndiff >>
rect 23420 57480 24020 57492
rect 23420 57446 23634 57480
rect 23806 57446 24020 57480
rect 23420 57434 24020 57446
rect 24114 57480 24714 57492
rect 24114 57446 24328 57480
rect 24500 57446 24714 57480
rect 24114 57434 24714 57446
rect 24808 57480 25408 57492
rect 24808 57446 25022 57480
rect 25194 57446 25408 57480
rect 24808 57434 25408 57446
rect 25502 57480 26102 57492
rect 25502 57446 25716 57480
rect 25888 57446 26102 57480
rect 25502 57434 26102 57446
rect 26196 57480 26796 57492
rect 26196 57446 26410 57480
rect 26582 57446 26796 57480
rect 26196 57434 26796 57446
rect 26890 57480 27490 57492
rect 26890 57446 27104 57480
rect 27276 57446 27490 57480
rect 26890 57434 27490 57446
rect 27584 57480 28184 57492
rect 27584 57446 27798 57480
rect 27970 57446 28184 57480
rect 27584 57434 28184 57446
rect 28278 57480 28878 57492
rect 28278 57446 28492 57480
rect 28664 57446 28878 57480
rect 28278 57434 28878 57446
rect 28972 57480 29572 57492
rect 28972 57446 29186 57480
rect 29358 57446 29572 57480
rect 28972 57434 29572 57446
rect 29666 57480 30266 57492
rect 29666 57446 29880 57480
rect 30052 57446 30266 57480
rect 29666 57434 30266 57446
rect 23420 56822 24020 56834
rect 23420 56788 23634 56822
rect 23806 56788 24020 56822
rect 23420 56776 24020 56788
rect 24114 56822 24714 56834
rect 24114 56788 24328 56822
rect 24500 56788 24714 56822
rect 24114 56776 24714 56788
rect 24808 56822 25408 56834
rect 24808 56788 25022 56822
rect 25194 56788 25408 56822
rect 24808 56776 25408 56788
rect 25502 56822 26102 56834
rect 25502 56788 25716 56822
rect 25888 56788 26102 56822
rect 25502 56776 26102 56788
rect 26196 56822 26796 56834
rect 26196 56788 26410 56822
rect 26582 56788 26796 56822
rect 26196 56776 26796 56788
rect 26890 56822 27490 56834
rect 26890 56788 27104 56822
rect 27276 56788 27490 56822
rect 26890 56776 27490 56788
rect 27584 56822 28184 56834
rect 27584 56788 27798 56822
rect 27970 56788 28184 56822
rect 27584 56776 28184 56788
rect 28278 56822 28878 56834
rect 28278 56788 28492 56822
rect 28664 56788 28878 56822
rect 28278 56776 28878 56788
rect 28972 56822 29572 56834
rect 28972 56788 29186 56822
rect 29358 56788 29572 56822
rect 28972 56776 29572 56788
rect 29666 56822 30266 56834
rect 29666 56788 29880 56822
rect 30052 56788 30266 56822
rect 29666 56776 30266 56788
rect 23420 56164 24020 56176
rect 23420 56130 23634 56164
rect 23806 56130 24020 56164
rect 23420 56118 24020 56130
rect 24114 56164 24714 56176
rect 24114 56130 24328 56164
rect 24500 56130 24714 56164
rect 24114 56118 24714 56130
rect 24808 56164 25408 56176
rect 24808 56130 25022 56164
rect 25194 56130 25408 56164
rect 24808 56118 25408 56130
rect 25502 56164 26102 56176
rect 25502 56130 25716 56164
rect 25888 56130 26102 56164
rect 25502 56118 26102 56130
rect 26196 56164 26796 56176
rect 26196 56130 26410 56164
rect 26582 56130 26796 56164
rect 26196 56118 26796 56130
rect 26890 56164 27490 56176
rect 26890 56130 27104 56164
rect 27276 56130 27490 56164
rect 26890 56118 27490 56130
rect 27584 56164 28184 56176
rect 27584 56130 27798 56164
rect 27970 56130 28184 56164
rect 27584 56118 28184 56130
rect 28278 56164 28878 56176
rect 28278 56130 28492 56164
rect 28664 56130 28878 56164
rect 28278 56118 28878 56130
rect 28972 56164 29572 56176
rect 28972 56130 29186 56164
rect 29358 56130 29572 56164
rect 28972 56118 29572 56130
rect 29666 56164 30266 56176
rect 29666 56130 29880 56164
rect 30052 56130 30266 56164
rect 29666 56118 30266 56130
rect 23426 55590 24026 55602
rect 23426 55556 23640 55590
rect 23812 55556 24026 55590
rect 23426 55544 24026 55556
rect 24120 55590 24720 55602
rect 24120 55556 24334 55590
rect 24506 55556 24720 55590
rect 24120 55544 24720 55556
rect 24814 55590 25414 55602
rect 24814 55556 25028 55590
rect 25200 55556 25414 55590
rect 24814 55544 25414 55556
rect 25508 55590 26108 55602
rect 25508 55556 25722 55590
rect 25894 55556 26108 55590
rect 25508 55544 26108 55556
rect 26202 55590 26802 55602
rect 26202 55556 26416 55590
rect 26588 55556 26802 55590
rect 26202 55544 26802 55556
rect 26896 55590 27496 55602
rect 26896 55556 27110 55590
rect 27282 55556 27496 55590
rect 26896 55544 27496 55556
rect 27590 55590 28190 55602
rect 27590 55556 27804 55590
rect 27976 55556 28190 55590
rect 27590 55544 28190 55556
rect 28284 55590 28884 55602
rect 28284 55556 28498 55590
rect 28670 55556 28884 55590
rect 28284 55544 28884 55556
rect 28978 55590 29578 55602
rect 28978 55556 29192 55590
rect 29364 55556 29578 55590
rect 28978 55544 29578 55556
rect 29672 55590 30272 55602
rect 29672 55556 29886 55590
rect 30058 55556 30272 55590
rect 29672 55544 30272 55556
rect 23426 54932 24026 54944
rect 23426 54898 23640 54932
rect 23812 54898 24026 54932
rect 23426 54886 24026 54898
rect 24120 54932 24720 54944
rect 24120 54898 24334 54932
rect 24506 54898 24720 54932
rect 24120 54886 24720 54898
rect 24814 54932 25414 54944
rect 24814 54898 25028 54932
rect 25200 54898 25414 54932
rect 24814 54886 25414 54898
rect 25508 54932 26108 54944
rect 25508 54898 25722 54932
rect 25894 54898 26108 54932
rect 25508 54886 26108 54898
rect 26202 54932 26802 54944
rect 26202 54898 26416 54932
rect 26588 54898 26802 54932
rect 26202 54886 26802 54898
rect 26896 54932 27496 54944
rect 26896 54898 27110 54932
rect 27282 54898 27496 54932
rect 26896 54886 27496 54898
rect 27590 54932 28190 54944
rect 27590 54898 27804 54932
rect 27976 54898 28190 54932
rect 27590 54886 28190 54898
rect 28284 54932 28884 54944
rect 28284 54898 28498 54932
rect 28670 54898 28884 54932
rect 28284 54886 28884 54898
rect 28978 54932 29578 54944
rect 28978 54898 29192 54932
rect 29364 54898 29578 54932
rect 28978 54886 29578 54898
rect 29672 54932 30272 54944
rect 29672 54898 29886 54932
rect 30058 54898 30272 54932
rect 29672 54886 30272 54898
rect 23426 54274 24026 54286
rect 23426 54240 23640 54274
rect 23812 54240 24026 54274
rect 23426 54228 24026 54240
rect 24120 54274 24720 54286
rect 24120 54240 24334 54274
rect 24506 54240 24720 54274
rect 24120 54228 24720 54240
rect 24814 54274 25414 54286
rect 24814 54240 25028 54274
rect 25200 54240 25414 54274
rect 24814 54228 25414 54240
rect 25508 54274 26108 54286
rect 25508 54240 25722 54274
rect 25894 54240 26108 54274
rect 25508 54228 26108 54240
rect 26202 54274 26802 54286
rect 26202 54240 26416 54274
rect 26588 54240 26802 54274
rect 26202 54228 26802 54240
rect 26896 54274 27496 54286
rect 26896 54240 27110 54274
rect 27282 54240 27496 54274
rect 26896 54228 27496 54240
rect 27590 54274 28190 54286
rect 27590 54240 27804 54274
rect 27976 54240 28190 54274
rect 27590 54228 28190 54240
rect 28284 54274 28884 54286
rect 28284 54240 28498 54274
rect 28670 54240 28884 54274
rect 28284 54228 28884 54240
rect 28978 54274 29578 54286
rect 28978 54240 29192 54274
rect 29364 54240 29578 54274
rect 28978 54228 29578 54240
rect 29672 54274 30272 54286
rect 29672 54240 29886 54274
rect 30058 54240 30272 54274
rect 29672 54228 30272 54240
rect 23442 53648 24042 53660
rect 23442 53614 23656 53648
rect 23828 53614 24042 53648
rect 23442 53602 24042 53614
rect 24136 53648 24736 53660
rect 24136 53614 24350 53648
rect 24522 53614 24736 53648
rect 24136 53602 24736 53614
rect 24830 53648 25430 53660
rect 24830 53614 25044 53648
rect 25216 53614 25430 53648
rect 24830 53602 25430 53614
rect 25524 53648 26124 53660
rect 25524 53614 25738 53648
rect 25910 53614 26124 53648
rect 25524 53602 26124 53614
rect 26218 53648 26818 53660
rect 26218 53614 26432 53648
rect 26604 53614 26818 53648
rect 26218 53602 26818 53614
rect 26912 53648 27512 53660
rect 26912 53614 27126 53648
rect 27298 53614 27512 53648
rect 26912 53602 27512 53614
rect 27606 53648 28206 53660
rect 27606 53614 27820 53648
rect 27992 53614 28206 53648
rect 27606 53602 28206 53614
rect 28300 53648 28900 53660
rect 28300 53614 28514 53648
rect 28686 53614 28900 53648
rect 28300 53602 28900 53614
rect 28994 53648 29594 53660
rect 28994 53614 29208 53648
rect 29380 53614 29594 53648
rect 28994 53602 29594 53614
rect 29688 53648 30288 53660
rect 29688 53614 29902 53648
rect 30074 53614 30288 53648
rect 29688 53602 30288 53614
rect 23442 52990 24042 53002
rect 23442 52956 23656 52990
rect 23828 52956 24042 52990
rect 23442 52944 24042 52956
rect 24136 52990 24736 53002
rect 24136 52956 24350 52990
rect 24522 52956 24736 52990
rect 24136 52944 24736 52956
rect 24830 52990 25430 53002
rect 24830 52956 25044 52990
rect 25216 52956 25430 52990
rect 24830 52944 25430 52956
rect 25524 52990 26124 53002
rect 25524 52956 25738 52990
rect 25910 52956 26124 52990
rect 25524 52944 26124 52956
rect 26218 52990 26818 53002
rect 26218 52956 26432 52990
rect 26604 52956 26818 52990
rect 26218 52944 26818 52956
rect 26912 52990 27512 53002
rect 26912 52956 27126 52990
rect 27298 52956 27512 52990
rect 26912 52944 27512 52956
rect 27606 52990 28206 53002
rect 27606 52956 27820 52990
rect 27992 52956 28206 52990
rect 27606 52944 28206 52956
rect 28300 52990 28900 53002
rect 28300 52956 28514 52990
rect 28686 52956 28900 52990
rect 28300 52944 28900 52956
rect 28994 52990 29594 53002
rect 28994 52956 29208 52990
rect 29380 52956 29594 52990
rect 28994 52944 29594 52956
rect 29688 52990 30288 53002
rect 29688 52956 29902 52990
rect 30074 52956 30288 52990
rect 29688 52944 30288 52956
rect 23442 52332 24042 52344
rect 23442 52298 23656 52332
rect 23828 52298 24042 52332
rect 23442 52286 24042 52298
rect 24136 52332 24736 52344
rect 24136 52298 24350 52332
rect 24522 52298 24736 52332
rect 24136 52286 24736 52298
rect 24830 52332 25430 52344
rect 24830 52298 25044 52332
rect 25216 52298 25430 52332
rect 24830 52286 25430 52298
rect 25524 52332 26124 52344
rect 25524 52298 25738 52332
rect 25910 52298 26124 52332
rect 25524 52286 26124 52298
rect 26218 52332 26818 52344
rect 26218 52298 26432 52332
rect 26604 52298 26818 52332
rect 26218 52286 26818 52298
rect 26912 52332 27512 52344
rect 26912 52298 27126 52332
rect 27298 52298 27512 52332
rect 26912 52286 27512 52298
rect 27606 52332 28206 52344
rect 27606 52298 27820 52332
rect 27992 52298 28206 52332
rect 27606 52286 28206 52298
rect 28300 52332 28900 52344
rect 28300 52298 28514 52332
rect 28686 52298 28900 52332
rect 28300 52286 28900 52298
rect 28994 52332 29594 52344
rect 28994 52298 29208 52332
rect 29380 52298 29594 52332
rect 28994 52286 29594 52298
rect 29688 52332 30288 52344
rect 29688 52298 29902 52332
rect 30074 52298 30288 52332
rect 29688 52286 30288 52298
rect 83752 53500 83809 53525
rect 83752 53466 83764 53500
rect 83798 53466 83809 53500
rect 83302 53434 83359 53459
rect 83302 53400 83314 53434
rect 83348 53400 83359 53434
rect 83302 53375 83359 53400
rect 83459 53434 83515 53459
rect 83459 53400 83470 53434
rect 83504 53400 83515 53434
rect 83459 53375 83515 53400
rect 83615 53434 83672 53459
rect 83752 53441 83809 53466
rect 83909 53441 83951 53525
rect 84051 53500 84107 53525
rect 84051 53466 84062 53500
rect 84096 53466 84107 53500
rect 84051 53441 84107 53466
rect 84207 53500 84263 53525
rect 84207 53466 84218 53500
rect 84252 53466 84263 53500
rect 84207 53441 84263 53466
rect 84363 53441 84405 53525
rect 84505 53441 84552 53525
rect 84652 53441 84905 53525
rect 83615 53400 83626 53434
rect 83660 53400 83672 53434
rect 84832 53437 84905 53441
rect 83615 53375 83672 53400
rect 84832 53403 84844 53437
rect 84878 53403 84905 53437
rect 84832 53375 84905 53403
rect 85005 53517 85061 53525
rect 85005 53483 85016 53517
rect 85050 53483 85061 53517
rect 85005 53425 85061 53483
rect 85005 53391 85016 53425
rect 85050 53391 85061 53425
rect 85005 53375 85061 53391
rect 85161 53517 85220 53525
rect 85161 53483 85174 53517
rect 85208 53483 85220 53517
rect 85161 53459 85220 53483
rect 85921 53534 85978 53559
rect 85921 53500 85933 53534
rect 85967 53500 85978 53534
rect 85921 53475 85978 53500
rect 86078 53551 86157 53559
rect 86078 53517 86112 53551
rect 86146 53517 86157 53551
rect 86078 53475 86157 53517
rect 85161 53425 85261 53459
rect 85161 53391 85174 53425
rect 85208 53391 85261 53425
rect 85161 53375 85261 53391
rect 85361 53375 85403 53459
rect 85503 53434 85559 53459
rect 85503 53400 85514 53434
rect 85548 53400 85559 53434
rect 85503 53375 85559 53400
rect 85659 53375 85701 53459
rect 85801 53434 85858 53459
rect 86100 53451 86157 53475
rect 85801 53400 85812 53434
rect 85846 53400 85858 53434
rect 86100 53417 86112 53451
rect 86146 53417 86157 53451
rect 86100 53409 86157 53417
rect 86257 53551 86314 53559
rect 86257 53517 86268 53551
rect 86302 53517 86314 53551
rect 86257 53451 86314 53517
rect 86257 53417 86268 53451
rect 86302 53417 86314 53451
rect 86257 53409 86314 53417
rect 85801 53375 85858 53400
rect 1946 43052 2004 43406
rect 1946 42760 1958 43052
rect 1992 42760 2004 43052
rect 1946 42406 2004 42760
rect 3004 43052 3062 43406
rect 3004 42760 3016 43052
rect 3050 42760 3062 43052
rect 3004 42406 3062 42760
rect 4062 43052 4120 43406
rect 4062 42760 4074 43052
rect 4108 42760 4120 43052
rect 4062 42406 4120 42760
rect 5120 43052 5178 43406
rect 5120 42760 5132 43052
rect 5166 42760 5178 43052
rect 5120 42406 5178 42760
rect 6178 43052 6236 43406
rect 6178 42760 6190 43052
rect 6224 42760 6236 43052
rect 6178 42406 6236 42760
rect 7236 43052 7294 43406
rect 7236 42760 7248 43052
rect 7282 42760 7294 43052
rect 7236 42406 7294 42760
rect 8460 43060 8518 43414
rect 8460 42768 8472 43060
rect 8506 42768 8518 43060
rect 8460 42414 8518 42768
rect 9518 43060 9576 43414
rect 9518 42768 9530 43060
rect 9564 42768 9576 43060
rect 9518 42414 9576 42768
rect 10576 43060 10634 43414
rect 10576 42768 10588 43060
rect 10622 42768 10634 43060
rect 10576 42414 10634 42768
rect 11634 43060 11692 43414
rect 11634 42768 11646 43060
rect 11680 42768 11692 43060
rect 11634 42414 11692 42768
rect 12692 43060 12750 43414
rect 12692 42768 12704 43060
rect 12738 42768 12750 43060
rect 12692 42414 12750 42768
rect 13750 43060 13808 43414
rect 13750 42768 13762 43060
rect 13796 42768 13808 43060
rect 13750 42414 13808 42768
rect 14966 43068 15024 43422
rect 14966 42776 14978 43068
rect 15012 42776 15024 43068
rect 14966 42422 15024 42776
rect 16024 43068 16082 43422
rect 16024 42776 16036 43068
rect 16070 42776 16082 43068
rect 16024 42422 16082 42776
rect 17082 43068 17140 43422
rect 17082 42776 17094 43068
rect 17128 42776 17140 43068
rect 17082 42422 17140 42776
rect 18140 43068 18198 43422
rect 18140 42776 18152 43068
rect 18186 42776 18198 43068
rect 18140 42422 18198 42776
rect 19198 43068 19256 43422
rect 19198 42776 19210 43068
rect 19244 42776 19256 43068
rect 19198 42422 19256 42776
rect 20256 43068 20314 43422
rect 20256 42776 20268 43068
rect 20302 42776 20314 43068
rect 20256 42422 20314 42776
rect 21456 43052 21514 43406
rect 21456 42760 21468 43052
rect 21502 42760 21514 43052
rect 21456 42406 21514 42760
rect 22514 43052 22572 43406
rect 22514 42760 22526 43052
rect 22560 42760 22572 43052
rect 22514 42406 22572 42760
rect 23572 43052 23630 43406
rect 23572 42760 23584 43052
rect 23618 42760 23630 43052
rect 23572 42406 23630 42760
rect 24630 43052 24688 43406
rect 24630 42760 24642 43052
rect 24676 42760 24688 43052
rect 24630 42406 24688 42760
rect 25688 43052 25746 43406
rect 25688 42760 25700 43052
rect 25734 42760 25746 43052
rect 25688 42406 25746 42760
rect 26746 43052 26804 43406
rect 26746 42760 26758 43052
rect 26792 42760 26804 43052
rect 26746 42406 26804 42760
rect 27978 43068 28036 43422
rect 27978 42776 27990 43068
rect 28024 42776 28036 43068
rect 27978 42422 28036 42776
rect 29036 43068 29094 43422
rect 29036 42776 29048 43068
rect 29082 42776 29094 43068
rect 29036 42422 29094 42776
rect 30094 43068 30152 43422
rect 30094 42776 30106 43068
rect 30140 42776 30152 43068
rect 30094 42422 30152 42776
rect 31152 43068 31210 43422
rect 31152 42776 31164 43068
rect 31198 42776 31210 43068
rect 31152 42422 31210 42776
rect 32210 43068 32268 43422
rect 32210 42776 32222 43068
rect 32256 42776 32268 43068
rect 32210 42422 32268 42776
rect 33268 43068 33326 43422
rect 33268 42776 33280 43068
rect 33314 42776 33326 43068
rect 33268 42422 33326 42776
rect 34488 43074 34546 43428
rect 34488 42782 34500 43074
rect 34534 42782 34546 43074
rect 34488 42428 34546 42782
rect 35546 43074 35604 43428
rect 35546 42782 35558 43074
rect 35592 42782 35604 43074
rect 35546 42428 35604 42782
rect 36604 43074 36662 43428
rect 36604 42782 36616 43074
rect 36650 42782 36662 43074
rect 36604 42428 36662 42782
rect 37662 43074 37720 43428
rect 37662 42782 37674 43074
rect 37708 42782 37720 43074
rect 37662 42428 37720 42782
rect 38720 43074 38778 43428
rect 38720 42782 38732 43074
rect 38766 42782 38778 43074
rect 38720 42428 38778 42782
rect 39778 43074 39836 43428
rect 39778 42782 39790 43074
rect 39824 42782 39836 43074
rect 39778 42428 39836 42782
rect 40978 43074 41036 43428
rect 40978 42782 40990 43074
rect 41024 42782 41036 43074
rect 40978 42428 41036 42782
rect 42036 43074 42094 43428
rect 42036 42782 42048 43074
rect 42082 42782 42094 43074
rect 42036 42428 42094 42782
rect 43094 43074 43152 43428
rect 43094 42782 43106 43074
rect 43140 42782 43152 43074
rect 43094 42428 43152 42782
rect 44152 43074 44210 43428
rect 44152 42782 44164 43074
rect 44198 42782 44210 43074
rect 44152 42428 44210 42782
rect 45210 43074 45268 43428
rect 45210 42782 45222 43074
rect 45256 42782 45268 43074
rect 45210 42428 45268 42782
rect 46268 43074 46326 43428
rect 46268 42782 46280 43074
rect 46314 42782 46326 43074
rect 46268 42428 46326 42782
rect 47566 43096 47624 43450
rect 47566 42804 47578 43096
rect 47612 42804 47624 43096
rect 47566 42450 47624 42804
rect 48624 43096 48682 43450
rect 48624 42804 48636 43096
rect 48670 42804 48682 43096
rect 48624 42450 48682 42804
rect 49682 43096 49740 43450
rect 49682 42804 49694 43096
rect 49728 42804 49740 43096
rect 49682 42450 49740 42804
rect 50740 43096 50798 43450
rect 50740 42804 50752 43096
rect 50786 42804 50798 43096
rect 50740 42450 50798 42804
rect 51798 43096 51856 43450
rect 51798 42804 51810 43096
rect 51844 42804 51856 43096
rect 51798 42450 51856 42804
rect 52856 43096 52914 43450
rect 52856 42804 52868 43096
rect 52902 42804 52914 43096
rect 52856 42450 52914 42804
rect 54080 43110 54138 43464
rect 54080 42818 54092 43110
rect 54126 42818 54138 43110
rect 54080 42464 54138 42818
rect 55138 43110 55196 43464
rect 55138 42818 55150 43110
rect 55184 42818 55196 43110
rect 55138 42464 55196 42818
rect 56196 43110 56254 43464
rect 56196 42818 56208 43110
rect 56242 42818 56254 43110
rect 56196 42464 56254 42818
rect 57254 43110 57312 43464
rect 57254 42818 57266 43110
rect 57300 42818 57312 43110
rect 57254 42464 57312 42818
rect 58312 43110 58370 43464
rect 58312 42818 58324 43110
rect 58358 42818 58370 43110
rect 58312 42464 58370 42818
rect 59370 43110 59428 43464
rect 59370 42818 59382 43110
rect 59416 42818 59428 43110
rect 59370 42464 59428 42818
rect 1946 41958 2004 42312
rect 1946 41666 1958 41958
rect 1992 41666 2004 41958
rect 1946 41312 2004 41666
rect 3004 41958 3062 42312
rect 3004 41666 3016 41958
rect 3050 41666 3062 41958
rect 3004 41312 3062 41666
rect 4062 41958 4120 42312
rect 4062 41666 4074 41958
rect 4108 41666 4120 41958
rect 4062 41312 4120 41666
rect 5120 41958 5178 42312
rect 5120 41666 5132 41958
rect 5166 41666 5178 41958
rect 5120 41312 5178 41666
rect 6178 41958 6236 42312
rect 6178 41666 6190 41958
rect 6224 41666 6236 41958
rect 6178 41312 6236 41666
rect 7236 41958 7294 42312
rect 7236 41666 7248 41958
rect 7282 41666 7294 41958
rect 8460 41966 8518 42320
rect 7236 41312 7294 41666
rect 1946 40864 2004 41218
rect 1946 40572 1958 40864
rect 1992 40572 2004 40864
rect 1946 40218 2004 40572
rect 3004 40864 3062 41218
rect 3004 40572 3016 40864
rect 3050 40572 3062 40864
rect 3004 40218 3062 40572
rect 4062 40864 4120 41218
rect 4062 40572 4074 40864
rect 4108 40572 4120 40864
rect 4062 40218 4120 40572
rect 5120 40864 5178 41218
rect 5120 40572 5132 40864
rect 5166 40572 5178 40864
rect 5120 40218 5178 40572
rect 6178 40864 6236 41218
rect 6178 40572 6190 40864
rect 6224 40572 6236 40864
rect 6178 40218 6236 40572
rect 7236 40864 7294 41218
rect 7236 40572 7248 40864
rect 7282 40572 7294 40864
rect 7236 40218 7294 40572
rect 8460 41674 8472 41966
rect 8506 41674 8518 41966
rect 8460 41320 8518 41674
rect 9518 41966 9576 42320
rect 9518 41674 9530 41966
rect 9564 41674 9576 41966
rect 9518 41320 9576 41674
rect 10576 41966 10634 42320
rect 10576 41674 10588 41966
rect 10622 41674 10634 41966
rect 10576 41320 10634 41674
rect 11634 41966 11692 42320
rect 11634 41674 11646 41966
rect 11680 41674 11692 41966
rect 11634 41320 11692 41674
rect 12692 41966 12750 42320
rect 12692 41674 12704 41966
rect 12738 41674 12750 41966
rect 12692 41320 12750 41674
rect 13750 41966 13808 42320
rect 13750 41674 13762 41966
rect 13796 41674 13808 41966
rect 14966 41974 15024 42328
rect 13750 41320 13808 41674
rect 1946 39770 2004 40124
rect 1946 39478 1958 39770
rect 1992 39478 2004 39770
rect 1946 39124 2004 39478
rect 3004 39770 3062 40124
rect 3004 39478 3016 39770
rect 3050 39478 3062 39770
rect 3004 39124 3062 39478
rect 4062 39770 4120 40124
rect 4062 39478 4074 39770
rect 4108 39478 4120 39770
rect 4062 39124 4120 39478
rect 5120 39770 5178 40124
rect 5120 39478 5132 39770
rect 5166 39478 5178 39770
rect 5120 39124 5178 39478
rect 6178 39770 6236 40124
rect 6178 39478 6190 39770
rect 6224 39478 6236 39770
rect 6178 39124 6236 39478
rect 7236 39770 7294 40124
rect 8460 40872 8518 41226
rect 8460 40580 8472 40872
rect 8506 40580 8518 40872
rect 8460 40226 8518 40580
rect 9518 40872 9576 41226
rect 9518 40580 9530 40872
rect 9564 40580 9576 40872
rect 9518 40226 9576 40580
rect 10576 40872 10634 41226
rect 10576 40580 10588 40872
rect 10622 40580 10634 40872
rect 10576 40226 10634 40580
rect 11634 40872 11692 41226
rect 11634 40580 11646 40872
rect 11680 40580 11692 40872
rect 11634 40226 11692 40580
rect 12692 40872 12750 41226
rect 12692 40580 12704 40872
rect 12738 40580 12750 40872
rect 12692 40226 12750 40580
rect 13750 40872 13808 41226
rect 13750 40580 13762 40872
rect 13796 40580 13808 40872
rect 13750 40226 13808 40580
rect 14966 41682 14978 41974
rect 15012 41682 15024 41974
rect 14966 41328 15024 41682
rect 16024 41974 16082 42328
rect 16024 41682 16036 41974
rect 16070 41682 16082 41974
rect 16024 41328 16082 41682
rect 17082 41974 17140 42328
rect 17082 41682 17094 41974
rect 17128 41682 17140 41974
rect 17082 41328 17140 41682
rect 18140 41974 18198 42328
rect 18140 41682 18152 41974
rect 18186 41682 18198 41974
rect 18140 41328 18198 41682
rect 19198 41974 19256 42328
rect 19198 41682 19210 41974
rect 19244 41682 19256 41974
rect 19198 41328 19256 41682
rect 20256 41974 20314 42328
rect 20256 41682 20268 41974
rect 20302 41682 20314 41974
rect 20256 41328 20314 41682
rect 21456 41958 21514 42312
rect 7236 39478 7248 39770
rect 7282 39478 7294 39770
rect 7236 39124 7294 39478
rect 8460 39778 8518 40132
rect 8460 39486 8472 39778
rect 8506 39486 8518 39778
rect 8460 39132 8518 39486
rect 9518 39778 9576 40132
rect 9518 39486 9530 39778
rect 9564 39486 9576 39778
rect 9518 39132 9576 39486
rect 10576 39778 10634 40132
rect 10576 39486 10588 39778
rect 10622 39486 10634 39778
rect 10576 39132 10634 39486
rect 11634 39778 11692 40132
rect 11634 39486 11646 39778
rect 11680 39486 11692 39778
rect 11634 39132 11692 39486
rect 12692 39778 12750 40132
rect 12692 39486 12704 39778
rect 12738 39486 12750 39778
rect 12692 39132 12750 39486
rect 13750 39778 13808 40132
rect 14966 40880 15024 41234
rect 14966 40588 14978 40880
rect 15012 40588 15024 40880
rect 14966 40234 15024 40588
rect 16024 40880 16082 41234
rect 16024 40588 16036 40880
rect 16070 40588 16082 40880
rect 16024 40234 16082 40588
rect 17082 40880 17140 41234
rect 17082 40588 17094 40880
rect 17128 40588 17140 40880
rect 17082 40234 17140 40588
rect 18140 40880 18198 41234
rect 18140 40588 18152 40880
rect 18186 40588 18198 40880
rect 18140 40234 18198 40588
rect 19198 40880 19256 41234
rect 19198 40588 19210 40880
rect 19244 40588 19256 40880
rect 19198 40234 19256 40588
rect 20256 40880 20314 41234
rect 20256 40588 20268 40880
rect 20302 40588 20314 40880
rect 20256 40234 20314 40588
rect 21456 41666 21468 41958
rect 21502 41666 21514 41958
rect 21456 41312 21514 41666
rect 22514 41958 22572 42312
rect 22514 41666 22526 41958
rect 22560 41666 22572 41958
rect 22514 41312 22572 41666
rect 23572 41958 23630 42312
rect 23572 41666 23584 41958
rect 23618 41666 23630 41958
rect 23572 41312 23630 41666
rect 24630 41958 24688 42312
rect 24630 41666 24642 41958
rect 24676 41666 24688 41958
rect 24630 41312 24688 41666
rect 25688 41958 25746 42312
rect 25688 41666 25700 41958
rect 25734 41666 25746 41958
rect 25688 41312 25746 41666
rect 26746 41958 26804 42312
rect 26746 41666 26758 41958
rect 26792 41666 26804 41958
rect 27978 41974 28036 42328
rect 26746 41312 26804 41666
rect 13750 39486 13762 39778
rect 13796 39486 13808 39778
rect 13750 39132 13808 39486
rect 14966 39786 15024 40140
rect 14966 39494 14978 39786
rect 15012 39494 15024 39786
rect 14966 39140 15024 39494
rect 16024 39786 16082 40140
rect 16024 39494 16036 39786
rect 16070 39494 16082 39786
rect 16024 39140 16082 39494
rect 17082 39786 17140 40140
rect 17082 39494 17094 39786
rect 17128 39494 17140 39786
rect 17082 39140 17140 39494
rect 18140 39786 18198 40140
rect 18140 39494 18152 39786
rect 18186 39494 18198 39786
rect 18140 39140 18198 39494
rect 19198 39786 19256 40140
rect 19198 39494 19210 39786
rect 19244 39494 19256 39786
rect 19198 39140 19256 39494
rect 20256 39786 20314 40140
rect 21456 40864 21514 41218
rect 21456 40572 21468 40864
rect 21502 40572 21514 40864
rect 21456 40218 21514 40572
rect 22514 40864 22572 41218
rect 22514 40572 22526 40864
rect 22560 40572 22572 40864
rect 22514 40218 22572 40572
rect 23572 40864 23630 41218
rect 23572 40572 23584 40864
rect 23618 40572 23630 40864
rect 23572 40218 23630 40572
rect 24630 40864 24688 41218
rect 24630 40572 24642 40864
rect 24676 40572 24688 40864
rect 24630 40218 24688 40572
rect 25688 40864 25746 41218
rect 25688 40572 25700 40864
rect 25734 40572 25746 40864
rect 25688 40218 25746 40572
rect 26746 40864 26804 41218
rect 26746 40572 26758 40864
rect 26792 40572 26804 40864
rect 26746 40218 26804 40572
rect 27978 41682 27990 41974
rect 28024 41682 28036 41974
rect 27978 41328 28036 41682
rect 29036 41974 29094 42328
rect 29036 41682 29048 41974
rect 29082 41682 29094 41974
rect 29036 41328 29094 41682
rect 30094 41974 30152 42328
rect 30094 41682 30106 41974
rect 30140 41682 30152 41974
rect 30094 41328 30152 41682
rect 31152 41974 31210 42328
rect 31152 41682 31164 41974
rect 31198 41682 31210 41974
rect 31152 41328 31210 41682
rect 32210 41974 32268 42328
rect 32210 41682 32222 41974
rect 32256 41682 32268 41974
rect 32210 41328 32268 41682
rect 33268 41974 33326 42328
rect 33268 41682 33280 41974
rect 33314 41682 33326 41974
rect 34488 41980 34546 42334
rect 33268 41328 33326 41682
rect 20256 39494 20268 39786
rect 20302 39494 20314 39786
rect 20256 39140 20314 39494
rect 21456 39770 21514 40124
rect 21456 39478 21468 39770
rect 21502 39478 21514 39770
rect 21456 39124 21514 39478
rect 22514 39770 22572 40124
rect 22514 39478 22526 39770
rect 22560 39478 22572 39770
rect 22514 39124 22572 39478
rect 23572 39770 23630 40124
rect 23572 39478 23584 39770
rect 23618 39478 23630 39770
rect 23572 39124 23630 39478
rect 24630 39770 24688 40124
rect 24630 39478 24642 39770
rect 24676 39478 24688 39770
rect 24630 39124 24688 39478
rect 25688 39770 25746 40124
rect 25688 39478 25700 39770
rect 25734 39478 25746 39770
rect 25688 39124 25746 39478
rect 26746 39770 26804 40124
rect 27978 40880 28036 41234
rect 27978 40588 27990 40880
rect 28024 40588 28036 40880
rect 27978 40234 28036 40588
rect 29036 40880 29094 41234
rect 29036 40588 29048 40880
rect 29082 40588 29094 40880
rect 29036 40234 29094 40588
rect 30094 40880 30152 41234
rect 30094 40588 30106 40880
rect 30140 40588 30152 40880
rect 30094 40234 30152 40588
rect 31152 40880 31210 41234
rect 31152 40588 31164 40880
rect 31198 40588 31210 40880
rect 31152 40234 31210 40588
rect 32210 40880 32268 41234
rect 32210 40588 32222 40880
rect 32256 40588 32268 40880
rect 32210 40234 32268 40588
rect 33268 40880 33326 41234
rect 33268 40588 33280 40880
rect 33314 40588 33326 40880
rect 33268 40234 33326 40588
rect 34488 41688 34500 41980
rect 34534 41688 34546 41980
rect 34488 41334 34546 41688
rect 35546 41980 35604 42334
rect 35546 41688 35558 41980
rect 35592 41688 35604 41980
rect 35546 41334 35604 41688
rect 36604 41980 36662 42334
rect 36604 41688 36616 41980
rect 36650 41688 36662 41980
rect 36604 41334 36662 41688
rect 37662 41980 37720 42334
rect 37662 41688 37674 41980
rect 37708 41688 37720 41980
rect 37662 41334 37720 41688
rect 38720 41980 38778 42334
rect 38720 41688 38732 41980
rect 38766 41688 38778 41980
rect 38720 41334 38778 41688
rect 39778 41980 39836 42334
rect 39778 41688 39790 41980
rect 39824 41688 39836 41980
rect 40978 41980 41036 42334
rect 39778 41334 39836 41688
rect 26746 39478 26758 39770
rect 26792 39478 26804 39770
rect 26746 39124 26804 39478
rect 27978 39786 28036 40140
rect 27978 39494 27990 39786
rect 28024 39494 28036 39786
rect 27978 39140 28036 39494
rect 29036 39786 29094 40140
rect 29036 39494 29048 39786
rect 29082 39494 29094 39786
rect 29036 39140 29094 39494
rect 30094 39786 30152 40140
rect 30094 39494 30106 39786
rect 30140 39494 30152 39786
rect 30094 39140 30152 39494
rect 31152 39786 31210 40140
rect 31152 39494 31164 39786
rect 31198 39494 31210 39786
rect 31152 39140 31210 39494
rect 32210 39786 32268 40140
rect 32210 39494 32222 39786
rect 32256 39494 32268 39786
rect 32210 39140 32268 39494
rect 33268 39786 33326 40140
rect 34488 40886 34546 41240
rect 34488 40594 34500 40886
rect 34534 40594 34546 40886
rect 34488 40240 34546 40594
rect 35546 40886 35604 41240
rect 35546 40594 35558 40886
rect 35592 40594 35604 40886
rect 35546 40240 35604 40594
rect 36604 40886 36662 41240
rect 36604 40594 36616 40886
rect 36650 40594 36662 40886
rect 36604 40240 36662 40594
rect 37662 40886 37720 41240
rect 37662 40594 37674 40886
rect 37708 40594 37720 40886
rect 37662 40240 37720 40594
rect 38720 40886 38778 41240
rect 38720 40594 38732 40886
rect 38766 40594 38778 40886
rect 38720 40240 38778 40594
rect 39778 40886 39836 41240
rect 39778 40594 39790 40886
rect 39824 40594 39836 40886
rect 39778 40240 39836 40594
rect 40978 41688 40990 41980
rect 41024 41688 41036 41980
rect 40978 41334 41036 41688
rect 42036 41980 42094 42334
rect 42036 41688 42048 41980
rect 42082 41688 42094 41980
rect 42036 41334 42094 41688
rect 43094 41980 43152 42334
rect 43094 41688 43106 41980
rect 43140 41688 43152 41980
rect 43094 41334 43152 41688
rect 44152 41980 44210 42334
rect 44152 41688 44164 41980
rect 44198 41688 44210 41980
rect 44152 41334 44210 41688
rect 45210 41980 45268 42334
rect 45210 41688 45222 41980
rect 45256 41688 45268 41980
rect 45210 41334 45268 41688
rect 46268 41980 46326 42334
rect 46268 41688 46280 41980
rect 46314 41688 46326 41980
rect 47566 42002 47624 42356
rect 46268 41334 46326 41688
rect 33268 39494 33280 39786
rect 33314 39494 33326 39786
rect 33268 39140 33326 39494
rect 34488 39792 34546 40146
rect 34488 39500 34500 39792
rect 34534 39500 34546 39792
rect 34488 39146 34546 39500
rect 35546 39792 35604 40146
rect 35546 39500 35558 39792
rect 35592 39500 35604 39792
rect 35546 39146 35604 39500
rect 36604 39792 36662 40146
rect 36604 39500 36616 39792
rect 36650 39500 36662 39792
rect 36604 39146 36662 39500
rect 37662 39792 37720 40146
rect 37662 39500 37674 39792
rect 37708 39500 37720 39792
rect 37662 39146 37720 39500
rect 38720 39792 38778 40146
rect 38720 39500 38732 39792
rect 38766 39500 38778 39792
rect 38720 39146 38778 39500
rect 39778 39792 39836 40146
rect 40978 40886 41036 41240
rect 40978 40594 40990 40886
rect 41024 40594 41036 40886
rect 40978 40240 41036 40594
rect 42036 40886 42094 41240
rect 42036 40594 42048 40886
rect 42082 40594 42094 40886
rect 42036 40240 42094 40594
rect 43094 40886 43152 41240
rect 43094 40594 43106 40886
rect 43140 40594 43152 40886
rect 43094 40240 43152 40594
rect 44152 40886 44210 41240
rect 44152 40594 44164 40886
rect 44198 40594 44210 40886
rect 44152 40240 44210 40594
rect 45210 40886 45268 41240
rect 45210 40594 45222 40886
rect 45256 40594 45268 40886
rect 45210 40240 45268 40594
rect 46268 40886 46326 41240
rect 46268 40594 46280 40886
rect 46314 40594 46326 40886
rect 46268 40240 46326 40594
rect 47566 41710 47578 42002
rect 47612 41710 47624 42002
rect 47566 41356 47624 41710
rect 48624 42002 48682 42356
rect 48624 41710 48636 42002
rect 48670 41710 48682 42002
rect 48624 41356 48682 41710
rect 49682 42002 49740 42356
rect 49682 41710 49694 42002
rect 49728 41710 49740 42002
rect 49682 41356 49740 41710
rect 50740 42002 50798 42356
rect 50740 41710 50752 42002
rect 50786 41710 50798 42002
rect 50740 41356 50798 41710
rect 51798 42002 51856 42356
rect 51798 41710 51810 42002
rect 51844 41710 51856 42002
rect 51798 41356 51856 41710
rect 52856 42002 52914 42356
rect 52856 41710 52868 42002
rect 52902 41710 52914 42002
rect 54080 42016 54138 42370
rect 52856 41356 52914 41710
rect 39778 39500 39790 39792
rect 39824 39500 39836 39792
rect 39778 39146 39836 39500
rect 40978 39792 41036 40146
rect 40978 39500 40990 39792
rect 41024 39500 41036 39792
rect 40978 39146 41036 39500
rect 42036 39792 42094 40146
rect 42036 39500 42048 39792
rect 42082 39500 42094 39792
rect 42036 39146 42094 39500
rect 43094 39792 43152 40146
rect 43094 39500 43106 39792
rect 43140 39500 43152 39792
rect 43094 39146 43152 39500
rect 44152 39792 44210 40146
rect 44152 39500 44164 39792
rect 44198 39500 44210 39792
rect 44152 39146 44210 39500
rect 45210 39792 45268 40146
rect 45210 39500 45222 39792
rect 45256 39500 45268 39792
rect 45210 39146 45268 39500
rect 46268 39792 46326 40146
rect 47566 40908 47624 41262
rect 47566 40616 47578 40908
rect 47612 40616 47624 40908
rect 47566 40262 47624 40616
rect 48624 40908 48682 41262
rect 48624 40616 48636 40908
rect 48670 40616 48682 40908
rect 48624 40262 48682 40616
rect 49682 40908 49740 41262
rect 49682 40616 49694 40908
rect 49728 40616 49740 40908
rect 49682 40262 49740 40616
rect 50740 40908 50798 41262
rect 50740 40616 50752 40908
rect 50786 40616 50798 40908
rect 50740 40262 50798 40616
rect 51798 40908 51856 41262
rect 51798 40616 51810 40908
rect 51844 40616 51856 40908
rect 51798 40262 51856 40616
rect 52856 40908 52914 41262
rect 52856 40616 52868 40908
rect 52902 40616 52914 40908
rect 52856 40262 52914 40616
rect 54080 41724 54092 42016
rect 54126 41724 54138 42016
rect 54080 41370 54138 41724
rect 55138 42016 55196 42370
rect 55138 41724 55150 42016
rect 55184 41724 55196 42016
rect 55138 41370 55196 41724
rect 56196 42016 56254 42370
rect 56196 41724 56208 42016
rect 56242 41724 56254 42016
rect 56196 41370 56254 41724
rect 57254 42016 57312 42370
rect 57254 41724 57266 42016
rect 57300 41724 57312 42016
rect 57254 41370 57312 41724
rect 58312 42016 58370 42370
rect 58312 41724 58324 42016
rect 58358 41724 58370 42016
rect 58312 41370 58370 41724
rect 59370 42016 59428 42370
rect 59370 41724 59382 42016
rect 59416 41724 59428 42016
rect 59370 41370 59428 41724
rect 46268 39500 46280 39792
rect 46314 39500 46326 39792
rect 46268 39146 46326 39500
rect 47566 39814 47624 40168
rect 47566 39522 47578 39814
rect 47612 39522 47624 39814
rect 47566 39168 47624 39522
rect 48624 39814 48682 40168
rect 48624 39522 48636 39814
rect 48670 39522 48682 39814
rect 48624 39168 48682 39522
rect 49682 39814 49740 40168
rect 49682 39522 49694 39814
rect 49728 39522 49740 39814
rect 49682 39168 49740 39522
rect 50740 39814 50798 40168
rect 50740 39522 50752 39814
rect 50786 39522 50798 39814
rect 50740 39168 50798 39522
rect 51798 39814 51856 40168
rect 51798 39522 51810 39814
rect 51844 39522 51856 39814
rect 51798 39168 51856 39522
rect 52856 39814 52914 40168
rect 54080 40922 54138 41276
rect 54080 40630 54092 40922
rect 54126 40630 54138 40922
rect 54080 40276 54138 40630
rect 55138 40922 55196 41276
rect 55138 40630 55150 40922
rect 55184 40630 55196 40922
rect 55138 40276 55196 40630
rect 56196 40922 56254 41276
rect 56196 40630 56208 40922
rect 56242 40630 56254 40922
rect 56196 40276 56254 40630
rect 57254 40922 57312 41276
rect 57254 40630 57266 40922
rect 57300 40630 57312 40922
rect 57254 40276 57312 40630
rect 58312 40922 58370 41276
rect 58312 40630 58324 40922
rect 58358 40630 58370 40922
rect 58312 40276 58370 40630
rect 59370 40922 59428 41276
rect 59370 40630 59382 40922
rect 59416 40630 59428 40922
rect 59370 40276 59428 40630
rect 52856 39522 52868 39814
rect 52902 39522 52914 39814
rect 52856 39168 52914 39522
rect 54080 39828 54138 40182
rect 54080 39536 54092 39828
rect 54126 39536 54138 39828
rect 54080 39182 54138 39536
rect 55138 39828 55196 40182
rect 55138 39536 55150 39828
rect 55184 39536 55196 39828
rect 55138 39182 55196 39536
rect 56196 39828 56254 40182
rect 56196 39536 56208 39828
rect 56242 39536 56254 39828
rect 56196 39182 56254 39536
rect 57254 39828 57312 40182
rect 57254 39536 57266 39828
rect 57300 39536 57312 39828
rect 57254 39182 57312 39536
rect 58312 39828 58370 40182
rect 58312 39536 58324 39828
rect 58358 39536 58370 39828
rect 58312 39182 58370 39536
rect 59370 39828 59428 40182
rect 59370 39536 59382 39828
rect 59416 39536 59428 39828
rect 59370 39182 59428 39536
rect 1946 38676 2004 39030
rect 1946 38384 1958 38676
rect 1992 38384 2004 38676
rect 1946 38030 2004 38384
rect 3004 38676 3062 39030
rect 3004 38384 3016 38676
rect 3050 38384 3062 38676
rect 3004 38030 3062 38384
rect 4062 38676 4120 39030
rect 4062 38384 4074 38676
rect 4108 38384 4120 38676
rect 4062 38030 4120 38384
rect 5120 38676 5178 39030
rect 5120 38384 5132 38676
rect 5166 38384 5178 38676
rect 5120 38030 5178 38384
rect 6178 38676 6236 39030
rect 6178 38384 6190 38676
rect 6224 38384 6236 38676
rect 6178 38030 6236 38384
rect 7236 38676 7294 39030
rect 7236 38384 7248 38676
rect 7282 38384 7294 38676
rect 7236 38030 7294 38384
rect 8460 38684 8518 39038
rect 8460 38392 8472 38684
rect 8506 38392 8518 38684
rect 8460 38038 8518 38392
rect 9518 38684 9576 39038
rect 9518 38392 9530 38684
rect 9564 38392 9576 38684
rect 9518 38038 9576 38392
rect 10576 38684 10634 39038
rect 10576 38392 10588 38684
rect 10622 38392 10634 38684
rect 10576 38038 10634 38392
rect 11634 38684 11692 39038
rect 11634 38392 11646 38684
rect 11680 38392 11692 38684
rect 11634 38038 11692 38392
rect 12692 38684 12750 39038
rect 12692 38392 12704 38684
rect 12738 38392 12750 38684
rect 12692 38038 12750 38392
rect 13750 38684 13808 39038
rect 13750 38392 13762 38684
rect 13796 38392 13808 38684
rect 13750 38038 13808 38392
rect 14966 38692 15024 39046
rect 14966 38400 14978 38692
rect 15012 38400 15024 38692
rect 14966 38046 15024 38400
rect 16024 38692 16082 39046
rect 16024 38400 16036 38692
rect 16070 38400 16082 38692
rect 16024 38046 16082 38400
rect 17082 38692 17140 39046
rect 17082 38400 17094 38692
rect 17128 38400 17140 38692
rect 17082 38046 17140 38400
rect 18140 38692 18198 39046
rect 18140 38400 18152 38692
rect 18186 38400 18198 38692
rect 18140 38046 18198 38400
rect 19198 38692 19256 39046
rect 19198 38400 19210 38692
rect 19244 38400 19256 38692
rect 19198 38046 19256 38400
rect 20256 38692 20314 39046
rect 20256 38400 20268 38692
rect 20302 38400 20314 38692
rect 20256 38046 20314 38400
rect 21456 38676 21514 39030
rect 21456 38384 21468 38676
rect 21502 38384 21514 38676
rect 21456 38030 21514 38384
rect 22514 38676 22572 39030
rect 22514 38384 22526 38676
rect 22560 38384 22572 38676
rect 22514 38030 22572 38384
rect 23572 38676 23630 39030
rect 23572 38384 23584 38676
rect 23618 38384 23630 38676
rect 23572 38030 23630 38384
rect 24630 38676 24688 39030
rect 24630 38384 24642 38676
rect 24676 38384 24688 38676
rect 24630 38030 24688 38384
rect 25688 38676 25746 39030
rect 25688 38384 25700 38676
rect 25734 38384 25746 38676
rect 25688 38030 25746 38384
rect 26746 38676 26804 39030
rect 26746 38384 26758 38676
rect 26792 38384 26804 38676
rect 26746 38030 26804 38384
rect 27978 38692 28036 39046
rect 27978 38400 27990 38692
rect 28024 38400 28036 38692
rect 27978 38046 28036 38400
rect 29036 38692 29094 39046
rect 29036 38400 29048 38692
rect 29082 38400 29094 38692
rect 29036 38046 29094 38400
rect 30094 38692 30152 39046
rect 30094 38400 30106 38692
rect 30140 38400 30152 38692
rect 30094 38046 30152 38400
rect 31152 38692 31210 39046
rect 31152 38400 31164 38692
rect 31198 38400 31210 38692
rect 31152 38046 31210 38400
rect 32210 38692 32268 39046
rect 32210 38400 32222 38692
rect 32256 38400 32268 38692
rect 32210 38046 32268 38400
rect 33268 38692 33326 39046
rect 33268 38400 33280 38692
rect 33314 38400 33326 38692
rect 33268 38046 33326 38400
rect 34488 38698 34546 39052
rect 34488 38406 34500 38698
rect 34534 38406 34546 38698
rect 34488 38052 34546 38406
rect 35546 38698 35604 39052
rect 35546 38406 35558 38698
rect 35592 38406 35604 38698
rect 35546 38052 35604 38406
rect 36604 38698 36662 39052
rect 36604 38406 36616 38698
rect 36650 38406 36662 38698
rect 36604 38052 36662 38406
rect 37662 38698 37720 39052
rect 37662 38406 37674 38698
rect 37708 38406 37720 38698
rect 37662 38052 37720 38406
rect 38720 38698 38778 39052
rect 38720 38406 38732 38698
rect 38766 38406 38778 38698
rect 38720 38052 38778 38406
rect 39778 38698 39836 39052
rect 39778 38406 39790 38698
rect 39824 38406 39836 38698
rect 39778 38052 39836 38406
rect 40978 38698 41036 39052
rect 40978 38406 40990 38698
rect 41024 38406 41036 38698
rect 40978 38052 41036 38406
rect 42036 38698 42094 39052
rect 42036 38406 42048 38698
rect 42082 38406 42094 38698
rect 42036 38052 42094 38406
rect 43094 38698 43152 39052
rect 43094 38406 43106 38698
rect 43140 38406 43152 38698
rect 43094 38052 43152 38406
rect 44152 38698 44210 39052
rect 44152 38406 44164 38698
rect 44198 38406 44210 38698
rect 44152 38052 44210 38406
rect 45210 38698 45268 39052
rect 45210 38406 45222 38698
rect 45256 38406 45268 38698
rect 45210 38052 45268 38406
rect 46268 38698 46326 39052
rect 46268 38406 46280 38698
rect 46314 38406 46326 38698
rect 46268 38052 46326 38406
rect 47566 38720 47624 39074
rect 47566 38428 47578 38720
rect 47612 38428 47624 38720
rect 47566 38074 47624 38428
rect 48624 38720 48682 39074
rect 48624 38428 48636 38720
rect 48670 38428 48682 38720
rect 48624 38074 48682 38428
rect 49682 38720 49740 39074
rect 49682 38428 49694 38720
rect 49728 38428 49740 38720
rect 49682 38074 49740 38428
rect 50740 38720 50798 39074
rect 50740 38428 50752 38720
rect 50786 38428 50798 38720
rect 50740 38074 50798 38428
rect 51798 38720 51856 39074
rect 51798 38428 51810 38720
rect 51844 38428 51856 38720
rect 51798 38074 51856 38428
rect 52856 38720 52914 39074
rect 52856 38428 52868 38720
rect 52902 38428 52914 38720
rect 52856 38074 52914 38428
rect 54080 38734 54138 39088
rect 54080 38442 54092 38734
rect 54126 38442 54138 38734
rect 54080 38088 54138 38442
rect 55138 38734 55196 39088
rect 55138 38442 55150 38734
rect 55184 38442 55196 38734
rect 55138 38088 55196 38442
rect 56196 38734 56254 39088
rect 56196 38442 56208 38734
rect 56242 38442 56254 38734
rect 56196 38088 56254 38442
rect 57254 38734 57312 39088
rect 57254 38442 57266 38734
rect 57300 38442 57312 38734
rect 57254 38088 57312 38442
rect 58312 38734 58370 39088
rect 58312 38442 58324 38734
rect 58358 38442 58370 38734
rect 58312 38088 58370 38442
rect 59370 38734 59428 39088
rect 59370 38442 59382 38734
rect 59416 38442 59428 38734
rect 59370 38088 59428 38442
rect 1946 37236 2004 37590
rect 1946 36944 1958 37236
rect 1992 36944 2004 37236
rect 1946 36590 2004 36944
rect 3004 37236 3062 37590
rect 3004 36944 3016 37236
rect 3050 36944 3062 37236
rect 3004 36590 3062 36944
rect 4062 37236 4120 37590
rect 4062 36944 4074 37236
rect 4108 36944 4120 37236
rect 4062 36590 4120 36944
rect 5120 37236 5178 37590
rect 5120 36944 5132 37236
rect 5166 36944 5178 37236
rect 5120 36590 5178 36944
rect 6178 37236 6236 37590
rect 6178 36944 6190 37236
rect 6224 36944 6236 37236
rect 6178 36590 6236 36944
rect 7236 37236 7294 37590
rect 7236 36944 7248 37236
rect 7282 36944 7294 37236
rect 7236 36590 7294 36944
rect 8460 37244 8518 37598
rect 8460 36952 8472 37244
rect 8506 36952 8518 37244
rect 8460 36598 8518 36952
rect 9518 37244 9576 37598
rect 9518 36952 9530 37244
rect 9564 36952 9576 37244
rect 9518 36598 9576 36952
rect 10576 37244 10634 37598
rect 10576 36952 10588 37244
rect 10622 36952 10634 37244
rect 10576 36598 10634 36952
rect 11634 37244 11692 37598
rect 11634 36952 11646 37244
rect 11680 36952 11692 37244
rect 11634 36598 11692 36952
rect 12692 37244 12750 37598
rect 12692 36952 12704 37244
rect 12738 36952 12750 37244
rect 12692 36598 12750 36952
rect 13750 37244 13808 37598
rect 13750 36952 13762 37244
rect 13796 36952 13808 37244
rect 13750 36598 13808 36952
rect 14966 37252 15024 37606
rect 14966 36960 14978 37252
rect 15012 36960 15024 37252
rect 14966 36606 15024 36960
rect 16024 37252 16082 37606
rect 16024 36960 16036 37252
rect 16070 36960 16082 37252
rect 16024 36606 16082 36960
rect 17082 37252 17140 37606
rect 17082 36960 17094 37252
rect 17128 36960 17140 37252
rect 17082 36606 17140 36960
rect 18140 37252 18198 37606
rect 18140 36960 18152 37252
rect 18186 36960 18198 37252
rect 18140 36606 18198 36960
rect 19198 37252 19256 37606
rect 19198 36960 19210 37252
rect 19244 36960 19256 37252
rect 19198 36606 19256 36960
rect 20256 37252 20314 37606
rect 20256 36960 20268 37252
rect 20302 36960 20314 37252
rect 20256 36606 20314 36960
rect 21456 37236 21514 37590
rect 21456 36944 21468 37236
rect 21502 36944 21514 37236
rect 21456 36590 21514 36944
rect 22514 37236 22572 37590
rect 22514 36944 22526 37236
rect 22560 36944 22572 37236
rect 22514 36590 22572 36944
rect 23572 37236 23630 37590
rect 23572 36944 23584 37236
rect 23618 36944 23630 37236
rect 23572 36590 23630 36944
rect 24630 37236 24688 37590
rect 24630 36944 24642 37236
rect 24676 36944 24688 37236
rect 24630 36590 24688 36944
rect 25688 37236 25746 37590
rect 25688 36944 25700 37236
rect 25734 36944 25746 37236
rect 25688 36590 25746 36944
rect 26746 37236 26804 37590
rect 26746 36944 26758 37236
rect 26792 36944 26804 37236
rect 26746 36590 26804 36944
rect 27978 37252 28036 37606
rect 27978 36960 27990 37252
rect 28024 36960 28036 37252
rect 27978 36606 28036 36960
rect 29036 37252 29094 37606
rect 29036 36960 29048 37252
rect 29082 36960 29094 37252
rect 29036 36606 29094 36960
rect 30094 37252 30152 37606
rect 30094 36960 30106 37252
rect 30140 36960 30152 37252
rect 30094 36606 30152 36960
rect 31152 37252 31210 37606
rect 31152 36960 31164 37252
rect 31198 36960 31210 37252
rect 31152 36606 31210 36960
rect 32210 37252 32268 37606
rect 32210 36960 32222 37252
rect 32256 36960 32268 37252
rect 32210 36606 32268 36960
rect 33268 37252 33326 37606
rect 33268 36960 33280 37252
rect 33314 36960 33326 37252
rect 33268 36606 33326 36960
rect 34488 37258 34546 37612
rect 34488 36966 34500 37258
rect 34534 36966 34546 37258
rect 34488 36612 34546 36966
rect 35546 37258 35604 37612
rect 35546 36966 35558 37258
rect 35592 36966 35604 37258
rect 35546 36612 35604 36966
rect 36604 37258 36662 37612
rect 36604 36966 36616 37258
rect 36650 36966 36662 37258
rect 36604 36612 36662 36966
rect 37662 37258 37720 37612
rect 37662 36966 37674 37258
rect 37708 36966 37720 37258
rect 37662 36612 37720 36966
rect 38720 37258 38778 37612
rect 38720 36966 38732 37258
rect 38766 36966 38778 37258
rect 38720 36612 38778 36966
rect 39778 37258 39836 37612
rect 39778 36966 39790 37258
rect 39824 36966 39836 37258
rect 39778 36612 39836 36966
rect 40978 37258 41036 37612
rect 40978 36966 40990 37258
rect 41024 36966 41036 37258
rect 40978 36612 41036 36966
rect 42036 37258 42094 37612
rect 42036 36966 42048 37258
rect 42082 36966 42094 37258
rect 42036 36612 42094 36966
rect 43094 37258 43152 37612
rect 43094 36966 43106 37258
rect 43140 36966 43152 37258
rect 43094 36612 43152 36966
rect 44152 37258 44210 37612
rect 44152 36966 44164 37258
rect 44198 36966 44210 37258
rect 44152 36612 44210 36966
rect 45210 37258 45268 37612
rect 45210 36966 45222 37258
rect 45256 36966 45268 37258
rect 45210 36612 45268 36966
rect 46268 37258 46326 37612
rect 46268 36966 46280 37258
rect 46314 36966 46326 37258
rect 46268 36612 46326 36966
rect 47566 37280 47624 37634
rect 47566 36988 47578 37280
rect 47612 36988 47624 37280
rect 47566 36634 47624 36988
rect 48624 37280 48682 37634
rect 48624 36988 48636 37280
rect 48670 36988 48682 37280
rect 48624 36634 48682 36988
rect 49682 37280 49740 37634
rect 49682 36988 49694 37280
rect 49728 36988 49740 37280
rect 49682 36634 49740 36988
rect 50740 37280 50798 37634
rect 50740 36988 50752 37280
rect 50786 36988 50798 37280
rect 50740 36634 50798 36988
rect 51798 37280 51856 37634
rect 51798 36988 51810 37280
rect 51844 36988 51856 37280
rect 51798 36634 51856 36988
rect 52856 37280 52914 37634
rect 52856 36988 52868 37280
rect 52902 36988 52914 37280
rect 52856 36634 52914 36988
rect 54080 37294 54138 37648
rect 54080 37002 54092 37294
rect 54126 37002 54138 37294
rect 54080 36648 54138 37002
rect 55138 37294 55196 37648
rect 55138 37002 55150 37294
rect 55184 37002 55196 37294
rect 55138 36648 55196 37002
rect 56196 37294 56254 37648
rect 56196 37002 56208 37294
rect 56242 37002 56254 37294
rect 56196 36648 56254 37002
rect 57254 37294 57312 37648
rect 57254 37002 57266 37294
rect 57300 37002 57312 37294
rect 57254 36648 57312 37002
rect 58312 37294 58370 37648
rect 58312 37002 58324 37294
rect 58358 37002 58370 37294
rect 58312 36648 58370 37002
rect 59370 37294 59428 37648
rect 59370 37002 59382 37294
rect 59416 37002 59428 37294
rect 59370 36648 59428 37002
rect 1946 36142 2004 36496
rect 1946 35850 1958 36142
rect 1992 35850 2004 36142
rect 1946 35496 2004 35850
rect 3004 36142 3062 36496
rect 3004 35850 3016 36142
rect 3050 35850 3062 36142
rect 3004 35496 3062 35850
rect 4062 36142 4120 36496
rect 4062 35850 4074 36142
rect 4108 35850 4120 36142
rect 4062 35496 4120 35850
rect 5120 36142 5178 36496
rect 5120 35850 5132 36142
rect 5166 35850 5178 36142
rect 5120 35496 5178 35850
rect 6178 36142 6236 36496
rect 6178 35850 6190 36142
rect 6224 35850 6236 36142
rect 6178 35496 6236 35850
rect 7236 36142 7294 36496
rect 7236 35850 7248 36142
rect 7282 35850 7294 36142
rect 8460 36150 8518 36504
rect 7236 35496 7294 35850
rect 1946 35048 2004 35402
rect 1946 34756 1958 35048
rect 1992 34756 2004 35048
rect 1946 34402 2004 34756
rect 3004 35048 3062 35402
rect 3004 34756 3016 35048
rect 3050 34756 3062 35048
rect 3004 34402 3062 34756
rect 4062 35048 4120 35402
rect 4062 34756 4074 35048
rect 4108 34756 4120 35048
rect 4062 34402 4120 34756
rect 5120 35048 5178 35402
rect 5120 34756 5132 35048
rect 5166 34756 5178 35048
rect 5120 34402 5178 34756
rect 6178 35048 6236 35402
rect 6178 34756 6190 35048
rect 6224 34756 6236 35048
rect 6178 34402 6236 34756
rect 7236 35048 7294 35402
rect 7236 34756 7248 35048
rect 7282 34756 7294 35048
rect 7236 34402 7294 34756
rect 8460 35858 8472 36150
rect 8506 35858 8518 36150
rect 8460 35504 8518 35858
rect 9518 36150 9576 36504
rect 9518 35858 9530 36150
rect 9564 35858 9576 36150
rect 9518 35504 9576 35858
rect 10576 36150 10634 36504
rect 10576 35858 10588 36150
rect 10622 35858 10634 36150
rect 10576 35504 10634 35858
rect 11634 36150 11692 36504
rect 11634 35858 11646 36150
rect 11680 35858 11692 36150
rect 11634 35504 11692 35858
rect 12692 36150 12750 36504
rect 12692 35858 12704 36150
rect 12738 35858 12750 36150
rect 12692 35504 12750 35858
rect 13750 36150 13808 36504
rect 13750 35858 13762 36150
rect 13796 35858 13808 36150
rect 14966 36158 15024 36512
rect 13750 35504 13808 35858
rect 1946 33954 2004 34308
rect 1946 33662 1958 33954
rect 1992 33662 2004 33954
rect 1946 33308 2004 33662
rect 3004 33954 3062 34308
rect 3004 33662 3016 33954
rect 3050 33662 3062 33954
rect 3004 33308 3062 33662
rect 4062 33954 4120 34308
rect 4062 33662 4074 33954
rect 4108 33662 4120 33954
rect 4062 33308 4120 33662
rect 5120 33954 5178 34308
rect 5120 33662 5132 33954
rect 5166 33662 5178 33954
rect 5120 33308 5178 33662
rect 6178 33954 6236 34308
rect 6178 33662 6190 33954
rect 6224 33662 6236 33954
rect 6178 33308 6236 33662
rect 7236 33954 7294 34308
rect 8460 35056 8518 35410
rect 8460 34764 8472 35056
rect 8506 34764 8518 35056
rect 8460 34410 8518 34764
rect 9518 35056 9576 35410
rect 9518 34764 9530 35056
rect 9564 34764 9576 35056
rect 9518 34410 9576 34764
rect 10576 35056 10634 35410
rect 10576 34764 10588 35056
rect 10622 34764 10634 35056
rect 10576 34410 10634 34764
rect 11634 35056 11692 35410
rect 11634 34764 11646 35056
rect 11680 34764 11692 35056
rect 11634 34410 11692 34764
rect 12692 35056 12750 35410
rect 12692 34764 12704 35056
rect 12738 34764 12750 35056
rect 12692 34410 12750 34764
rect 13750 35056 13808 35410
rect 13750 34764 13762 35056
rect 13796 34764 13808 35056
rect 13750 34410 13808 34764
rect 14966 35866 14978 36158
rect 15012 35866 15024 36158
rect 14966 35512 15024 35866
rect 16024 36158 16082 36512
rect 16024 35866 16036 36158
rect 16070 35866 16082 36158
rect 16024 35512 16082 35866
rect 17082 36158 17140 36512
rect 17082 35866 17094 36158
rect 17128 35866 17140 36158
rect 17082 35512 17140 35866
rect 18140 36158 18198 36512
rect 18140 35866 18152 36158
rect 18186 35866 18198 36158
rect 18140 35512 18198 35866
rect 19198 36158 19256 36512
rect 19198 35866 19210 36158
rect 19244 35866 19256 36158
rect 19198 35512 19256 35866
rect 20256 36158 20314 36512
rect 20256 35866 20268 36158
rect 20302 35866 20314 36158
rect 20256 35512 20314 35866
rect 21456 36142 21514 36496
rect 7236 33662 7248 33954
rect 7282 33662 7294 33954
rect 7236 33308 7294 33662
rect 8460 33962 8518 34316
rect 8460 33670 8472 33962
rect 8506 33670 8518 33962
rect 8460 33316 8518 33670
rect 9518 33962 9576 34316
rect 9518 33670 9530 33962
rect 9564 33670 9576 33962
rect 9518 33316 9576 33670
rect 10576 33962 10634 34316
rect 10576 33670 10588 33962
rect 10622 33670 10634 33962
rect 10576 33316 10634 33670
rect 11634 33962 11692 34316
rect 11634 33670 11646 33962
rect 11680 33670 11692 33962
rect 11634 33316 11692 33670
rect 12692 33962 12750 34316
rect 12692 33670 12704 33962
rect 12738 33670 12750 33962
rect 12692 33316 12750 33670
rect 13750 33962 13808 34316
rect 14966 35064 15024 35418
rect 14966 34772 14978 35064
rect 15012 34772 15024 35064
rect 14966 34418 15024 34772
rect 16024 35064 16082 35418
rect 16024 34772 16036 35064
rect 16070 34772 16082 35064
rect 16024 34418 16082 34772
rect 17082 35064 17140 35418
rect 17082 34772 17094 35064
rect 17128 34772 17140 35064
rect 17082 34418 17140 34772
rect 18140 35064 18198 35418
rect 18140 34772 18152 35064
rect 18186 34772 18198 35064
rect 18140 34418 18198 34772
rect 19198 35064 19256 35418
rect 19198 34772 19210 35064
rect 19244 34772 19256 35064
rect 19198 34418 19256 34772
rect 20256 35064 20314 35418
rect 20256 34772 20268 35064
rect 20302 34772 20314 35064
rect 20256 34418 20314 34772
rect 21456 35850 21468 36142
rect 21502 35850 21514 36142
rect 21456 35496 21514 35850
rect 22514 36142 22572 36496
rect 22514 35850 22526 36142
rect 22560 35850 22572 36142
rect 22514 35496 22572 35850
rect 23572 36142 23630 36496
rect 23572 35850 23584 36142
rect 23618 35850 23630 36142
rect 23572 35496 23630 35850
rect 24630 36142 24688 36496
rect 24630 35850 24642 36142
rect 24676 35850 24688 36142
rect 24630 35496 24688 35850
rect 25688 36142 25746 36496
rect 25688 35850 25700 36142
rect 25734 35850 25746 36142
rect 25688 35496 25746 35850
rect 26746 36142 26804 36496
rect 26746 35850 26758 36142
rect 26792 35850 26804 36142
rect 27978 36158 28036 36512
rect 26746 35496 26804 35850
rect 13750 33670 13762 33962
rect 13796 33670 13808 33962
rect 13750 33316 13808 33670
rect 14966 33970 15024 34324
rect 14966 33678 14978 33970
rect 15012 33678 15024 33970
rect 14966 33324 15024 33678
rect 16024 33970 16082 34324
rect 16024 33678 16036 33970
rect 16070 33678 16082 33970
rect 16024 33324 16082 33678
rect 17082 33970 17140 34324
rect 17082 33678 17094 33970
rect 17128 33678 17140 33970
rect 17082 33324 17140 33678
rect 18140 33970 18198 34324
rect 18140 33678 18152 33970
rect 18186 33678 18198 33970
rect 18140 33324 18198 33678
rect 19198 33970 19256 34324
rect 19198 33678 19210 33970
rect 19244 33678 19256 33970
rect 19198 33324 19256 33678
rect 20256 33970 20314 34324
rect 21456 35048 21514 35402
rect 21456 34756 21468 35048
rect 21502 34756 21514 35048
rect 21456 34402 21514 34756
rect 22514 35048 22572 35402
rect 22514 34756 22526 35048
rect 22560 34756 22572 35048
rect 22514 34402 22572 34756
rect 23572 35048 23630 35402
rect 23572 34756 23584 35048
rect 23618 34756 23630 35048
rect 23572 34402 23630 34756
rect 24630 35048 24688 35402
rect 24630 34756 24642 35048
rect 24676 34756 24688 35048
rect 24630 34402 24688 34756
rect 25688 35048 25746 35402
rect 25688 34756 25700 35048
rect 25734 34756 25746 35048
rect 25688 34402 25746 34756
rect 26746 35048 26804 35402
rect 26746 34756 26758 35048
rect 26792 34756 26804 35048
rect 26746 34402 26804 34756
rect 27978 35866 27990 36158
rect 28024 35866 28036 36158
rect 27978 35512 28036 35866
rect 29036 36158 29094 36512
rect 29036 35866 29048 36158
rect 29082 35866 29094 36158
rect 29036 35512 29094 35866
rect 30094 36158 30152 36512
rect 30094 35866 30106 36158
rect 30140 35866 30152 36158
rect 30094 35512 30152 35866
rect 31152 36158 31210 36512
rect 31152 35866 31164 36158
rect 31198 35866 31210 36158
rect 31152 35512 31210 35866
rect 32210 36158 32268 36512
rect 32210 35866 32222 36158
rect 32256 35866 32268 36158
rect 32210 35512 32268 35866
rect 33268 36158 33326 36512
rect 33268 35866 33280 36158
rect 33314 35866 33326 36158
rect 34488 36164 34546 36518
rect 33268 35512 33326 35866
rect 20256 33678 20268 33970
rect 20302 33678 20314 33970
rect 20256 33324 20314 33678
rect 21456 33954 21514 34308
rect 21456 33662 21468 33954
rect 21502 33662 21514 33954
rect 21456 33308 21514 33662
rect 22514 33954 22572 34308
rect 22514 33662 22526 33954
rect 22560 33662 22572 33954
rect 22514 33308 22572 33662
rect 23572 33954 23630 34308
rect 23572 33662 23584 33954
rect 23618 33662 23630 33954
rect 23572 33308 23630 33662
rect 24630 33954 24688 34308
rect 24630 33662 24642 33954
rect 24676 33662 24688 33954
rect 24630 33308 24688 33662
rect 25688 33954 25746 34308
rect 25688 33662 25700 33954
rect 25734 33662 25746 33954
rect 25688 33308 25746 33662
rect 26746 33954 26804 34308
rect 27978 35064 28036 35418
rect 27978 34772 27990 35064
rect 28024 34772 28036 35064
rect 27978 34418 28036 34772
rect 29036 35064 29094 35418
rect 29036 34772 29048 35064
rect 29082 34772 29094 35064
rect 29036 34418 29094 34772
rect 30094 35064 30152 35418
rect 30094 34772 30106 35064
rect 30140 34772 30152 35064
rect 30094 34418 30152 34772
rect 31152 35064 31210 35418
rect 31152 34772 31164 35064
rect 31198 34772 31210 35064
rect 31152 34418 31210 34772
rect 32210 35064 32268 35418
rect 32210 34772 32222 35064
rect 32256 34772 32268 35064
rect 32210 34418 32268 34772
rect 33268 35064 33326 35418
rect 33268 34772 33280 35064
rect 33314 34772 33326 35064
rect 33268 34418 33326 34772
rect 34488 35872 34500 36164
rect 34534 35872 34546 36164
rect 34488 35518 34546 35872
rect 35546 36164 35604 36518
rect 35546 35872 35558 36164
rect 35592 35872 35604 36164
rect 35546 35518 35604 35872
rect 36604 36164 36662 36518
rect 36604 35872 36616 36164
rect 36650 35872 36662 36164
rect 36604 35518 36662 35872
rect 37662 36164 37720 36518
rect 37662 35872 37674 36164
rect 37708 35872 37720 36164
rect 37662 35518 37720 35872
rect 38720 36164 38778 36518
rect 38720 35872 38732 36164
rect 38766 35872 38778 36164
rect 38720 35518 38778 35872
rect 39778 36164 39836 36518
rect 39778 35872 39790 36164
rect 39824 35872 39836 36164
rect 40978 36164 41036 36518
rect 39778 35518 39836 35872
rect 26746 33662 26758 33954
rect 26792 33662 26804 33954
rect 26746 33308 26804 33662
rect 27978 33970 28036 34324
rect 27978 33678 27990 33970
rect 28024 33678 28036 33970
rect 27978 33324 28036 33678
rect 29036 33970 29094 34324
rect 29036 33678 29048 33970
rect 29082 33678 29094 33970
rect 29036 33324 29094 33678
rect 30094 33970 30152 34324
rect 30094 33678 30106 33970
rect 30140 33678 30152 33970
rect 30094 33324 30152 33678
rect 31152 33970 31210 34324
rect 31152 33678 31164 33970
rect 31198 33678 31210 33970
rect 31152 33324 31210 33678
rect 32210 33970 32268 34324
rect 32210 33678 32222 33970
rect 32256 33678 32268 33970
rect 32210 33324 32268 33678
rect 33268 33970 33326 34324
rect 34488 35070 34546 35424
rect 34488 34778 34500 35070
rect 34534 34778 34546 35070
rect 34488 34424 34546 34778
rect 35546 35070 35604 35424
rect 35546 34778 35558 35070
rect 35592 34778 35604 35070
rect 35546 34424 35604 34778
rect 36604 35070 36662 35424
rect 36604 34778 36616 35070
rect 36650 34778 36662 35070
rect 36604 34424 36662 34778
rect 37662 35070 37720 35424
rect 37662 34778 37674 35070
rect 37708 34778 37720 35070
rect 37662 34424 37720 34778
rect 38720 35070 38778 35424
rect 38720 34778 38732 35070
rect 38766 34778 38778 35070
rect 38720 34424 38778 34778
rect 39778 35070 39836 35424
rect 39778 34778 39790 35070
rect 39824 34778 39836 35070
rect 39778 34424 39836 34778
rect 40978 35872 40990 36164
rect 41024 35872 41036 36164
rect 40978 35518 41036 35872
rect 42036 36164 42094 36518
rect 42036 35872 42048 36164
rect 42082 35872 42094 36164
rect 42036 35518 42094 35872
rect 43094 36164 43152 36518
rect 43094 35872 43106 36164
rect 43140 35872 43152 36164
rect 43094 35518 43152 35872
rect 44152 36164 44210 36518
rect 44152 35872 44164 36164
rect 44198 35872 44210 36164
rect 44152 35518 44210 35872
rect 45210 36164 45268 36518
rect 45210 35872 45222 36164
rect 45256 35872 45268 36164
rect 45210 35518 45268 35872
rect 46268 36164 46326 36518
rect 46268 35872 46280 36164
rect 46314 35872 46326 36164
rect 47566 36186 47624 36540
rect 46268 35518 46326 35872
rect 33268 33678 33280 33970
rect 33314 33678 33326 33970
rect 33268 33324 33326 33678
rect 34488 33976 34546 34330
rect 34488 33684 34500 33976
rect 34534 33684 34546 33976
rect 34488 33330 34546 33684
rect 35546 33976 35604 34330
rect 35546 33684 35558 33976
rect 35592 33684 35604 33976
rect 35546 33330 35604 33684
rect 36604 33976 36662 34330
rect 36604 33684 36616 33976
rect 36650 33684 36662 33976
rect 36604 33330 36662 33684
rect 37662 33976 37720 34330
rect 37662 33684 37674 33976
rect 37708 33684 37720 33976
rect 37662 33330 37720 33684
rect 38720 33976 38778 34330
rect 38720 33684 38732 33976
rect 38766 33684 38778 33976
rect 38720 33330 38778 33684
rect 39778 33976 39836 34330
rect 40978 35070 41036 35424
rect 40978 34778 40990 35070
rect 41024 34778 41036 35070
rect 40978 34424 41036 34778
rect 42036 35070 42094 35424
rect 42036 34778 42048 35070
rect 42082 34778 42094 35070
rect 42036 34424 42094 34778
rect 43094 35070 43152 35424
rect 43094 34778 43106 35070
rect 43140 34778 43152 35070
rect 43094 34424 43152 34778
rect 44152 35070 44210 35424
rect 44152 34778 44164 35070
rect 44198 34778 44210 35070
rect 44152 34424 44210 34778
rect 45210 35070 45268 35424
rect 45210 34778 45222 35070
rect 45256 34778 45268 35070
rect 45210 34424 45268 34778
rect 46268 35070 46326 35424
rect 46268 34778 46280 35070
rect 46314 34778 46326 35070
rect 46268 34424 46326 34778
rect 47566 35894 47578 36186
rect 47612 35894 47624 36186
rect 47566 35540 47624 35894
rect 48624 36186 48682 36540
rect 48624 35894 48636 36186
rect 48670 35894 48682 36186
rect 48624 35540 48682 35894
rect 49682 36186 49740 36540
rect 49682 35894 49694 36186
rect 49728 35894 49740 36186
rect 49682 35540 49740 35894
rect 50740 36186 50798 36540
rect 50740 35894 50752 36186
rect 50786 35894 50798 36186
rect 50740 35540 50798 35894
rect 51798 36186 51856 36540
rect 51798 35894 51810 36186
rect 51844 35894 51856 36186
rect 51798 35540 51856 35894
rect 52856 36186 52914 36540
rect 52856 35894 52868 36186
rect 52902 35894 52914 36186
rect 54080 36200 54138 36554
rect 52856 35540 52914 35894
rect 39778 33684 39790 33976
rect 39824 33684 39836 33976
rect 39778 33330 39836 33684
rect 40978 33976 41036 34330
rect 40978 33684 40990 33976
rect 41024 33684 41036 33976
rect 40978 33330 41036 33684
rect 42036 33976 42094 34330
rect 42036 33684 42048 33976
rect 42082 33684 42094 33976
rect 42036 33330 42094 33684
rect 43094 33976 43152 34330
rect 43094 33684 43106 33976
rect 43140 33684 43152 33976
rect 43094 33330 43152 33684
rect 44152 33976 44210 34330
rect 44152 33684 44164 33976
rect 44198 33684 44210 33976
rect 44152 33330 44210 33684
rect 45210 33976 45268 34330
rect 45210 33684 45222 33976
rect 45256 33684 45268 33976
rect 45210 33330 45268 33684
rect 46268 33976 46326 34330
rect 47566 35092 47624 35446
rect 47566 34800 47578 35092
rect 47612 34800 47624 35092
rect 47566 34446 47624 34800
rect 48624 35092 48682 35446
rect 48624 34800 48636 35092
rect 48670 34800 48682 35092
rect 48624 34446 48682 34800
rect 49682 35092 49740 35446
rect 49682 34800 49694 35092
rect 49728 34800 49740 35092
rect 49682 34446 49740 34800
rect 50740 35092 50798 35446
rect 50740 34800 50752 35092
rect 50786 34800 50798 35092
rect 50740 34446 50798 34800
rect 51798 35092 51856 35446
rect 51798 34800 51810 35092
rect 51844 34800 51856 35092
rect 51798 34446 51856 34800
rect 52856 35092 52914 35446
rect 52856 34800 52868 35092
rect 52902 34800 52914 35092
rect 52856 34446 52914 34800
rect 54080 35908 54092 36200
rect 54126 35908 54138 36200
rect 54080 35554 54138 35908
rect 55138 36200 55196 36554
rect 55138 35908 55150 36200
rect 55184 35908 55196 36200
rect 55138 35554 55196 35908
rect 56196 36200 56254 36554
rect 56196 35908 56208 36200
rect 56242 35908 56254 36200
rect 56196 35554 56254 35908
rect 57254 36200 57312 36554
rect 57254 35908 57266 36200
rect 57300 35908 57312 36200
rect 57254 35554 57312 35908
rect 58312 36200 58370 36554
rect 58312 35908 58324 36200
rect 58358 35908 58370 36200
rect 58312 35554 58370 35908
rect 59370 36200 59428 36554
rect 59370 35908 59382 36200
rect 59416 35908 59428 36200
rect 59370 35554 59428 35908
rect 62496 43108 62554 43322
rect 62496 42936 62508 43108
rect 62542 42936 62554 43108
rect 62496 42722 62554 42936
rect 63154 43108 63212 43322
rect 63154 42936 63166 43108
rect 63200 42936 63212 43108
rect 63154 42722 63212 42936
rect 63812 43108 63870 43322
rect 63812 42936 63824 43108
rect 63858 42936 63870 43108
rect 63812 42722 63870 42936
rect 64470 43108 64528 43322
rect 64470 42936 64482 43108
rect 64516 42936 64528 43108
rect 64470 42722 64528 42936
rect 65128 43108 65186 43322
rect 65128 42936 65140 43108
rect 65174 42936 65186 43108
rect 65128 42722 65186 42936
rect 65786 43108 65844 43322
rect 65786 42936 65798 43108
rect 65832 42936 65844 43108
rect 65786 42722 65844 42936
rect 66290 43110 66348 43324
rect 66290 42938 66302 43110
rect 66336 42938 66348 43110
rect 66290 42724 66348 42938
rect 66948 43110 67006 43324
rect 66948 42938 66960 43110
rect 66994 42938 67006 43110
rect 66948 42724 67006 42938
rect 67606 43110 67664 43324
rect 67606 42938 67618 43110
rect 67652 42938 67664 43110
rect 67606 42724 67664 42938
rect 68264 43110 68322 43324
rect 68264 42938 68276 43110
rect 68310 42938 68322 43110
rect 68264 42724 68322 42938
rect 68922 43110 68980 43324
rect 68922 42938 68934 43110
rect 68968 42938 68980 43110
rect 68922 42724 68980 42938
rect 69580 43110 69638 43324
rect 69580 42938 69592 43110
rect 69626 42938 69638 43110
rect 69580 42724 69638 42938
rect 70098 43124 70156 43338
rect 70098 42952 70110 43124
rect 70144 42952 70156 43124
rect 70098 42738 70156 42952
rect 70756 43124 70814 43338
rect 70756 42952 70768 43124
rect 70802 42952 70814 43124
rect 70756 42738 70814 42952
rect 71414 43124 71472 43338
rect 71414 42952 71426 43124
rect 71460 42952 71472 43124
rect 71414 42738 71472 42952
rect 72072 43124 72130 43338
rect 72072 42952 72084 43124
rect 72118 42952 72130 43124
rect 72072 42738 72130 42952
rect 72730 43124 72788 43338
rect 72730 42952 72742 43124
rect 72776 42952 72788 43124
rect 72730 42738 72788 42952
rect 73388 43124 73446 43338
rect 73388 42952 73400 43124
rect 73434 42952 73446 43124
rect 73388 42738 73446 42952
rect 62496 42414 62554 42628
rect 62496 42242 62508 42414
rect 62542 42242 62554 42414
rect 62496 42028 62554 42242
rect 63154 42414 63212 42628
rect 63154 42242 63166 42414
rect 63200 42242 63212 42414
rect 63154 42028 63212 42242
rect 63812 42414 63870 42628
rect 63812 42242 63824 42414
rect 63858 42242 63870 42414
rect 63812 42028 63870 42242
rect 64470 42414 64528 42628
rect 64470 42242 64482 42414
rect 64516 42242 64528 42414
rect 64470 42028 64528 42242
rect 65128 42414 65186 42628
rect 65128 42242 65140 42414
rect 65174 42242 65186 42414
rect 65128 42028 65186 42242
rect 65786 42414 65844 42628
rect 65786 42242 65798 42414
rect 65832 42242 65844 42414
rect 65786 42028 65844 42242
rect 62496 41720 62554 41934
rect 62496 41548 62508 41720
rect 62542 41548 62554 41720
rect 62496 41334 62554 41548
rect 63154 41720 63212 41934
rect 63154 41548 63166 41720
rect 63200 41548 63212 41720
rect 63154 41334 63212 41548
rect 63812 41720 63870 41934
rect 63812 41548 63824 41720
rect 63858 41548 63870 41720
rect 63812 41334 63870 41548
rect 64470 41720 64528 41934
rect 64470 41548 64482 41720
rect 64516 41548 64528 41720
rect 64470 41334 64528 41548
rect 65128 41720 65186 41934
rect 65128 41548 65140 41720
rect 65174 41548 65186 41720
rect 65128 41334 65186 41548
rect 65786 41720 65844 41934
rect 65786 41548 65798 41720
rect 65832 41548 65844 41720
rect 65786 41334 65844 41548
rect 62496 41026 62554 41240
rect 62496 40854 62508 41026
rect 62542 40854 62554 41026
rect 62496 40640 62554 40854
rect 63154 41026 63212 41240
rect 63154 40854 63166 41026
rect 63200 40854 63212 41026
rect 63154 40640 63212 40854
rect 63812 41026 63870 41240
rect 63812 40854 63824 41026
rect 63858 40854 63870 41026
rect 63812 40640 63870 40854
rect 64470 41026 64528 41240
rect 64470 40854 64482 41026
rect 64516 40854 64528 41026
rect 64470 40640 64528 40854
rect 65128 41026 65186 41240
rect 65128 40854 65140 41026
rect 65174 40854 65186 41026
rect 65128 40640 65186 40854
rect 65786 41026 65844 41240
rect 65786 40854 65798 41026
rect 65832 40854 65844 41026
rect 65786 40640 65844 40854
rect 66290 42416 66348 42630
rect 66290 42244 66302 42416
rect 66336 42244 66348 42416
rect 66290 42030 66348 42244
rect 66948 42416 67006 42630
rect 66948 42244 66960 42416
rect 66994 42244 67006 42416
rect 66948 42030 67006 42244
rect 67606 42416 67664 42630
rect 67606 42244 67618 42416
rect 67652 42244 67664 42416
rect 67606 42030 67664 42244
rect 68264 42416 68322 42630
rect 68264 42244 68276 42416
rect 68310 42244 68322 42416
rect 68264 42030 68322 42244
rect 68922 42416 68980 42630
rect 68922 42244 68934 42416
rect 68968 42244 68980 42416
rect 68922 42030 68980 42244
rect 69580 42416 69638 42630
rect 69580 42244 69592 42416
rect 69626 42244 69638 42416
rect 69580 42030 69638 42244
rect 66290 41722 66348 41936
rect 66290 41550 66302 41722
rect 66336 41550 66348 41722
rect 66290 41336 66348 41550
rect 66948 41722 67006 41936
rect 66948 41550 66960 41722
rect 66994 41550 67006 41722
rect 66948 41336 67006 41550
rect 67606 41722 67664 41936
rect 67606 41550 67618 41722
rect 67652 41550 67664 41722
rect 67606 41336 67664 41550
rect 68264 41722 68322 41936
rect 68264 41550 68276 41722
rect 68310 41550 68322 41722
rect 68264 41336 68322 41550
rect 68922 41722 68980 41936
rect 68922 41550 68934 41722
rect 68968 41550 68980 41722
rect 68922 41336 68980 41550
rect 69580 41722 69638 41936
rect 69580 41550 69592 41722
rect 69626 41550 69638 41722
rect 69580 41336 69638 41550
rect 66290 41028 66348 41242
rect 66290 40856 66302 41028
rect 66336 40856 66348 41028
rect 66290 40642 66348 40856
rect 66948 41028 67006 41242
rect 66948 40856 66960 41028
rect 66994 40856 67006 41028
rect 66948 40642 67006 40856
rect 67606 41028 67664 41242
rect 67606 40856 67618 41028
rect 67652 40856 67664 41028
rect 67606 40642 67664 40856
rect 68264 41028 68322 41242
rect 68264 40856 68276 41028
rect 68310 40856 68322 41028
rect 68264 40642 68322 40856
rect 68922 41028 68980 41242
rect 68922 40856 68934 41028
rect 68968 40856 68980 41028
rect 68922 40642 68980 40856
rect 69580 41028 69638 41242
rect 69580 40856 69592 41028
rect 69626 40856 69638 41028
rect 69580 40642 69638 40856
rect 70098 42430 70156 42644
rect 70098 42258 70110 42430
rect 70144 42258 70156 42430
rect 70098 42044 70156 42258
rect 70756 42430 70814 42644
rect 70756 42258 70768 42430
rect 70802 42258 70814 42430
rect 70756 42044 70814 42258
rect 71414 42430 71472 42644
rect 71414 42258 71426 42430
rect 71460 42258 71472 42430
rect 71414 42044 71472 42258
rect 72072 42430 72130 42644
rect 72072 42258 72084 42430
rect 72118 42258 72130 42430
rect 72072 42044 72130 42258
rect 72730 42430 72788 42644
rect 72730 42258 72742 42430
rect 72776 42258 72788 42430
rect 72730 42044 72788 42258
rect 73388 42430 73446 42644
rect 73388 42258 73400 42430
rect 73434 42258 73446 42430
rect 73388 42044 73446 42258
rect 70098 41736 70156 41950
rect 70098 41564 70110 41736
rect 70144 41564 70156 41736
rect 70098 41350 70156 41564
rect 70756 41736 70814 41950
rect 70756 41564 70768 41736
rect 70802 41564 70814 41736
rect 70756 41350 70814 41564
rect 71414 41736 71472 41950
rect 71414 41564 71426 41736
rect 71460 41564 71472 41736
rect 71414 41350 71472 41564
rect 72072 41736 72130 41950
rect 72072 41564 72084 41736
rect 72118 41564 72130 41736
rect 72072 41350 72130 41564
rect 72730 41736 72788 41950
rect 72730 41564 72742 41736
rect 72776 41564 72788 41736
rect 72730 41350 72788 41564
rect 73388 41736 73446 41950
rect 73388 41564 73400 41736
rect 73434 41564 73446 41736
rect 73388 41350 73446 41564
rect 70098 41042 70156 41256
rect 70098 40870 70110 41042
rect 70144 40870 70156 41042
rect 70098 40656 70156 40870
rect 70756 41042 70814 41256
rect 70756 40870 70768 41042
rect 70802 40870 70814 41042
rect 70756 40656 70814 40870
rect 71414 41042 71472 41256
rect 71414 40870 71426 41042
rect 71460 40870 71472 41042
rect 71414 40656 71472 40870
rect 72072 41042 72130 41256
rect 72072 40870 72084 41042
rect 72118 40870 72130 41042
rect 72072 40656 72130 40870
rect 72730 41042 72788 41256
rect 72730 40870 72742 41042
rect 72776 40870 72788 41042
rect 72730 40656 72788 40870
rect 73388 41042 73446 41256
rect 73388 40870 73400 41042
rect 73434 40870 73446 41042
rect 73388 40656 73446 40870
rect 62496 40332 62554 40546
rect 62496 40160 62508 40332
rect 62542 40160 62554 40332
rect 62496 39946 62554 40160
rect 63154 40332 63212 40546
rect 63154 40160 63166 40332
rect 63200 40160 63212 40332
rect 63154 39946 63212 40160
rect 63812 40332 63870 40546
rect 63812 40160 63824 40332
rect 63858 40160 63870 40332
rect 63812 39946 63870 40160
rect 64470 40332 64528 40546
rect 64470 40160 64482 40332
rect 64516 40160 64528 40332
rect 64470 39946 64528 40160
rect 65128 40332 65186 40546
rect 65128 40160 65140 40332
rect 65174 40160 65186 40332
rect 65128 39946 65186 40160
rect 65786 40332 65844 40546
rect 65786 40160 65798 40332
rect 65832 40160 65844 40332
rect 65786 39946 65844 40160
rect 66290 40334 66348 40548
rect 66290 40162 66302 40334
rect 66336 40162 66348 40334
rect 66290 39948 66348 40162
rect 66948 40334 67006 40548
rect 66948 40162 66960 40334
rect 66994 40162 67006 40334
rect 66948 39948 67006 40162
rect 67606 40334 67664 40548
rect 67606 40162 67618 40334
rect 67652 40162 67664 40334
rect 67606 39948 67664 40162
rect 68264 40334 68322 40548
rect 68264 40162 68276 40334
rect 68310 40162 68322 40334
rect 68264 39948 68322 40162
rect 68922 40334 68980 40548
rect 68922 40162 68934 40334
rect 68968 40162 68980 40334
rect 68922 39948 68980 40162
rect 69580 40334 69638 40548
rect 69580 40162 69592 40334
rect 69626 40162 69638 40334
rect 69580 39948 69638 40162
rect 70098 40348 70156 40562
rect 70098 40176 70110 40348
rect 70144 40176 70156 40348
rect 70098 39962 70156 40176
rect 70756 40348 70814 40562
rect 70756 40176 70768 40348
rect 70802 40176 70814 40348
rect 70756 39962 70814 40176
rect 71414 40348 71472 40562
rect 71414 40176 71426 40348
rect 71460 40176 71472 40348
rect 71414 39962 71472 40176
rect 72072 40348 72130 40562
rect 72072 40176 72084 40348
rect 72118 40176 72130 40348
rect 72072 39962 72130 40176
rect 72730 40348 72788 40562
rect 72730 40176 72742 40348
rect 72776 40176 72788 40348
rect 72730 39962 72788 40176
rect 73388 40348 73446 40562
rect 73388 40176 73400 40348
rect 73434 40176 73446 40348
rect 73388 39962 73446 40176
rect 46268 33684 46280 33976
rect 46314 33684 46326 33976
rect 46268 33330 46326 33684
rect 47566 33998 47624 34352
rect 47566 33706 47578 33998
rect 47612 33706 47624 33998
rect 47566 33352 47624 33706
rect 48624 33998 48682 34352
rect 48624 33706 48636 33998
rect 48670 33706 48682 33998
rect 48624 33352 48682 33706
rect 49682 33998 49740 34352
rect 49682 33706 49694 33998
rect 49728 33706 49740 33998
rect 49682 33352 49740 33706
rect 50740 33998 50798 34352
rect 50740 33706 50752 33998
rect 50786 33706 50798 33998
rect 50740 33352 50798 33706
rect 51798 33998 51856 34352
rect 51798 33706 51810 33998
rect 51844 33706 51856 33998
rect 51798 33352 51856 33706
rect 52856 33998 52914 34352
rect 54080 35106 54138 35460
rect 54080 34814 54092 35106
rect 54126 34814 54138 35106
rect 54080 34460 54138 34814
rect 55138 35106 55196 35460
rect 55138 34814 55150 35106
rect 55184 34814 55196 35106
rect 55138 34460 55196 34814
rect 56196 35106 56254 35460
rect 56196 34814 56208 35106
rect 56242 34814 56254 35106
rect 56196 34460 56254 34814
rect 57254 35106 57312 35460
rect 57254 34814 57266 35106
rect 57300 34814 57312 35106
rect 57254 34460 57312 34814
rect 58312 35106 58370 35460
rect 58312 34814 58324 35106
rect 58358 34814 58370 35106
rect 58312 34460 58370 34814
rect 59370 35106 59428 35460
rect 59370 34814 59382 35106
rect 59416 34814 59428 35106
rect 59370 34460 59428 34814
rect 77158 39094 77216 39308
rect 77158 38922 77170 39094
rect 77204 38922 77216 39094
rect 77158 38708 77216 38922
rect 77816 39094 77874 39308
rect 77816 38922 77828 39094
rect 77862 38922 77874 39094
rect 77816 38708 77874 38922
rect 78474 39094 78532 39308
rect 78474 38922 78486 39094
rect 78520 38922 78532 39094
rect 78474 38708 78532 38922
rect 79132 39094 79190 39308
rect 79132 38922 79144 39094
rect 79178 38922 79190 39094
rect 79132 38708 79190 38922
rect 79790 39094 79848 39308
rect 79790 38922 79802 39094
rect 79836 38922 79848 39094
rect 80484 39088 80542 39302
rect 79790 38708 79848 38922
rect 77158 38400 77216 38614
rect 77158 38228 77170 38400
rect 77204 38228 77216 38400
rect 77158 38014 77216 38228
rect 77816 38400 77874 38614
rect 77816 38228 77828 38400
rect 77862 38228 77874 38400
rect 77816 38014 77874 38228
rect 78474 38400 78532 38614
rect 78474 38228 78486 38400
rect 78520 38228 78532 38400
rect 78474 38014 78532 38228
rect 79132 38400 79190 38614
rect 79132 38228 79144 38400
rect 79178 38228 79190 38400
rect 79132 38014 79190 38228
rect 79790 38400 79848 38614
rect 79790 38228 79802 38400
rect 79836 38228 79848 38400
rect 79790 38014 79848 38228
rect 77158 37706 77216 37920
rect 77158 37534 77170 37706
rect 77204 37534 77216 37706
rect 77158 37320 77216 37534
rect 77816 37706 77874 37920
rect 77816 37534 77828 37706
rect 77862 37534 77874 37706
rect 77816 37320 77874 37534
rect 78474 37706 78532 37920
rect 78474 37534 78486 37706
rect 78520 37534 78532 37706
rect 78474 37320 78532 37534
rect 79132 37706 79190 37920
rect 79132 37534 79144 37706
rect 79178 37534 79190 37706
rect 79132 37320 79190 37534
rect 79790 37706 79848 37920
rect 79790 37534 79802 37706
rect 79836 37534 79848 37706
rect 79790 37320 79848 37534
rect 77158 37012 77216 37226
rect 77158 36840 77170 37012
rect 77204 36840 77216 37012
rect 77158 36626 77216 36840
rect 77816 37012 77874 37226
rect 77816 36840 77828 37012
rect 77862 36840 77874 37012
rect 77816 36626 77874 36840
rect 78474 37012 78532 37226
rect 78474 36840 78486 37012
rect 78520 36840 78532 37012
rect 78474 36626 78532 36840
rect 79132 37012 79190 37226
rect 79132 36840 79144 37012
rect 79178 36840 79190 37012
rect 79132 36626 79190 36840
rect 79790 37012 79848 37226
rect 79790 36840 79802 37012
rect 79836 36840 79848 37012
rect 79790 36626 79848 36840
rect 77158 36318 77216 36532
rect 77158 36146 77170 36318
rect 77204 36146 77216 36318
rect 77158 35932 77216 36146
rect 77816 36318 77874 36532
rect 77816 36146 77828 36318
rect 77862 36146 77874 36318
rect 77816 35932 77874 36146
rect 78474 36318 78532 36532
rect 78474 36146 78486 36318
rect 78520 36146 78532 36318
rect 78474 35932 78532 36146
rect 79132 36318 79190 36532
rect 79132 36146 79144 36318
rect 79178 36146 79190 36318
rect 79132 35932 79190 36146
rect 79790 36318 79848 36532
rect 79790 36146 79802 36318
rect 79836 36146 79848 36318
rect 79790 35932 79848 36146
rect 77158 35624 77216 35838
rect 77158 35452 77170 35624
rect 77204 35452 77216 35624
rect 77158 35238 77216 35452
rect 77816 35624 77874 35838
rect 77816 35452 77828 35624
rect 77862 35452 77874 35624
rect 77816 35238 77874 35452
rect 78474 35624 78532 35838
rect 78474 35452 78486 35624
rect 78520 35452 78532 35624
rect 78474 35238 78532 35452
rect 79132 35624 79190 35838
rect 79132 35452 79144 35624
rect 79178 35452 79190 35624
rect 79132 35238 79190 35452
rect 79790 35624 79848 35838
rect 79790 35452 79802 35624
rect 79836 35452 79848 35624
rect 80484 38916 80496 39088
rect 80530 38916 80542 39088
rect 80484 38702 80542 38916
rect 81142 39088 81200 39302
rect 81142 38916 81154 39088
rect 81188 38916 81200 39088
rect 81142 38702 81200 38916
rect 81800 39088 81858 39302
rect 81800 38916 81812 39088
rect 81846 38916 81858 39088
rect 81800 38702 81858 38916
rect 82458 39088 82516 39302
rect 82458 38916 82470 39088
rect 82504 38916 82516 39088
rect 82458 38702 82516 38916
rect 83116 39088 83174 39302
rect 83116 38916 83128 39088
rect 83162 38916 83174 39088
rect 83794 39088 83852 39302
rect 83116 38702 83174 38916
rect 80484 38394 80542 38608
rect 80484 38222 80496 38394
rect 80530 38222 80542 38394
rect 80484 38008 80542 38222
rect 81142 38394 81200 38608
rect 81142 38222 81154 38394
rect 81188 38222 81200 38394
rect 81142 38008 81200 38222
rect 81800 38394 81858 38608
rect 81800 38222 81812 38394
rect 81846 38222 81858 38394
rect 81800 38008 81858 38222
rect 82458 38394 82516 38608
rect 82458 38222 82470 38394
rect 82504 38222 82516 38394
rect 82458 38008 82516 38222
rect 83116 38394 83174 38608
rect 83116 38222 83128 38394
rect 83162 38222 83174 38394
rect 83116 38008 83174 38222
rect 80484 37700 80542 37914
rect 80484 37528 80496 37700
rect 80530 37528 80542 37700
rect 80484 37314 80542 37528
rect 81142 37700 81200 37914
rect 81142 37528 81154 37700
rect 81188 37528 81200 37700
rect 81142 37314 81200 37528
rect 81800 37700 81858 37914
rect 81800 37528 81812 37700
rect 81846 37528 81858 37700
rect 81800 37314 81858 37528
rect 82458 37700 82516 37914
rect 82458 37528 82470 37700
rect 82504 37528 82516 37700
rect 82458 37314 82516 37528
rect 83116 37700 83174 37914
rect 83116 37528 83128 37700
rect 83162 37528 83174 37700
rect 83116 37314 83174 37528
rect 80484 37006 80542 37220
rect 80484 36834 80496 37006
rect 80530 36834 80542 37006
rect 80484 36620 80542 36834
rect 81142 37006 81200 37220
rect 81142 36834 81154 37006
rect 81188 36834 81200 37006
rect 81142 36620 81200 36834
rect 81800 37006 81858 37220
rect 81800 36834 81812 37006
rect 81846 36834 81858 37006
rect 81800 36620 81858 36834
rect 82458 37006 82516 37220
rect 82458 36834 82470 37006
rect 82504 36834 82516 37006
rect 82458 36620 82516 36834
rect 83116 37006 83174 37220
rect 83116 36834 83128 37006
rect 83162 36834 83174 37006
rect 83116 36620 83174 36834
rect 80484 36312 80542 36526
rect 80484 36140 80496 36312
rect 80530 36140 80542 36312
rect 80484 35926 80542 36140
rect 81142 36312 81200 36526
rect 81142 36140 81154 36312
rect 81188 36140 81200 36312
rect 81142 35926 81200 36140
rect 81800 36312 81858 36526
rect 81800 36140 81812 36312
rect 81846 36140 81858 36312
rect 81800 35926 81858 36140
rect 82458 36312 82516 36526
rect 82458 36140 82470 36312
rect 82504 36140 82516 36312
rect 82458 35926 82516 36140
rect 83116 36312 83174 36526
rect 83116 36140 83128 36312
rect 83162 36140 83174 36312
rect 83116 35926 83174 36140
rect 80484 35618 80542 35832
rect 79790 35238 79848 35452
rect 80484 35446 80496 35618
rect 80530 35446 80542 35618
rect 80484 35232 80542 35446
rect 81142 35618 81200 35832
rect 81142 35446 81154 35618
rect 81188 35446 81200 35618
rect 81142 35232 81200 35446
rect 81800 35618 81858 35832
rect 81800 35446 81812 35618
rect 81846 35446 81858 35618
rect 81800 35232 81858 35446
rect 82458 35618 82516 35832
rect 82458 35446 82470 35618
rect 82504 35446 82516 35618
rect 82458 35232 82516 35446
rect 83116 35618 83174 35832
rect 83116 35446 83128 35618
rect 83162 35446 83174 35618
rect 83794 38916 83806 39088
rect 83840 38916 83852 39088
rect 83794 38702 83852 38916
rect 84452 39088 84510 39302
rect 84452 38916 84464 39088
rect 84498 38916 84510 39088
rect 84452 38702 84510 38916
rect 85110 39088 85168 39302
rect 85110 38916 85122 39088
rect 85156 38916 85168 39088
rect 85110 38702 85168 38916
rect 85768 39088 85826 39302
rect 85768 38916 85780 39088
rect 85814 38916 85826 39088
rect 85768 38702 85826 38916
rect 86426 39088 86484 39302
rect 86426 38916 86438 39088
rect 86472 38916 86484 39088
rect 86426 38702 86484 38916
rect 83794 38394 83852 38608
rect 83794 38222 83806 38394
rect 83840 38222 83852 38394
rect 83794 38008 83852 38222
rect 84452 38394 84510 38608
rect 84452 38222 84464 38394
rect 84498 38222 84510 38394
rect 84452 38008 84510 38222
rect 85110 38394 85168 38608
rect 85110 38222 85122 38394
rect 85156 38222 85168 38394
rect 85110 38008 85168 38222
rect 85768 38394 85826 38608
rect 85768 38222 85780 38394
rect 85814 38222 85826 38394
rect 85768 38008 85826 38222
rect 86426 38394 86484 38608
rect 86426 38222 86438 38394
rect 86472 38222 86484 38394
rect 86426 38008 86484 38222
rect 83794 37700 83852 37914
rect 83794 37528 83806 37700
rect 83840 37528 83852 37700
rect 83794 37314 83852 37528
rect 84452 37700 84510 37914
rect 84452 37528 84464 37700
rect 84498 37528 84510 37700
rect 84452 37314 84510 37528
rect 85110 37700 85168 37914
rect 85110 37528 85122 37700
rect 85156 37528 85168 37700
rect 85110 37314 85168 37528
rect 85768 37700 85826 37914
rect 85768 37528 85780 37700
rect 85814 37528 85826 37700
rect 85768 37314 85826 37528
rect 86426 37700 86484 37914
rect 86426 37528 86438 37700
rect 86472 37528 86484 37700
rect 86426 37314 86484 37528
rect 83794 37006 83852 37220
rect 83794 36834 83806 37006
rect 83840 36834 83852 37006
rect 83794 36620 83852 36834
rect 84452 37006 84510 37220
rect 84452 36834 84464 37006
rect 84498 36834 84510 37006
rect 84452 36620 84510 36834
rect 85110 37006 85168 37220
rect 85110 36834 85122 37006
rect 85156 36834 85168 37006
rect 85110 36620 85168 36834
rect 85768 37006 85826 37220
rect 85768 36834 85780 37006
rect 85814 36834 85826 37006
rect 85768 36620 85826 36834
rect 86426 37006 86484 37220
rect 86426 36834 86438 37006
rect 86472 36834 86484 37006
rect 86426 36620 86484 36834
rect 83794 36312 83852 36526
rect 83794 36140 83806 36312
rect 83840 36140 83852 36312
rect 83794 35926 83852 36140
rect 84452 36312 84510 36526
rect 84452 36140 84464 36312
rect 84498 36140 84510 36312
rect 84452 35926 84510 36140
rect 85110 36312 85168 36526
rect 85110 36140 85122 36312
rect 85156 36140 85168 36312
rect 85110 35926 85168 36140
rect 85768 36312 85826 36526
rect 85768 36140 85780 36312
rect 85814 36140 85826 36312
rect 85768 35926 85826 36140
rect 86426 36312 86484 36526
rect 86426 36140 86438 36312
rect 86472 36140 86484 36312
rect 86426 35926 86484 36140
rect 83794 35618 83852 35832
rect 83116 35232 83174 35446
rect 83794 35446 83806 35618
rect 83840 35446 83852 35618
rect 83794 35232 83852 35446
rect 84452 35618 84510 35832
rect 84452 35446 84464 35618
rect 84498 35446 84510 35618
rect 84452 35232 84510 35446
rect 85110 35618 85168 35832
rect 85110 35446 85122 35618
rect 85156 35446 85168 35618
rect 85110 35232 85168 35446
rect 85768 35618 85826 35832
rect 85768 35446 85780 35618
rect 85814 35446 85826 35618
rect 85768 35232 85826 35446
rect 86426 35618 86484 35832
rect 86426 35446 86438 35618
rect 86472 35446 86484 35618
rect 86426 35232 86484 35446
rect 52856 33706 52868 33998
rect 52902 33706 52914 33998
rect 52856 33352 52914 33706
rect 54080 34012 54138 34366
rect 54080 33720 54092 34012
rect 54126 33720 54138 34012
rect 54080 33366 54138 33720
rect 55138 34012 55196 34366
rect 55138 33720 55150 34012
rect 55184 33720 55196 34012
rect 55138 33366 55196 33720
rect 56196 34012 56254 34366
rect 56196 33720 56208 34012
rect 56242 33720 56254 34012
rect 56196 33366 56254 33720
rect 57254 34012 57312 34366
rect 57254 33720 57266 34012
rect 57300 33720 57312 34012
rect 57254 33366 57312 33720
rect 58312 34012 58370 34366
rect 58312 33720 58324 34012
rect 58358 33720 58370 34012
rect 58312 33366 58370 33720
rect 59370 34012 59428 34366
rect 59370 33720 59382 34012
rect 59416 33720 59428 34012
rect 59370 33366 59428 33720
rect 1946 32860 2004 33214
rect 1946 32568 1958 32860
rect 1992 32568 2004 32860
rect 1946 32214 2004 32568
rect 3004 32860 3062 33214
rect 3004 32568 3016 32860
rect 3050 32568 3062 32860
rect 3004 32214 3062 32568
rect 4062 32860 4120 33214
rect 4062 32568 4074 32860
rect 4108 32568 4120 32860
rect 4062 32214 4120 32568
rect 5120 32860 5178 33214
rect 5120 32568 5132 32860
rect 5166 32568 5178 32860
rect 5120 32214 5178 32568
rect 6178 32860 6236 33214
rect 6178 32568 6190 32860
rect 6224 32568 6236 32860
rect 6178 32214 6236 32568
rect 7236 32860 7294 33214
rect 7236 32568 7248 32860
rect 7282 32568 7294 32860
rect 7236 32214 7294 32568
rect 8460 32868 8518 33222
rect 8460 32576 8472 32868
rect 8506 32576 8518 32868
rect 8460 32222 8518 32576
rect 9518 32868 9576 33222
rect 9518 32576 9530 32868
rect 9564 32576 9576 32868
rect 9518 32222 9576 32576
rect 10576 32868 10634 33222
rect 10576 32576 10588 32868
rect 10622 32576 10634 32868
rect 10576 32222 10634 32576
rect 11634 32868 11692 33222
rect 11634 32576 11646 32868
rect 11680 32576 11692 32868
rect 11634 32222 11692 32576
rect 12692 32868 12750 33222
rect 12692 32576 12704 32868
rect 12738 32576 12750 32868
rect 12692 32222 12750 32576
rect 13750 32868 13808 33222
rect 13750 32576 13762 32868
rect 13796 32576 13808 32868
rect 13750 32222 13808 32576
rect 14966 32876 15024 33230
rect 14966 32584 14978 32876
rect 15012 32584 15024 32876
rect 14966 32230 15024 32584
rect 16024 32876 16082 33230
rect 16024 32584 16036 32876
rect 16070 32584 16082 32876
rect 16024 32230 16082 32584
rect 17082 32876 17140 33230
rect 17082 32584 17094 32876
rect 17128 32584 17140 32876
rect 17082 32230 17140 32584
rect 18140 32876 18198 33230
rect 18140 32584 18152 32876
rect 18186 32584 18198 32876
rect 18140 32230 18198 32584
rect 19198 32876 19256 33230
rect 19198 32584 19210 32876
rect 19244 32584 19256 32876
rect 19198 32230 19256 32584
rect 20256 32876 20314 33230
rect 20256 32584 20268 32876
rect 20302 32584 20314 32876
rect 20256 32230 20314 32584
rect 21456 32860 21514 33214
rect 21456 32568 21468 32860
rect 21502 32568 21514 32860
rect 21456 32214 21514 32568
rect 22514 32860 22572 33214
rect 22514 32568 22526 32860
rect 22560 32568 22572 32860
rect 22514 32214 22572 32568
rect 23572 32860 23630 33214
rect 23572 32568 23584 32860
rect 23618 32568 23630 32860
rect 23572 32214 23630 32568
rect 24630 32860 24688 33214
rect 24630 32568 24642 32860
rect 24676 32568 24688 32860
rect 24630 32214 24688 32568
rect 25688 32860 25746 33214
rect 25688 32568 25700 32860
rect 25734 32568 25746 32860
rect 25688 32214 25746 32568
rect 26746 32860 26804 33214
rect 26746 32568 26758 32860
rect 26792 32568 26804 32860
rect 26746 32214 26804 32568
rect 27978 32876 28036 33230
rect 27978 32584 27990 32876
rect 28024 32584 28036 32876
rect 27978 32230 28036 32584
rect 29036 32876 29094 33230
rect 29036 32584 29048 32876
rect 29082 32584 29094 32876
rect 29036 32230 29094 32584
rect 30094 32876 30152 33230
rect 30094 32584 30106 32876
rect 30140 32584 30152 32876
rect 30094 32230 30152 32584
rect 31152 32876 31210 33230
rect 31152 32584 31164 32876
rect 31198 32584 31210 32876
rect 31152 32230 31210 32584
rect 32210 32876 32268 33230
rect 32210 32584 32222 32876
rect 32256 32584 32268 32876
rect 32210 32230 32268 32584
rect 33268 32876 33326 33230
rect 33268 32584 33280 32876
rect 33314 32584 33326 32876
rect 33268 32230 33326 32584
rect 34488 32882 34546 33236
rect 34488 32590 34500 32882
rect 34534 32590 34546 32882
rect 34488 32236 34546 32590
rect 35546 32882 35604 33236
rect 35546 32590 35558 32882
rect 35592 32590 35604 32882
rect 35546 32236 35604 32590
rect 36604 32882 36662 33236
rect 36604 32590 36616 32882
rect 36650 32590 36662 32882
rect 36604 32236 36662 32590
rect 37662 32882 37720 33236
rect 37662 32590 37674 32882
rect 37708 32590 37720 32882
rect 37662 32236 37720 32590
rect 38720 32882 38778 33236
rect 38720 32590 38732 32882
rect 38766 32590 38778 32882
rect 38720 32236 38778 32590
rect 39778 32882 39836 33236
rect 39778 32590 39790 32882
rect 39824 32590 39836 32882
rect 39778 32236 39836 32590
rect 40978 32882 41036 33236
rect 40978 32590 40990 32882
rect 41024 32590 41036 32882
rect 40978 32236 41036 32590
rect 42036 32882 42094 33236
rect 42036 32590 42048 32882
rect 42082 32590 42094 32882
rect 42036 32236 42094 32590
rect 43094 32882 43152 33236
rect 43094 32590 43106 32882
rect 43140 32590 43152 32882
rect 43094 32236 43152 32590
rect 44152 32882 44210 33236
rect 44152 32590 44164 32882
rect 44198 32590 44210 32882
rect 44152 32236 44210 32590
rect 45210 32882 45268 33236
rect 45210 32590 45222 32882
rect 45256 32590 45268 32882
rect 45210 32236 45268 32590
rect 46268 32882 46326 33236
rect 46268 32590 46280 32882
rect 46314 32590 46326 32882
rect 46268 32236 46326 32590
rect 47566 32904 47624 33258
rect 47566 32612 47578 32904
rect 47612 32612 47624 32904
rect 47566 32258 47624 32612
rect 48624 32904 48682 33258
rect 48624 32612 48636 32904
rect 48670 32612 48682 32904
rect 48624 32258 48682 32612
rect 49682 32904 49740 33258
rect 49682 32612 49694 32904
rect 49728 32612 49740 32904
rect 49682 32258 49740 32612
rect 50740 32904 50798 33258
rect 50740 32612 50752 32904
rect 50786 32612 50798 32904
rect 50740 32258 50798 32612
rect 51798 32904 51856 33258
rect 51798 32612 51810 32904
rect 51844 32612 51856 32904
rect 51798 32258 51856 32612
rect 52856 32904 52914 33258
rect 52856 32612 52868 32904
rect 52902 32612 52914 32904
rect 52856 32258 52914 32612
rect 54080 32918 54138 33272
rect 54080 32626 54092 32918
rect 54126 32626 54138 32918
rect 54080 32272 54138 32626
rect 55138 32918 55196 33272
rect 55138 32626 55150 32918
rect 55184 32626 55196 32918
rect 55138 32272 55196 32626
rect 56196 32918 56254 33272
rect 56196 32626 56208 32918
rect 56242 32626 56254 32918
rect 56196 32272 56254 32626
rect 57254 32918 57312 33272
rect 57254 32626 57266 32918
rect 57300 32626 57312 32918
rect 57254 32272 57312 32626
rect 58312 32918 58370 33272
rect 58312 32626 58324 32918
rect 58358 32626 58370 32918
rect 58312 32272 58370 32626
rect 59370 32918 59428 33272
rect 59370 32626 59382 32918
rect 59416 32626 59428 32918
rect 59370 32272 59428 32626
rect 1946 31402 2004 31756
rect 1946 31110 1958 31402
rect 1992 31110 2004 31402
rect 1946 30756 2004 31110
rect 3004 31402 3062 31756
rect 3004 31110 3016 31402
rect 3050 31110 3062 31402
rect 3004 30756 3062 31110
rect 4062 31402 4120 31756
rect 4062 31110 4074 31402
rect 4108 31110 4120 31402
rect 4062 30756 4120 31110
rect 5120 31402 5178 31756
rect 5120 31110 5132 31402
rect 5166 31110 5178 31402
rect 5120 30756 5178 31110
rect 6178 31402 6236 31756
rect 6178 31110 6190 31402
rect 6224 31110 6236 31402
rect 6178 30756 6236 31110
rect 7236 31402 7294 31756
rect 7236 31110 7248 31402
rect 7282 31110 7294 31402
rect 7236 30756 7294 31110
rect 8460 31410 8518 31764
rect 8460 31118 8472 31410
rect 8506 31118 8518 31410
rect 8460 30764 8518 31118
rect 9518 31410 9576 31764
rect 9518 31118 9530 31410
rect 9564 31118 9576 31410
rect 9518 30764 9576 31118
rect 10576 31410 10634 31764
rect 10576 31118 10588 31410
rect 10622 31118 10634 31410
rect 10576 30764 10634 31118
rect 11634 31410 11692 31764
rect 11634 31118 11646 31410
rect 11680 31118 11692 31410
rect 11634 30764 11692 31118
rect 12692 31410 12750 31764
rect 12692 31118 12704 31410
rect 12738 31118 12750 31410
rect 12692 30764 12750 31118
rect 13750 31410 13808 31764
rect 13750 31118 13762 31410
rect 13796 31118 13808 31410
rect 13750 30764 13808 31118
rect 14966 31418 15024 31772
rect 14966 31126 14978 31418
rect 15012 31126 15024 31418
rect 14966 30772 15024 31126
rect 16024 31418 16082 31772
rect 16024 31126 16036 31418
rect 16070 31126 16082 31418
rect 16024 30772 16082 31126
rect 17082 31418 17140 31772
rect 17082 31126 17094 31418
rect 17128 31126 17140 31418
rect 17082 30772 17140 31126
rect 18140 31418 18198 31772
rect 18140 31126 18152 31418
rect 18186 31126 18198 31418
rect 18140 30772 18198 31126
rect 19198 31418 19256 31772
rect 19198 31126 19210 31418
rect 19244 31126 19256 31418
rect 19198 30772 19256 31126
rect 20256 31418 20314 31772
rect 20256 31126 20268 31418
rect 20302 31126 20314 31418
rect 20256 30772 20314 31126
rect 21456 31402 21514 31756
rect 21456 31110 21468 31402
rect 21502 31110 21514 31402
rect 21456 30756 21514 31110
rect 22514 31402 22572 31756
rect 22514 31110 22526 31402
rect 22560 31110 22572 31402
rect 22514 30756 22572 31110
rect 23572 31402 23630 31756
rect 23572 31110 23584 31402
rect 23618 31110 23630 31402
rect 23572 30756 23630 31110
rect 24630 31402 24688 31756
rect 24630 31110 24642 31402
rect 24676 31110 24688 31402
rect 24630 30756 24688 31110
rect 25688 31402 25746 31756
rect 25688 31110 25700 31402
rect 25734 31110 25746 31402
rect 25688 30756 25746 31110
rect 26746 31402 26804 31756
rect 26746 31110 26758 31402
rect 26792 31110 26804 31402
rect 26746 30756 26804 31110
rect 27978 31418 28036 31772
rect 27978 31126 27990 31418
rect 28024 31126 28036 31418
rect 27978 30772 28036 31126
rect 29036 31418 29094 31772
rect 29036 31126 29048 31418
rect 29082 31126 29094 31418
rect 29036 30772 29094 31126
rect 30094 31418 30152 31772
rect 30094 31126 30106 31418
rect 30140 31126 30152 31418
rect 30094 30772 30152 31126
rect 31152 31418 31210 31772
rect 31152 31126 31164 31418
rect 31198 31126 31210 31418
rect 31152 30772 31210 31126
rect 32210 31418 32268 31772
rect 32210 31126 32222 31418
rect 32256 31126 32268 31418
rect 32210 30772 32268 31126
rect 33268 31418 33326 31772
rect 33268 31126 33280 31418
rect 33314 31126 33326 31418
rect 33268 30772 33326 31126
rect 34488 31424 34546 31778
rect 34488 31132 34500 31424
rect 34534 31132 34546 31424
rect 34488 30778 34546 31132
rect 35546 31424 35604 31778
rect 35546 31132 35558 31424
rect 35592 31132 35604 31424
rect 35546 30778 35604 31132
rect 36604 31424 36662 31778
rect 36604 31132 36616 31424
rect 36650 31132 36662 31424
rect 36604 30778 36662 31132
rect 37662 31424 37720 31778
rect 37662 31132 37674 31424
rect 37708 31132 37720 31424
rect 37662 30778 37720 31132
rect 38720 31424 38778 31778
rect 38720 31132 38732 31424
rect 38766 31132 38778 31424
rect 38720 30778 38778 31132
rect 39778 31424 39836 31778
rect 39778 31132 39790 31424
rect 39824 31132 39836 31424
rect 39778 30778 39836 31132
rect 40978 31424 41036 31778
rect 40978 31132 40990 31424
rect 41024 31132 41036 31424
rect 40978 30778 41036 31132
rect 42036 31424 42094 31778
rect 42036 31132 42048 31424
rect 42082 31132 42094 31424
rect 42036 30778 42094 31132
rect 43094 31424 43152 31778
rect 43094 31132 43106 31424
rect 43140 31132 43152 31424
rect 43094 30778 43152 31132
rect 44152 31424 44210 31778
rect 44152 31132 44164 31424
rect 44198 31132 44210 31424
rect 44152 30778 44210 31132
rect 45210 31424 45268 31778
rect 45210 31132 45222 31424
rect 45256 31132 45268 31424
rect 45210 30778 45268 31132
rect 46268 31424 46326 31778
rect 46268 31132 46280 31424
rect 46314 31132 46326 31424
rect 46268 30778 46326 31132
rect 47566 31446 47624 31800
rect 47566 31154 47578 31446
rect 47612 31154 47624 31446
rect 47566 30800 47624 31154
rect 48624 31446 48682 31800
rect 48624 31154 48636 31446
rect 48670 31154 48682 31446
rect 48624 30800 48682 31154
rect 49682 31446 49740 31800
rect 49682 31154 49694 31446
rect 49728 31154 49740 31446
rect 49682 30800 49740 31154
rect 50740 31446 50798 31800
rect 50740 31154 50752 31446
rect 50786 31154 50798 31446
rect 50740 30800 50798 31154
rect 51798 31446 51856 31800
rect 51798 31154 51810 31446
rect 51844 31154 51856 31446
rect 51798 30800 51856 31154
rect 52856 31446 52914 31800
rect 52856 31154 52868 31446
rect 52902 31154 52914 31446
rect 52856 30800 52914 31154
rect 54080 31460 54138 31814
rect 54080 31168 54092 31460
rect 54126 31168 54138 31460
rect 54080 30814 54138 31168
rect 55138 31460 55196 31814
rect 55138 31168 55150 31460
rect 55184 31168 55196 31460
rect 55138 30814 55196 31168
rect 56196 31460 56254 31814
rect 56196 31168 56208 31460
rect 56242 31168 56254 31460
rect 56196 30814 56254 31168
rect 57254 31460 57312 31814
rect 57254 31168 57266 31460
rect 57300 31168 57312 31460
rect 57254 30814 57312 31168
rect 58312 31460 58370 31814
rect 58312 31168 58324 31460
rect 58358 31168 58370 31460
rect 58312 30814 58370 31168
rect 59370 31460 59428 31814
rect 59370 31168 59382 31460
rect 59416 31168 59428 31460
rect 59370 30814 59428 31168
rect 1946 30308 2004 30662
rect 1946 30016 1958 30308
rect 1992 30016 2004 30308
rect 1946 29662 2004 30016
rect 3004 30308 3062 30662
rect 3004 30016 3016 30308
rect 3050 30016 3062 30308
rect 3004 29662 3062 30016
rect 4062 30308 4120 30662
rect 4062 30016 4074 30308
rect 4108 30016 4120 30308
rect 4062 29662 4120 30016
rect 5120 30308 5178 30662
rect 5120 30016 5132 30308
rect 5166 30016 5178 30308
rect 5120 29662 5178 30016
rect 6178 30308 6236 30662
rect 6178 30016 6190 30308
rect 6224 30016 6236 30308
rect 6178 29662 6236 30016
rect 7236 30308 7294 30662
rect 7236 30016 7248 30308
rect 7282 30016 7294 30308
rect 8460 30316 8518 30670
rect 7236 29662 7294 30016
rect 1946 29214 2004 29568
rect 1946 28922 1958 29214
rect 1992 28922 2004 29214
rect 1946 28568 2004 28922
rect 3004 29214 3062 29568
rect 3004 28922 3016 29214
rect 3050 28922 3062 29214
rect 3004 28568 3062 28922
rect 4062 29214 4120 29568
rect 4062 28922 4074 29214
rect 4108 28922 4120 29214
rect 4062 28568 4120 28922
rect 5120 29214 5178 29568
rect 5120 28922 5132 29214
rect 5166 28922 5178 29214
rect 5120 28568 5178 28922
rect 6178 29214 6236 29568
rect 6178 28922 6190 29214
rect 6224 28922 6236 29214
rect 6178 28568 6236 28922
rect 7236 29214 7294 29568
rect 7236 28922 7248 29214
rect 7282 28922 7294 29214
rect 7236 28568 7294 28922
rect 8460 30024 8472 30316
rect 8506 30024 8518 30316
rect 8460 29670 8518 30024
rect 9518 30316 9576 30670
rect 9518 30024 9530 30316
rect 9564 30024 9576 30316
rect 9518 29670 9576 30024
rect 10576 30316 10634 30670
rect 10576 30024 10588 30316
rect 10622 30024 10634 30316
rect 10576 29670 10634 30024
rect 11634 30316 11692 30670
rect 11634 30024 11646 30316
rect 11680 30024 11692 30316
rect 11634 29670 11692 30024
rect 12692 30316 12750 30670
rect 12692 30024 12704 30316
rect 12738 30024 12750 30316
rect 12692 29670 12750 30024
rect 13750 30316 13808 30670
rect 13750 30024 13762 30316
rect 13796 30024 13808 30316
rect 14966 30324 15024 30678
rect 13750 29670 13808 30024
rect 1946 28120 2004 28474
rect 1946 27828 1958 28120
rect 1992 27828 2004 28120
rect 1946 27474 2004 27828
rect 3004 28120 3062 28474
rect 3004 27828 3016 28120
rect 3050 27828 3062 28120
rect 3004 27474 3062 27828
rect 4062 28120 4120 28474
rect 4062 27828 4074 28120
rect 4108 27828 4120 28120
rect 4062 27474 4120 27828
rect 5120 28120 5178 28474
rect 5120 27828 5132 28120
rect 5166 27828 5178 28120
rect 5120 27474 5178 27828
rect 6178 28120 6236 28474
rect 6178 27828 6190 28120
rect 6224 27828 6236 28120
rect 6178 27474 6236 27828
rect 7236 28120 7294 28474
rect 8460 29222 8518 29576
rect 8460 28930 8472 29222
rect 8506 28930 8518 29222
rect 8460 28576 8518 28930
rect 9518 29222 9576 29576
rect 9518 28930 9530 29222
rect 9564 28930 9576 29222
rect 9518 28576 9576 28930
rect 10576 29222 10634 29576
rect 10576 28930 10588 29222
rect 10622 28930 10634 29222
rect 10576 28576 10634 28930
rect 11634 29222 11692 29576
rect 11634 28930 11646 29222
rect 11680 28930 11692 29222
rect 11634 28576 11692 28930
rect 12692 29222 12750 29576
rect 12692 28930 12704 29222
rect 12738 28930 12750 29222
rect 12692 28576 12750 28930
rect 13750 29222 13808 29576
rect 13750 28930 13762 29222
rect 13796 28930 13808 29222
rect 13750 28576 13808 28930
rect 14966 30032 14978 30324
rect 15012 30032 15024 30324
rect 14966 29678 15024 30032
rect 16024 30324 16082 30678
rect 16024 30032 16036 30324
rect 16070 30032 16082 30324
rect 16024 29678 16082 30032
rect 17082 30324 17140 30678
rect 17082 30032 17094 30324
rect 17128 30032 17140 30324
rect 17082 29678 17140 30032
rect 18140 30324 18198 30678
rect 18140 30032 18152 30324
rect 18186 30032 18198 30324
rect 18140 29678 18198 30032
rect 19198 30324 19256 30678
rect 19198 30032 19210 30324
rect 19244 30032 19256 30324
rect 19198 29678 19256 30032
rect 20256 30324 20314 30678
rect 20256 30032 20268 30324
rect 20302 30032 20314 30324
rect 20256 29678 20314 30032
rect 21456 30308 21514 30662
rect 7236 27828 7248 28120
rect 7282 27828 7294 28120
rect 7236 27474 7294 27828
rect 8460 28128 8518 28482
rect 8460 27836 8472 28128
rect 8506 27836 8518 28128
rect 8460 27482 8518 27836
rect 9518 28128 9576 28482
rect 9518 27836 9530 28128
rect 9564 27836 9576 28128
rect 9518 27482 9576 27836
rect 10576 28128 10634 28482
rect 10576 27836 10588 28128
rect 10622 27836 10634 28128
rect 10576 27482 10634 27836
rect 11634 28128 11692 28482
rect 11634 27836 11646 28128
rect 11680 27836 11692 28128
rect 11634 27482 11692 27836
rect 12692 28128 12750 28482
rect 12692 27836 12704 28128
rect 12738 27836 12750 28128
rect 12692 27482 12750 27836
rect 13750 28128 13808 28482
rect 14966 29230 15024 29584
rect 14966 28938 14978 29230
rect 15012 28938 15024 29230
rect 14966 28584 15024 28938
rect 16024 29230 16082 29584
rect 16024 28938 16036 29230
rect 16070 28938 16082 29230
rect 16024 28584 16082 28938
rect 17082 29230 17140 29584
rect 17082 28938 17094 29230
rect 17128 28938 17140 29230
rect 17082 28584 17140 28938
rect 18140 29230 18198 29584
rect 18140 28938 18152 29230
rect 18186 28938 18198 29230
rect 18140 28584 18198 28938
rect 19198 29230 19256 29584
rect 19198 28938 19210 29230
rect 19244 28938 19256 29230
rect 19198 28584 19256 28938
rect 20256 29230 20314 29584
rect 20256 28938 20268 29230
rect 20302 28938 20314 29230
rect 20256 28584 20314 28938
rect 21456 30016 21468 30308
rect 21502 30016 21514 30308
rect 21456 29662 21514 30016
rect 22514 30308 22572 30662
rect 22514 30016 22526 30308
rect 22560 30016 22572 30308
rect 22514 29662 22572 30016
rect 23572 30308 23630 30662
rect 23572 30016 23584 30308
rect 23618 30016 23630 30308
rect 23572 29662 23630 30016
rect 24630 30308 24688 30662
rect 24630 30016 24642 30308
rect 24676 30016 24688 30308
rect 24630 29662 24688 30016
rect 25688 30308 25746 30662
rect 25688 30016 25700 30308
rect 25734 30016 25746 30308
rect 25688 29662 25746 30016
rect 26746 30308 26804 30662
rect 26746 30016 26758 30308
rect 26792 30016 26804 30308
rect 27978 30324 28036 30678
rect 26746 29662 26804 30016
rect 13750 27836 13762 28128
rect 13796 27836 13808 28128
rect 13750 27482 13808 27836
rect 14966 28136 15024 28490
rect 14966 27844 14978 28136
rect 15012 27844 15024 28136
rect 14966 27490 15024 27844
rect 16024 28136 16082 28490
rect 16024 27844 16036 28136
rect 16070 27844 16082 28136
rect 16024 27490 16082 27844
rect 17082 28136 17140 28490
rect 17082 27844 17094 28136
rect 17128 27844 17140 28136
rect 17082 27490 17140 27844
rect 18140 28136 18198 28490
rect 18140 27844 18152 28136
rect 18186 27844 18198 28136
rect 18140 27490 18198 27844
rect 19198 28136 19256 28490
rect 19198 27844 19210 28136
rect 19244 27844 19256 28136
rect 19198 27490 19256 27844
rect 20256 28136 20314 28490
rect 21456 29214 21514 29568
rect 21456 28922 21468 29214
rect 21502 28922 21514 29214
rect 21456 28568 21514 28922
rect 22514 29214 22572 29568
rect 22514 28922 22526 29214
rect 22560 28922 22572 29214
rect 22514 28568 22572 28922
rect 23572 29214 23630 29568
rect 23572 28922 23584 29214
rect 23618 28922 23630 29214
rect 23572 28568 23630 28922
rect 24630 29214 24688 29568
rect 24630 28922 24642 29214
rect 24676 28922 24688 29214
rect 24630 28568 24688 28922
rect 25688 29214 25746 29568
rect 25688 28922 25700 29214
rect 25734 28922 25746 29214
rect 25688 28568 25746 28922
rect 26746 29214 26804 29568
rect 26746 28922 26758 29214
rect 26792 28922 26804 29214
rect 26746 28568 26804 28922
rect 27978 30032 27990 30324
rect 28024 30032 28036 30324
rect 27978 29678 28036 30032
rect 29036 30324 29094 30678
rect 29036 30032 29048 30324
rect 29082 30032 29094 30324
rect 29036 29678 29094 30032
rect 30094 30324 30152 30678
rect 30094 30032 30106 30324
rect 30140 30032 30152 30324
rect 30094 29678 30152 30032
rect 31152 30324 31210 30678
rect 31152 30032 31164 30324
rect 31198 30032 31210 30324
rect 31152 29678 31210 30032
rect 32210 30324 32268 30678
rect 32210 30032 32222 30324
rect 32256 30032 32268 30324
rect 32210 29678 32268 30032
rect 33268 30324 33326 30678
rect 33268 30032 33280 30324
rect 33314 30032 33326 30324
rect 34488 30330 34546 30684
rect 33268 29678 33326 30032
rect 20256 27844 20268 28136
rect 20302 27844 20314 28136
rect 20256 27490 20314 27844
rect 21456 28120 21514 28474
rect 21456 27828 21468 28120
rect 21502 27828 21514 28120
rect 21456 27474 21514 27828
rect 22514 28120 22572 28474
rect 22514 27828 22526 28120
rect 22560 27828 22572 28120
rect 22514 27474 22572 27828
rect 23572 28120 23630 28474
rect 23572 27828 23584 28120
rect 23618 27828 23630 28120
rect 23572 27474 23630 27828
rect 24630 28120 24688 28474
rect 24630 27828 24642 28120
rect 24676 27828 24688 28120
rect 24630 27474 24688 27828
rect 25688 28120 25746 28474
rect 25688 27828 25700 28120
rect 25734 27828 25746 28120
rect 25688 27474 25746 27828
rect 26746 28120 26804 28474
rect 27978 29230 28036 29584
rect 27978 28938 27990 29230
rect 28024 28938 28036 29230
rect 27978 28584 28036 28938
rect 29036 29230 29094 29584
rect 29036 28938 29048 29230
rect 29082 28938 29094 29230
rect 29036 28584 29094 28938
rect 30094 29230 30152 29584
rect 30094 28938 30106 29230
rect 30140 28938 30152 29230
rect 30094 28584 30152 28938
rect 31152 29230 31210 29584
rect 31152 28938 31164 29230
rect 31198 28938 31210 29230
rect 31152 28584 31210 28938
rect 32210 29230 32268 29584
rect 32210 28938 32222 29230
rect 32256 28938 32268 29230
rect 32210 28584 32268 28938
rect 33268 29230 33326 29584
rect 33268 28938 33280 29230
rect 33314 28938 33326 29230
rect 33268 28584 33326 28938
rect 34488 30038 34500 30330
rect 34534 30038 34546 30330
rect 34488 29684 34546 30038
rect 35546 30330 35604 30684
rect 35546 30038 35558 30330
rect 35592 30038 35604 30330
rect 35546 29684 35604 30038
rect 36604 30330 36662 30684
rect 36604 30038 36616 30330
rect 36650 30038 36662 30330
rect 36604 29684 36662 30038
rect 37662 30330 37720 30684
rect 37662 30038 37674 30330
rect 37708 30038 37720 30330
rect 37662 29684 37720 30038
rect 38720 30330 38778 30684
rect 38720 30038 38732 30330
rect 38766 30038 38778 30330
rect 38720 29684 38778 30038
rect 39778 30330 39836 30684
rect 39778 30038 39790 30330
rect 39824 30038 39836 30330
rect 40978 30330 41036 30684
rect 39778 29684 39836 30038
rect 26746 27828 26758 28120
rect 26792 27828 26804 28120
rect 26746 27474 26804 27828
rect 27978 28136 28036 28490
rect 27978 27844 27990 28136
rect 28024 27844 28036 28136
rect 27978 27490 28036 27844
rect 29036 28136 29094 28490
rect 29036 27844 29048 28136
rect 29082 27844 29094 28136
rect 29036 27490 29094 27844
rect 30094 28136 30152 28490
rect 30094 27844 30106 28136
rect 30140 27844 30152 28136
rect 30094 27490 30152 27844
rect 31152 28136 31210 28490
rect 31152 27844 31164 28136
rect 31198 27844 31210 28136
rect 31152 27490 31210 27844
rect 32210 28136 32268 28490
rect 32210 27844 32222 28136
rect 32256 27844 32268 28136
rect 32210 27490 32268 27844
rect 33268 28136 33326 28490
rect 34488 29236 34546 29590
rect 34488 28944 34500 29236
rect 34534 28944 34546 29236
rect 34488 28590 34546 28944
rect 35546 29236 35604 29590
rect 35546 28944 35558 29236
rect 35592 28944 35604 29236
rect 35546 28590 35604 28944
rect 36604 29236 36662 29590
rect 36604 28944 36616 29236
rect 36650 28944 36662 29236
rect 36604 28590 36662 28944
rect 37662 29236 37720 29590
rect 37662 28944 37674 29236
rect 37708 28944 37720 29236
rect 37662 28590 37720 28944
rect 38720 29236 38778 29590
rect 38720 28944 38732 29236
rect 38766 28944 38778 29236
rect 38720 28590 38778 28944
rect 39778 29236 39836 29590
rect 39778 28944 39790 29236
rect 39824 28944 39836 29236
rect 39778 28590 39836 28944
rect 40978 30038 40990 30330
rect 41024 30038 41036 30330
rect 40978 29684 41036 30038
rect 42036 30330 42094 30684
rect 42036 30038 42048 30330
rect 42082 30038 42094 30330
rect 42036 29684 42094 30038
rect 43094 30330 43152 30684
rect 43094 30038 43106 30330
rect 43140 30038 43152 30330
rect 43094 29684 43152 30038
rect 44152 30330 44210 30684
rect 44152 30038 44164 30330
rect 44198 30038 44210 30330
rect 44152 29684 44210 30038
rect 45210 30330 45268 30684
rect 45210 30038 45222 30330
rect 45256 30038 45268 30330
rect 45210 29684 45268 30038
rect 46268 30330 46326 30684
rect 46268 30038 46280 30330
rect 46314 30038 46326 30330
rect 47566 30352 47624 30706
rect 46268 29684 46326 30038
rect 33268 27844 33280 28136
rect 33314 27844 33326 28136
rect 33268 27490 33326 27844
rect 34488 28142 34546 28496
rect 34488 27850 34500 28142
rect 34534 27850 34546 28142
rect 34488 27496 34546 27850
rect 35546 28142 35604 28496
rect 35546 27850 35558 28142
rect 35592 27850 35604 28142
rect 35546 27496 35604 27850
rect 36604 28142 36662 28496
rect 36604 27850 36616 28142
rect 36650 27850 36662 28142
rect 36604 27496 36662 27850
rect 37662 28142 37720 28496
rect 37662 27850 37674 28142
rect 37708 27850 37720 28142
rect 37662 27496 37720 27850
rect 38720 28142 38778 28496
rect 38720 27850 38732 28142
rect 38766 27850 38778 28142
rect 38720 27496 38778 27850
rect 39778 28142 39836 28496
rect 40978 29236 41036 29590
rect 40978 28944 40990 29236
rect 41024 28944 41036 29236
rect 40978 28590 41036 28944
rect 42036 29236 42094 29590
rect 42036 28944 42048 29236
rect 42082 28944 42094 29236
rect 42036 28590 42094 28944
rect 43094 29236 43152 29590
rect 43094 28944 43106 29236
rect 43140 28944 43152 29236
rect 43094 28590 43152 28944
rect 44152 29236 44210 29590
rect 44152 28944 44164 29236
rect 44198 28944 44210 29236
rect 44152 28590 44210 28944
rect 45210 29236 45268 29590
rect 45210 28944 45222 29236
rect 45256 28944 45268 29236
rect 45210 28590 45268 28944
rect 46268 29236 46326 29590
rect 46268 28944 46280 29236
rect 46314 28944 46326 29236
rect 46268 28590 46326 28944
rect 47566 30060 47578 30352
rect 47612 30060 47624 30352
rect 47566 29706 47624 30060
rect 48624 30352 48682 30706
rect 48624 30060 48636 30352
rect 48670 30060 48682 30352
rect 48624 29706 48682 30060
rect 49682 30352 49740 30706
rect 49682 30060 49694 30352
rect 49728 30060 49740 30352
rect 49682 29706 49740 30060
rect 50740 30352 50798 30706
rect 50740 30060 50752 30352
rect 50786 30060 50798 30352
rect 50740 29706 50798 30060
rect 51798 30352 51856 30706
rect 51798 30060 51810 30352
rect 51844 30060 51856 30352
rect 51798 29706 51856 30060
rect 52856 30352 52914 30706
rect 52856 30060 52868 30352
rect 52902 30060 52914 30352
rect 54080 30366 54138 30720
rect 52856 29706 52914 30060
rect 39778 27850 39790 28142
rect 39824 27850 39836 28142
rect 39778 27496 39836 27850
rect 40978 28142 41036 28496
rect 40978 27850 40990 28142
rect 41024 27850 41036 28142
rect 40978 27496 41036 27850
rect 42036 28142 42094 28496
rect 42036 27850 42048 28142
rect 42082 27850 42094 28142
rect 42036 27496 42094 27850
rect 43094 28142 43152 28496
rect 43094 27850 43106 28142
rect 43140 27850 43152 28142
rect 43094 27496 43152 27850
rect 44152 28142 44210 28496
rect 44152 27850 44164 28142
rect 44198 27850 44210 28142
rect 44152 27496 44210 27850
rect 45210 28142 45268 28496
rect 45210 27850 45222 28142
rect 45256 27850 45268 28142
rect 45210 27496 45268 27850
rect 46268 28142 46326 28496
rect 47566 29258 47624 29612
rect 47566 28966 47578 29258
rect 47612 28966 47624 29258
rect 47566 28612 47624 28966
rect 48624 29258 48682 29612
rect 48624 28966 48636 29258
rect 48670 28966 48682 29258
rect 48624 28612 48682 28966
rect 49682 29258 49740 29612
rect 49682 28966 49694 29258
rect 49728 28966 49740 29258
rect 49682 28612 49740 28966
rect 50740 29258 50798 29612
rect 50740 28966 50752 29258
rect 50786 28966 50798 29258
rect 50740 28612 50798 28966
rect 51798 29258 51856 29612
rect 51798 28966 51810 29258
rect 51844 28966 51856 29258
rect 51798 28612 51856 28966
rect 52856 29258 52914 29612
rect 52856 28966 52868 29258
rect 52902 28966 52914 29258
rect 52856 28612 52914 28966
rect 54080 30074 54092 30366
rect 54126 30074 54138 30366
rect 54080 29720 54138 30074
rect 55138 30366 55196 30720
rect 55138 30074 55150 30366
rect 55184 30074 55196 30366
rect 55138 29720 55196 30074
rect 56196 30366 56254 30720
rect 56196 30074 56208 30366
rect 56242 30074 56254 30366
rect 56196 29720 56254 30074
rect 57254 30366 57312 30720
rect 57254 30074 57266 30366
rect 57300 30074 57312 30366
rect 57254 29720 57312 30074
rect 58312 30366 58370 30720
rect 58312 30074 58324 30366
rect 58358 30074 58370 30366
rect 58312 29720 58370 30074
rect 59370 30366 59428 30720
rect 59370 30074 59382 30366
rect 59416 30074 59428 30366
rect 59370 29720 59428 30074
rect 46268 27850 46280 28142
rect 46314 27850 46326 28142
rect 46268 27496 46326 27850
rect 47566 28164 47624 28518
rect 47566 27872 47578 28164
rect 47612 27872 47624 28164
rect 47566 27518 47624 27872
rect 48624 28164 48682 28518
rect 48624 27872 48636 28164
rect 48670 27872 48682 28164
rect 48624 27518 48682 27872
rect 49682 28164 49740 28518
rect 49682 27872 49694 28164
rect 49728 27872 49740 28164
rect 49682 27518 49740 27872
rect 50740 28164 50798 28518
rect 50740 27872 50752 28164
rect 50786 27872 50798 28164
rect 50740 27518 50798 27872
rect 51798 28164 51856 28518
rect 51798 27872 51810 28164
rect 51844 27872 51856 28164
rect 51798 27518 51856 27872
rect 52856 28164 52914 28518
rect 54080 29272 54138 29626
rect 54080 28980 54092 29272
rect 54126 28980 54138 29272
rect 54080 28626 54138 28980
rect 55138 29272 55196 29626
rect 55138 28980 55150 29272
rect 55184 28980 55196 29272
rect 55138 28626 55196 28980
rect 56196 29272 56254 29626
rect 56196 28980 56208 29272
rect 56242 28980 56254 29272
rect 56196 28626 56254 28980
rect 57254 29272 57312 29626
rect 57254 28980 57266 29272
rect 57300 28980 57312 29272
rect 57254 28626 57312 28980
rect 58312 29272 58370 29626
rect 58312 28980 58324 29272
rect 58358 28980 58370 29272
rect 58312 28626 58370 28980
rect 59370 29272 59428 29626
rect 59370 28980 59382 29272
rect 59416 28980 59428 29272
rect 59370 28626 59428 28980
rect 52856 27872 52868 28164
rect 52902 27872 52914 28164
rect 52856 27518 52914 27872
rect 54080 28178 54138 28532
rect 54080 27886 54092 28178
rect 54126 27886 54138 28178
rect 54080 27532 54138 27886
rect 55138 28178 55196 28532
rect 55138 27886 55150 28178
rect 55184 27886 55196 28178
rect 55138 27532 55196 27886
rect 56196 28178 56254 28532
rect 56196 27886 56208 28178
rect 56242 27886 56254 28178
rect 56196 27532 56254 27886
rect 57254 28178 57312 28532
rect 57254 27886 57266 28178
rect 57300 27886 57312 28178
rect 57254 27532 57312 27886
rect 58312 28178 58370 28532
rect 58312 27886 58324 28178
rect 58358 27886 58370 28178
rect 58312 27532 58370 27886
rect 59370 28178 59428 28532
rect 59370 27886 59382 28178
rect 59416 27886 59428 28178
rect 59370 27532 59428 27886
rect 1946 27026 2004 27380
rect 1946 26734 1958 27026
rect 1992 26734 2004 27026
rect 1946 26380 2004 26734
rect 3004 27026 3062 27380
rect 3004 26734 3016 27026
rect 3050 26734 3062 27026
rect 3004 26380 3062 26734
rect 4062 27026 4120 27380
rect 4062 26734 4074 27026
rect 4108 26734 4120 27026
rect 4062 26380 4120 26734
rect 5120 27026 5178 27380
rect 5120 26734 5132 27026
rect 5166 26734 5178 27026
rect 5120 26380 5178 26734
rect 6178 27026 6236 27380
rect 6178 26734 6190 27026
rect 6224 26734 6236 27026
rect 6178 26380 6236 26734
rect 7236 27026 7294 27380
rect 7236 26734 7248 27026
rect 7282 26734 7294 27026
rect 7236 26380 7294 26734
rect 8460 27034 8518 27388
rect 8460 26742 8472 27034
rect 8506 26742 8518 27034
rect 8460 26388 8518 26742
rect 9518 27034 9576 27388
rect 9518 26742 9530 27034
rect 9564 26742 9576 27034
rect 9518 26388 9576 26742
rect 10576 27034 10634 27388
rect 10576 26742 10588 27034
rect 10622 26742 10634 27034
rect 10576 26388 10634 26742
rect 11634 27034 11692 27388
rect 11634 26742 11646 27034
rect 11680 26742 11692 27034
rect 11634 26388 11692 26742
rect 12692 27034 12750 27388
rect 12692 26742 12704 27034
rect 12738 26742 12750 27034
rect 12692 26388 12750 26742
rect 13750 27034 13808 27388
rect 13750 26742 13762 27034
rect 13796 26742 13808 27034
rect 13750 26388 13808 26742
rect 14966 27042 15024 27396
rect 14966 26750 14978 27042
rect 15012 26750 15024 27042
rect 14966 26396 15024 26750
rect 16024 27042 16082 27396
rect 16024 26750 16036 27042
rect 16070 26750 16082 27042
rect 16024 26396 16082 26750
rect 17082 27042 17140 27396
rect 17082 26750 17094 27042
rect 17128 26750 17140 27042
rect 17082 26396 17140 26750
rect 18140 27042 18198 27396
rect 18140 26750 18152 27042
rect 18186 26750 18198 27042
rect 18140 26396 18198 26750
rect 19198 27042 19256 27396
rect 19198 26750 19210 27042
rect 19244 26750 19256 27042
rect 19198 26396 19256 26750
rect 20256 27042 20314 27396
rect 20256 26750 20268 27042
rect 20302 26750 20314 27042
rect 20256 26396 20314 26750
rect 21456 27026 21514 27380
rect 21456 26734 21468 27026
rect 21502 26734 21514 27026
rect 21456 26380 21514 26734
rect 22514 27026 22572 27380
rect 22514 26734 22526 27026
rect 22560 26734 22572 27026
rect 22514 26380 22572 26734
rect 23572 27026 23630 27380
rect 23572 26734 23584 27026
rect 23618 26734 23630 27026
rect 23572 26380 23630 26734
rect 24630 27026 24688 27380
rect 24630 26734 24642 27026
rect 24676 26734 24688 27026
rect 24630 26380 24688 26734
rect 25688 27026 25746 27380
rect 25688 26734 25700 27026
rect 25734 26734 25746 27026
rect 25688 26380 25746 26734
rect 26746 27026 26804 27380
rect 26746 26734 26758 27026
rect 26792 26734 26804 27026
rect 26746 26380 26804 26734
rect 27978 27042 28036 27396
rect 27978 26750 27990 27042
rect 28024 26750 28036 27042
rect 27978 26396 28036 26750
rect 29036 27042 29094 27396
rect 29036 26750 29048 27042
rect 29082 26750 29094 27042
rect 29036 26396 29094 26750
rect 30094 27042 30152 27396
rect 30094 26750 30106 27042
rect 30140 26750 30152 27042
rect 30094 26396 30152 26750
rect 31152 27042 31210 27396
rect 31152 26750 31164 27042
rect 31198 26750 31210 27042
rect 31152 26396 31210 26750
rect 32210 27042 32268 27396
rect 32210 26750 32222 27042
rect 32256 26750 32268 27042
rect 32210 26396 32268 26750
rect 33268 27042 33326 27396
rect 33268 26750 33280 27042
rect 33314 26750 33326 27042
rect 33268 26396 33326 26750
rect 34488 27048 34546 27402
rect 34488 26756 34500 27048
rect 34534 26756 34546 27048
rect 34488 26402 34546 26756
rect 35546 27048 35604 27402
rect 35546 26756 35558 27048
rect 35592 26756 35604 27048
rect 35546 26402 35604 26756
rect 36604 27048 36662 27402
rect 36604 26756 36616 27048
rect 36650 26756 36662 27048
rect 36604 26402 36662 26756
rect 37662 27048 37720 27402
rect 37662 26756 37674 27048
rect 37708 26756 37720 27048
rect 37662 26402 37720 26756
rect 38720 27048 38778 27402
rect 38720 26756 38732 27048
rect 38766 26756 38778 27048
rect 38720 26402 38778 26756
rect 39778 27048 39836 27402
rect 39778 26756 39790 27048
rect 39824 26756 39836 27048
rect 39778 26402 39836 26756
rect 40978 27048 41036 27402
rect 40978 26756 40990 27048
rect 41024 26756 41036 27048
rect 40978 26402 41036 26756
rect 42036 27048 42094 27402
rect 42036 26756 42048 27048
rect 42082 26756 42094 27048
rect 42036 26402 42094 26756
rect 43094 27048 43152 27402
rect 43094 26756 43106 27048
rect 43140 26756 43152 27048
rect 43094 26402 43152 26756
rect 44152 27048 44210 27402
rect 44152 26756 44164 27048
rect 44198 26756 44210 27048
rect 44152 26402 44210 26756
rect 45210 27048 45268 27402
rect 45210 26756 45222 27048
rect 45256 26756 45268 27048
rect 45210 26402 45268 26756
rect 46268 27048 46326 27402
rect 46268 26756 46280 27048
rect 46314 26756 46326 27048
rect 46268 26402 46326 26756
rect 47566 27070 47624 27424
rect 47566 26778 47578 27070
rect 47612 26778 47624 27070
rect 47566 26424 47624 26778
rect 48624 27070 48682 27424
rect 48624 26778 48636 27070
rect 48670 26778 48682 27070
rect 48624 26424 48682 26778
rect 49682 27070 49740 27424
rect 49682 26778 49694 27070
rect 49728 26778 49740 27070
rect 49682 26424 49740 26778
rect 50740 27070 50798 27424
rect 50740 26778 50752 27070
rect 50786 26778 50798 27070
rect 50740 26424 50798 26778
rect 51798 27070 51856 27424
rect 51798 26778 51810 27070
rect 51844 26778 51856 27070
rect 51798 26424 51856 26778
rect 52856 27070 52914 27424
rect 52856 26778 52868 27070
rect 52902 26778 52914 27070
rect 52856 26424 52914 26778
rect 54080 27084 54138 27438
rect 54080 26792 54092 27084
rect 54126 26792 54138 27084
rect 54080 26438 54138 26792
rect 55138 27084 55196 27438
rect 55138 26792 55150 27084
rect 55184 26792 55196 27084
rect 55138 26438 55196 26792
rect 56196 27084 56254 27438
rect 56196 26792 56208 27084
rect 56242 26792 56254 27084
rect 56196 26438 56254 26792
rect 57254 27084 57312 27438
rect 57254 26792 57266 27084
rect 57300 26792 57312 27084
rect 57254 26438 57312 26792
rect 58312 27084 58370 27438
rect 58312 26792 58324 27084
rect 58358 26792 58370 27084
rect 58312 26438 58370 26792
rect 59370 27084 59428 27438
rect 59370 26792 59382 27084
rect 59416 26792 59428 27084
rect 59370 26438 59428 26792
rect 1946 25566 2004 25920
rect 1946 25274 1958 25566
rect 1992 25274 2004 25566
rect 1946 24920 2004 25274
rect 3004 25566 3062 25920
rect 3004 25274 3016 25566
rect 3050 25274 3062 25566
rect 3004 24920 3062 25274
rect 4062 25566 4120 25920
rect 4062 25274 4074 25566
rect 4108 25274 4120 25566
rect 4062 24920 4120 25274
rect 5120 25566 5178 25920
rect 5120 25274 5132 25566
rect 5166 25274 5178 25566
rect 5120 24920 5178 25274
rect 6178 25566 6236 25920
rect 6178 25274 6190 25566
rect 6224 25274 6236 25566
rect 6178 24920 6236 25274
rect 7236 25566 7294 25920
rect 7236 25274 7248 25566
rect 7282 25274 7294 25566
rect 7236 24920 7294 25274
rect 8460 25574 8518 25928
rect 8460 25282 8472 25574
rect 8506 25282 8518 25574
rect 8460 24928 8518 25282
rect 9518 25574 9576 25928
rect 9518 25282 9530 25574
rect 9564 25282 9576 25574
rect 9518 24928 9576 25282
rect 10576 25574 10634 25928
rect 10576 25282 10588 25574
rect 10622 25282 10634 25574
rect 10576 24928 10634 25282
rect 11634 25574 11692 25928
rect 11634 25282 11646 25574
rect 11680 25282 11692 25574
rect 11634 24928 11692 25282
rect 12692 25574 12750 25928
rect 12692 25282 12704 25574
rect 12738 25282 12750 25574
rect 12692 24928 12750 25282
rect 13750 25574 13808 25928
rect 13750 25282 13762 25574
rect 13796 25282 13808 25574
rect 13750 24928 13808 25282
rect 14966 25582 15024 25936
rect 14966 25290 14978 25582
rect 15012 25290 15024 25582
rect 14966 24936 15024 25290
rect 16024 25582 16082 25936
rect 16024 25290 16036 25582
rect 16070 25290 16082 25582
rect 16024 24936 16082 25290
rect 17082 25582 17140 25936
rect 17082 25290 17094 25582
rect 17128 25290 17140 25582
rect 17082 24936 17140 25290
rect 18140 25582 18198 25936
rect 18140 25290 18152 25582
rect 18186 25290 18198 25582
rect 18140 24936 18198 25290
rect 19198 25582 19256 25936
rect 19198 25290 19210 25582
rect 19244 25290 19256 25582
rect 19198 24936 19256 25290
rect 20256 25582 20314 25936
rect 20256 25290 20268 25582
rect 20302 25290 20314 25582
rect 20256 24936 20314 25290
rect 21456 25566 21514 25920
rect 21456 25274 21468 25566
rect 21502 25274 21514 25566
rect 21456 24920 21514 25274
rect 22514 25566 22572 25920
rect 22514 25274 22526 25566
rect 22560 25274 22572 25566
rect 22514 24920 22572 25274
rect 23572 25566 23630 25920
rect 23572 25274 23584 25566
rect 23618 25274 23630 25566
rect 23572 24920 23630 25274
rect 24630 25566 24688 25920
rect 24630 25274 24642 25566
rect 24676 25274 24688 25566
rect 24630 24920 24688 25274
rect 25688 25566 25746 25920
rect 25688 25274 25700 25566
rect 25734 25274 25746 25566
rect 25688 24920 25746 25274
rect 26746 25566 26804 25920
rect 26746 25274 26758 25566
rect 26792 25274 26804 25566
rect 26746 24920 26804 25274
rect 27978 25582 28036 25936
rect 27978 25290 27990 25582
rect 28024 25290 28036 25582
rect 27978 24936 28036 25290
rect 29036 25582 29094 25936
rect 29036 25290 29048 25582
rect 29082 25290 29094 25582
rect 29036 24936 29094 25290
rect 30094 25582 30152 25936
rect 30094 25290 30106 25582
rect 30140 25290 30152 25582
rect 30094 24936 30152 25290
rect 31152 25582 31210 25936
rect 31152 25290 31164 25582
rect 31198 25290 31210 25582
rect 31152 24936 31210 25290
rect 32210 25582 32268 25936
rect 32210 25290 32222 25582
rect 32256 25290 32268 25582
rect 32210 24936 32268 25290
rect 33268 25582 33326 25936
rect 33268 25290 33280 25582
rect 33314 25290 33326 25582
rect 33268 24936 33326 25290
rect 34488 25588 34546 25942
rect 34488 25296 34500 25588
rect 34534 25296 34546 25588
rect 34488 24942 34546 25296
rect 35546 25588 35604 25942
rect 35546 25296 35558 25588
rect 35592 25296 35604 25588
rect 35546 24942 35604 25296
rect 36604 25588 36662 25942
rect 36604 25296 36616 25588
rect 36650 25296 36662 25588
rect 36604 24942 36662 25296
rect 37662 25588 37720 25942
rect 37662 25296 37674 25588
rect 37708 25296 37720 25588
rect 37662 24942 37720 25296
rect 38720 25588 38778 25942
rect 38720 25296 38732 25588
rect 38766 25296 38778 25588
rect 38720 24942 38778 25296
rect 39778 25588 39836 25942
rect 39778 25296 39790 25588
rect 39824 25296 39836 25588
rect 39778 24942 39836 25296
rect 40978 25588 41036 25942
rect 40978 25296 40990 25588
rect 41024 25296 41036 25588
rect 40978 24942 41036 25296
rect 42036 25588 42094 25942
rect 42036 25296 42048 25588
rect 42082 25296 42094 25588
rect 42036 24942 42094 25296
rect 43094 25588 43152 25942
rect 43094 25296 43106 25588
rect 43140 25296 43152 25588
rect 43094 24942 43152 25296
rect 44152 25588 44210 25942
rect 44152 25296 44164 25588
rect 44198 25296 44210 25588
rect 44152 24942 44210 25296
rect 45210 25588 45268 25942
rect 45210 25296 45222 25588
rect 45256 25296 45268 25588
rect 45210 24942 45268 25296
rect 46268 25588 46326 25942
rect 46268 25296 46280 25588
rect 46314 25296 46326 25588
rect 46268 24942 46326 25296
rect 47566 25610 47624 25964
rect 47566 25318 47578 25610
rect 47612 25318 47624 25610
rect 47566 24964 47624 25318
rect 48624 25610 48682 25964
rect 48624 25318 48636 25610
rect 48670 25318 48682 25610
rect 48624 24964 48682 25318
rect 49682 25610 49740 25964
rect 49682 25318 49694 25610
rect 49728 25318 49740 25610
rect 49682 24964 49740 25318
rect 50740 25610 50798 25964
rect 50740 25318 50752 25610
rect 50786 25318 50798 25610
rect 50740 24964 50798 25318
rect 51798 25610 51856 25964
rect 51798 25318 51810 25610
rect 51844 25318 51856 25610
rect 51798 24964 51856 25318
rect 52856 25610 52914 25964
rect 52856 25318 52868 25610
rect 52902 25318 52914 25610
rect 52856 24964 52914 25318
rect 54080 25624 54138 25978
rect 54080 25332 54092 25624
rect 54126 25332 54138 25624
rect 54080 24978 54138 25332
rect 55138 25624 55196 25978
rect 55138 25332 55150 25624
rect 55184 25332 55196 25624
rect 55138 24978 55196 25332
rect 56196 25624 56254 25978
rect 56196 25332 56208 25624
rect 56242 25332 56254 25624
rect 56196 24978 56254 25332
rect 57254 25624 57312 25978
rect 57254 25332 57266 25624
rect 57300 25332 57312 25624
rect 57254 24978 57312 25332
rect 58312 25624 58370 25978
rect 58312 25332 58324 25624
rect 58358 25332 58370 25624
rect 58312 24978 58370 25332
rect 59370 25624 59428 25978
rect 59370 25332 59382 25624
rect 59416 25332 59428 25624
rect 59370 24978 59428 25332
rect 1946 24472 2004 24826
rect 1946 24180 1958 24472
rect 1992 24180 2004 24472
rect 1946 23826 2004 24180
rect 3004 24472 3062 24826
rect 3004 24180 3016 24472
rect 3050 24180 3062 24472
rect 3004 23826 3062 24180
rect 4062 24472 4120 24826
rect 4062 24180 4074 24472
rect 4108 24180 4120 24472
rect 4062 23826 4120 24180
rect 5120 24472 5178 24826
rect 5120 24180 5132 24472
rect 5166 24180 5178 24472
rect 5120 23826 5178 24180
rect 6178 24472 6236 24826
rect 6178 24180 6190 24472
rect 6224 24180 6236 24472
rect 6178 23826 6236 24180
rect 7236 24472 7294 24826
rect 7236 24180 7248 24472
rect 7282 24180 7294 24472
rect 8460 24480 8518 24834
rect 7236 23826 7294 24180
rect 1946 23378 2004 23732
rect 1946 23086 1958 23378
rect 1992 23086 2004 23378
rect 1946 22732 2004 23086
rect 3004 23378 3062 23732
rect 3004 23086 3016 23378
rect 3050 23086 3062 23378
rect 3004 22732 3062 23086
rect 4062 23378 4120 23732
rect 4062 23086 4074 23378
rect 4108 23086 4120 23378
rect 4062 22732 4120 23086
rect 5120 23378 5178 23732
rect 5120 23086 5132 23378
rect 5166 23086 5178 23378
rect 5120 22732 5178 23086
rect 6178 23378 6236 23732
rect 6178 23086 6190 23378
rect 6224 23086 6236 23378
rect 6178 22732 6236 23086
rect 7236 23378 7294 23732
rect 7236 23086 7248 23378
rect 7282 23086 7294 23378
rect 7236 22732 7294 23086
rect 8460 24188 8472 24480
rect 8506 24188 8518 24480
rect 8460 23834 8518 24188
rect 9518 24480 9576 24834
rect 9518 24188 9530 24480
rect 9564 24188 9576 24480
rect 9518 23834 9576 24188
rect 10576 24480 10634 24834
rect 10576 24188 10588 24480
rect 10622 24188 10634 24480
rect 10576 23834 10634 24188
rect 11634 24480 11692 24834
rect 11634 24188 11646 24480
rect 11680 24188 11692 24480
rect 11634 23834 11692 24188
rect 12692 24480 12750 24834
rect 12692 24188 12704 24480
rect 12738 24188 12750 24480
rect 12692 23834 12750 24188
rect 13750 24480 13808 24834
rect 13750 24188 13762 24480
rect 13796 24188 13808 24480
rect 14966 24488 15024 24842
rect 13750 23834 13808 24188
rect 1946 22284 2004 22638
rect 1946 21992 1958 22284
rect 1992 21992 2004 22284
rect 1946 21638 2004 21992
rect 3004 22284 3062 22638
rect 3004 21992 3016 22284
rect 3050 21992 3062 22284
rect 3004 21638 3062 21992
rect 4062 22284 4120 22638
rect 4062 21992 4074 22284
rect 4108 21992 4120 22284
rect 4062 21638 4120 21992
rect 5120 22284 5178 22638
rect 5120 21992 5132 22284
rect 5166 21992 5178 22284
rect 5120 21638 5178 21992
rect 6178 22284 6236 22638
rect 6178 21992 6190 22284
rect 6224 21992 6236 22284
rect 6178 21638 6236 21992
rect 7236 22284 7294 22638
rect 8460 23386 8518 23740
rect 8460 23094 8472 23386
rect 8506 23094 8518 23386
rect 8460 22740 8518 23094
rect 9518 23386 9576 23740
rect 9518 23094 9530 23386
rect 9564 23094 9576 23386
rect 9518 22740 9576 23094
rect 10576 23386 10634 23740
rect 10576 23094 10588 23386
rect 10622 23094 10634 23386
rect 10576 22740 10634 23094
rect 11634 23386 11692 23740
rect 11634 23094 11646 23386
rect 11680 23094 11692 23386
rect 11634 22740 11692 23094
rect 12692 23386 12750 23740
rect 12692 23094 12704 23386
rect 12738 23094 12750 23386
rect 12692 22740 12750 23094
rect 13750 23386 13808 23740
rect 13750 23094 13762 23386
rect 13796 23094 13808 23386
rect 13750 22740 13808 23094
rect 14966 24196 14978 24488
rect 15012 24196 15024 24488
rect 14966 23842 15024 24196
rect 16024 24488 16082 24842
rect 16024 24196 16036 24488
rect 16070 24196 16082 24488
rect 16024 23842 16082 24196
rect 17082 24488 17140 24842
rect 17082 24196 17094 24488
rect 17128 24196 17140 24488
rect 17082 23842 17140 24196
rect 18140 24488 18198 24842
rect 18140 24196 18152 24488
rect 18186 24196 18198 24488
rect 18140 23842 18198 24196
rect 19198 24488 19256 24842
rect 19198 24196 19210 24488
rect 19244 24196 19256 24488
rect 19198 23842 19256 24196
rect 20256 24488 20314 24842
rect 20256 24196 20268 24488
rect 20302 24196 20314 24488
rect 20256 23842 20314 24196
rect 21456 24472 21514 24826
rect 7236 21992 7248 22284
rect 7282 21992 7294 22284
rect 7236 21638 7294 21992
rect 8460 22292 8518 22646
rect 8460 22000 8472 22292
rect 8506 22000 8518 22292
rect 8460 21646 8518 22000
rect 9518 22292 9576 22646
rect 9518 22000 9530 22292
rect 9564 22000 9576 22292
rect 9518 21646 9576 22000
rect 10576 22292 10634 22646
rect 10576 22000 10588 22292
rect 10622 22000 10634 22292
rect 10576 21646 10634 22000
rect 11634 22292 11692 22646
rect 11634 22000 11646 22292
rect 11680 22000 11692 22292
rect 11634 21646 11692 22000
rect 12692 22292 12750 22646
rect 12692 22000 12704 22292
rect 12738 22000 12750 22292
rect 12692 21646 12750 22000
rect 13750 22292 13808 22646
rect 14966 23394 15024 23748
rect 14966 23102 14978 23394
rect 15012 23102 15024 23394
rect 14966 22748 15024 23102
rect 16024 23394 16082 23748
rect 16024 23102 16036 23394
rect 16070 23102 16082 23394
rect 16024 22748 16082 23102
rect 17082 23394 17140 23748
rect 17082 23102 17094 23394
rect 17128 23102 17140 23394
rect 17082 22748 17140 23102
rect 18140 23394 18198 23748
rect 18140 23102 18152 23394
rect 18186 23102 18198 23394
rect 18140 22748 18198 23102
rect 19198 23394 19256 23748
rect 19198 23102 19210 23394
rect 19244 23102 19256 23394
rect 19198 22748 19256 23102
rect 20256 23394 20314 23748
rect 20256 23102 20268 23394
rect 20302 23102 20314 23394
rect 20256 22748 20314 23102
rect 21456 24180 21468 24472
rect 21502 24180 21514 24472
rect 21456 23826 21514 24180
rect 22514 24472 22572 24826
rect 22514 24180 22526 24472
rect 22560 24180 22572 24472
rect 22514 23826 22572 24180
rect 23572 24472 23630 24826
rect 23572 24180 23584 24472
rect 23618 24180 23630 24472
rect 23572 23826 23630 24180
rect 24630 24472 24688 24826
rect 24630 24180 24642 24472
rect 24676 24180 24688 24472
rect 24630 23826 24688 24180
rect 25688 24472 25746 24826
rect 25688 24180 25700 24472
rect 25734 24180 25746 24472
rect 25688 23826 25746 24180
rect 26746 24472 26804 24826
rect 26746 24180 26758 24472
rect 26792 24180 26804 24472
rect 27978 24488 28036 24842
rect 26746 23826 26804 24180
rect 13750 22000 13762 22292
rect 13796 22000 13808 22292
rect 13750 21646 13808 22000
rect 14966 22300 15024 22654
rect 14966 22008 14978 22300
rect 15012 22008 15024 22300
rect 14966 21654 15024 22008
rect 16024 22300 16082 22654
rect 16024 22008 16036 22300
rect 16070 22008 16082 22300
rect 16024 21654 16082 22008
rect 17082 22300 17140 22654
rect 17082 22008 17094 22300
rect 17128 22008 17140 22300
rect 17082 21654 17140 22008
rect 18140 22300 18198 22654
rect 18140 22008 18152 22300
rect 18186 22008 18198 22300
rect 18140 21654 18198 22008
rect 19198 22300 19256 22654
rect 19198 22008 19210 22300
rect 19244 22008 19256 22300
rect 19198 21654 19256 22008
rect 20256 22300 20314 22654
rect 21456 23378 21514 23732
rect 21456 23086 21468 23378
rect 21502 23086 21514 23378
rect 21456 22732 21514 23086
rect 22514 23378 22572 23732
rect 22514 23086 22526 23378
rect 22560 23086 22572 23378
rect 22514 22732 22572 23086
rect 23572 23378 23630 23732
rect 23572 23086 23584 23378
rect 23618 23086 23630 23378
rect 23572 22732 23630 23086
rect 24630 23378 24688 23732
rect 24630 23086 24642 23378
rect 24676 23086 24688 23378
rect 24630 22732 24688 23086
rect 25688 23378 25746 23732
rect 25688 23086 25700 23378
rect 25734 23086 25746 23378
rect 25688 22732 25746 23086
rect 26746 23378 26804 23732
rect 26746 23086 26758 23378
rect 26792 23086 26804 23378
rect 26746 22732 26804 23086
rect 27978 24196 27990 24488
rect 28024 24196 28036 24488
rect 27978 23842 28036 24196
rect 29036 24488 29094 24842
rect 29036 24196 29048 24488
rect 29082 24196 29094 24488
rect 29036 23842 29094 24196
rect 30094 24488 30152 24842
rect 30094 24196 30106 24488
rect 30140 24196 30152 24488
rect 30094 23842 30152 24196
rect 31152 24488 31210 24842
rect 31152 24196 31164 24488
rect 31198 24196 31210 24488
rect 31152 23842 31210 24196
rect 32210 24488 32268 24842
rect 32210 24196 32222 24488
rect 32256 24196 32268 24488
rect 32210 23842 32268 24196
rect 33268 24488 33326 24842
rect 33268 24196 33280 24488
rect 33314 24196 33326 24488
rect 34488 24494 34546 24848
rect 33268 23842 33326 24196
rect 20256 22008 20268 22300
rect 20302 22008 20314 22300
rect 20256 21654 20314 22008
rect 21456 22284 21514 22638
rect 21456 21992 21468 22284
rect 21502 21992 21514 22284
rect 21456 21638 21514 21992
rect 22514 22284 22572 22638
rect 22514 21992 22526 22284
rect 22560 21992 22572 22284
rect 22514 21638 22572 21992
rect 23572 22284 23630 22638
rect 23572 21992 23584 22284
rect 23618 21992 23630 22284
rect 23572 21638 23630 21992
rect 24630 22284 24688 22638
rect 24630 21992 24642 22284
rect 24676 21992 24688 22284
rect 24630 21638 24688 21992
rect 25688 22284 25746 22638
rect 25688 21992 25700 22284
rect 25734 21992 25746 22284
rect 25688 21638 25746 21992
rect 26746 22284 26804 22638
rect 27978 23394 28036 23748
rect 27978 23102 27990 23394
rect 28024 23102 28036 23394
rect 27978 22748 28036 23102
rect 29036 23394 29094 23748
rect 29036 23102 29048 23394
rect 29082 23102 29094 23394
rect 29036 22748 29094 23102
rect 30094 23394 30152 23748
rect 30094 23102 30106 23394
rect 30140 23102 30152 23394
rect 30094 22748 30152 23102
rect 31152 23394 31210 23748
rect 31152 23102 31164 23394
rect 31198 23102 31210 23394
rect 31152 22748 31210 23102
rect 32210 23394 32268 23748
rect 32210 23102 32222 23394
rect 32256 23102 32268 23394
rect 32210 22748 32268 23102
rect 33268 23394 33326 23748
rect 33268 23102 33280 23394
rect 33314 23102 33326 23394
rect 33268 22748 33326 23102
rect 34488 24202 34500 24494
rect 34534 24202 34546 24494
rect 34488 23848 34546 24202
rect 35546 24494 35604 24848
rect 35546 24202 35558 24494
rect 35592 24202 35604 24494
rect 35546 23848 35604 24202
rect 36604 24494 36662 24848
rect 36604 24202 36616 24494
rect 36650 24202 36662 24494
rect 36604 23848 36662 24202
rect 37662 24494 37720 24848
rect 37662 24202 37674 24494
rect 37708 24202 37720 24494
rect 37662 23848 37720 24202
rect 38720 24494 38778 24848
rect 38720 24202 38732 24494
rect 38766 24202 38778 24494
rect 38720 23848 38778 24202
rect 39778 24494 39836 24848
rect 39778 24202 39790 24494
rect 39824 24202 39836 24494
rect 40978 24494 41036 24848
rect 39778 23848 39836 24202
rect 26746 21992 26758 22284
rect 26792 21992 26804 22284
rect 26746 21638 26804 21992
rect 27978 22300 28036 22654
rect 27978 22008 27990 22300
rect 28024 22008 28036 22300
rect 27978 21654 28036 22008
rect 29036 22300 29094 22654
rect 29036 22008 29048 22300
rect 29082 22008 29094 22300
rect 29036 21654 29094 22008
rect 30094 22300 30152 22654
rect 30094 22008 30106 22300
rect 30140 22008 30152 22300
rect 30094 21654 30152 22008
rect 31152 22300 31210 22654
rect 31152 22008 31164 22300
rect 31198 22008 31210 22300
rect 31152 21654 31210 22008
rect 32210 22300 32268 22654
rect 32210 22008 32222 22300
rect 32256 22008 32268 22300
rect 32210 21654 32268 22008
rect 33268 22300 33326 22654
rect 34488 23400 34546 23754
rect 34488 23108 34500 23400
rect 34534 23108 34546 23400
rect 34488 22754 34546 23108
rect 35546 23400 35604 23754
rect 35546 23108 35558 23400
rect 35592 23108 35604 23400
rect 35546 22754 35604 23108
rect 36604 23400 36662 23754
rect 36604 23108 36616 23400
rect 36650 23108 36662 23400
rect 36604 22754 36662 23108
rect 37662 23400 37720 23754
rect 37662 23108 37674 23400
rect 37708 23108 37720 23400
rect 37662 22754 37720 23108
rect 38720 23400 38778 23754
rect 38720 23108 38732 23400
rect 38766 23108 38778 23400
rect 38720 22754 38778 23108
rect 39778 23400 39836 23754
rect 39778 23108 39790 23400
rect 39824 23108 39836 23400
rect 39778 22754 39836 23108
rect 40978 24202 40990 24494
rect 41024 24202 41036 24494
rect 40978 23848 41036 24202
rect 42036 24494 42094 24848
rect 42036 24202 42048 24494
rect 42082 24202 42094 24494
rect 42036 23848 42094 24202
rect 43094 24494 43152 24848
rect 43094 24202 43106 24494
rect 43140 24202 43152 24494
rect 43094 23848 43152 24202
rect 44152 24494 44210 24848
rect 44152 24202 44164 24494
rect 44198 24202 44210 24494
rect 44152 23848 44210 24202
rect 45210 24494 45268 24848
rect 45210 24202 45222 24494
rect 45256 24202 45268 24494
rect 45210 23848 45268 24202
rect 46268 24494 46326 24848
rect 46268 24202 46280 24494
rect 46314 24202 46326 24494
rect 47566 24516 47624 24870
rect 46268 23848 46326 24202
rect 33268 22008 33280 22300
rect 33314 22008 33326 22300
rect 33268 21654 33326 22008
rect 34488 22306 34546 22660
rect 34488 22014 34500 22306
rect 34534 22014 34546 22306
rect 34488 21660 34546 22014
rect 35546 22306 35604 22660
rect 35546 22014 35558 22306
rect 35592 22014 35604 22306
rect 35546 21660 35604 22014
rect 36604 22306 36662 22660
rect 36604 22014 36616 22306
rect 36650 22014 36662 22306
rect 36604 21660 36662 22014
rect 37662 22306 37720 22660
rect 37662 22014 37674 22306
rect 37708 22014 37720 22306
rect 37662 21660 37720 22014
rect 38720 22306 38778 22660
rect 38720 22014 38732 22306
rect 38766 22014 38778 22306
rect 38720 21660 38778 22014
rect 39778 22306 39836 22660
rect 40978 23400 41036 23754
rect 40978 23108 40990 23400
rect 41024 23108 41036 23400
rect 40978 22754 41036 23108
rect 42036 23400 42094 23754
rect 42036 23108 42048 23400
rect 42082 23108 42094 23400
rect 42036 22754 42094 23108
rect 43094 23400 43152 23754
rect 43094 23108 43106 23400
rect 43140 23108 43152 23400
rect 43094 22754 43152 23108
rect 44152 23400 44210 23754
rect 44152 23108 44164 23400
rect 44198 23108 44210 23400
rect 44152 22754 44210 23108
rect 45210 23400 45268 23754
rect 45210 23108 45222 23400
rect 45256 23108 45268 23400
rect 45210 22754 45268 23108
rect 46268 23400 46326 23754
rect 46268 23108 46280 23400
rect 46314 23108 46326 23400
rect 46268 22754 46326 23108
rect 47566 24224 47578 24516
rect 47612 24224 47624 24516
rect 47566 23870 47624 24224
rect 48624 24516 48682 24870
rect 48624 24224 48636 24516
rect 48670 24224 48682 24516
rect 48624 23870 48682 24224
rect 49682 24516 49740 24870
rect 49682 24224 49694 24516
rect 49728 24224 49740 24516
rect 49682 23870 49740 24224
rect 50740 24516 50798 24870
rect 50740 24224 50752 24516
rect 50786 24224 50798 24516
rect 50740 23870 50798 24224
rect 51798 24516 51856 24870
rect 51798 24224 51810 24516
rect 51844 24224 51856 24516
rect 51798 23870 51856 24224
rect 52856 24516 52914 24870
rect 52856 24224 52868 24516
rect 52902 24224 52914 24516
rect 54080 24530 54138 24884
rect 52856 23870 52914 24224
rect 39778 22014 39790 22306
rect 39824 22014 39836 22306
rect 39778 21660 39836 22014
rect 40978 22306 41036 22660
rect 40978 22014 40990 22306
rect 41024 22014 41036 22306
rect 40978 21660 41036 22014
rect 42036 22306 42094 22660
rect 42036 22014 42048 22306
rect 42082 22014 42094 22306
rect 42036 21660 42094 22014
rect 43094 22306 43152 22660
rect 43094 22014 43106 22306
rect 43140 22014 43152 22306
rect 43094 21660 43152 22014
rect 44152 22306 44210 22660
rect 44152 22014 44164 22306
rect 44198 22014 44210 22306
rect 44152 21660 44210 22014
rect 45210 22306 45268 22660
rect 45210 22014 45222 22306
rect 45256 22014 45268 22306
rect 45210 21660 45268 22014
rect 46268 22306 46326 22660
rect 47566 23422 47624 23776
rect 47566 23130 47578 23422
rect 47612 23130 47624 23422
rect 47566 22776 47624 23130
rect 48624 23422 48682 23776
rect 48624 23130 48636 23422
rect 48670 23130 48682 23422
rect 48624 22776 48682 23130
rect 49682 23422 49740 23776
rect 49682 23130 49694 23422
rect 49728 23130 49740 23422
rect 49682 22776 49740 23130
rect 50740 23422 50798 23776
rect 50740 23130 50752 23422
rect 50786 23130 50798 23422
rect 50740 22776 50798 23130
rect 51798 23422 51856 23776
rect 51798 23130 51810 23422
rect 51844 23130 51856 23422
rect 51798 22776 51856 23130
rect 52856 23422 52914 23776
rect 52856 23130 52868 23422
rect 52902 23130 52914 23422
rect 52856 22776 52914 23130
rect 54080 24238 54092 24530
rect 54126 24238 54138 24530
rect 54080 23884 54138 24238
rect 55138 24530 55196 24884
rect 55138 24238 55150 24530
rect 55184 24238 55196 24530
rect 55138 23884 55196 24238
rect 56196 24530 56254 24884
rect 56196 24238 56208 24530
rect 56242 24238 56254 24530
rect 56196 23884 56254 24238
rect 57254 24530 57312 24884
rect 57254 24238 57266 24530
rect 57300 24238 57312 24530
rect 57254 23884 57312 24238
rect 58312 24530 58370 24884
rect 58312 24238 58324 24530
rect 58358 24238 58370 24530
rect 58312 23884 58370 24238
rect 59370 24530 59428 24884
rect 59370 24238 59382 24530
rect 59416 24238 59428 24530
rect 59370 23884 59428 24238
rect 46268 22014 46280 22306
rect 46314 22014 46326 22306
rect 46268 21660 46326 22014
rect 47566 22328 47624 22682
rect 47566 22036 47578 22328
rect 47612 22036 47624 22328
rect 47566 21682 47624 22036
rect 48624 22328 48682 22682
rect 48624 22036 48636 22328
rect 48670 22036 48682 22328
rect 48624 21682 48682 22036
rect 49682 22328 49740 22682
rect 49682 22036 49694 22328
rect 49728 22036 49740 22328
rect 49682 21682 49740 22036
rect 50740 22328 50798 22682
rect 50740 22036 50752 22328
rect 50786 22036 50798 22328
rect 50740 21682 50798 22036
rect 51798 22328 51856 22682
rect 51798 22036 51810 22328
rect 51844 22036 51856 22328
rect 51798 21682 51856 22036
rect 52856 22328 52914 22682
rect 54080 23436 54138 23790
rect 54080 23144 54092 23436
rect 54126 23144 54138 23436
rect 54080 22790 54138 23144
rect 55138 23436 55196 23790
rect 55138 23144 55150 23436
rect 55184 23144 55196 23436
rect 55138 22790 55196 23144
rect 56196 23436 56254 23790
rect 56196 23144 56208 23436
rect 56242 23144 56254 23436
rect 56196 22790 56254 23144
rect 57254 23436 57312 23790
rect 57254 23144 57266 23436
rect 57300 23144 57312 23436
rect 57254 22790 57312 23144
rect 58312 23436 58370 23790
rect 58312 23144 58324 23436
rect 58358 23144 58370 23436
rect 58312 22790 58370 23144
rect 59370 23436 59428 23790
rect 59370 23144 59382 23436
rect 59416 23144 59428 23436
rect 59370 22790 59428 23144
rect 52856 22036 52868 22328
rect 52902 22036 52914 22328
rect 52856 21682 52914 22036
rect 54080 22342 54138 22696
rect 54080 22050 54092 22342
rect 54126 22050 54138 22342
rect 54080 21696 54138 22050
rect 55138 22342 55196 22696
rect 55138 22050 55150 22342
rect 55184 22050 55196 22342
rect 55138 21696 55196 22050
rect 56196 22342 56254 22696
rect 56196 22050 56208 22342
rect 56242 22050 56254 22342
rect 56196 21696 56254 22050
rect 57254 22342 57312 22696
rect 57254 22050 57266 22342
rect 57300 22050 57312 22342
rect 57254 21696 57312 22050
rect 58312 22342 58370 22696
rect 58312 22050 58324 22342
rect 58358 22050 58370 22342
rect 58312 21696 58370 22050
rect 59370 22342 59428 22696
rect 59370 22050 59382 22342
rect 59416 22050 59428 22342
rect 59370 21696 59428 22050
rect 1946 21190 2004 21544
rect 1946 20898 1958 21190
rect 1992 20898 2004 21190
rect 1946 20544 2004 20898
rect 3004 21190 3062 21544
rect 3004 20898 3016 21190
rect 3050 20898 3062 21190
rect 3004 20544 3062 20898
rect 4062 21190 4120 21544
rect 4062 20898 4074 21190
rect 4108 20898 4120 21190
rect 4062 20544 4120 20898
rect 5120 21190 5178 21544
rect 5120 20898 5132 21190
rect 5166 20898 5178 21190
rect 5120 20544 5178 20898
rect 6178 21190 6236 21544
rect 6178 20898 6190 21190
rect 6224 20898 6236 21190
rect 6178 20544 6236 20898
rect 7236 21190 7294 21544
rect 7236 20898 7248 21190
rect 7282 20898 7294 21190
rect 7236 20544 7294 20898
rect 8460 21198 8518 21552
rect 8460 20906 8472 21198
rect 8506 20906 8518 21198
rect 8460 20552 8518 20906
rect 9518 21198 9576 21552
rect 9518 20906 9530 21198
rect 9564 20906 9576 21198
rect 9518 20552 9576 20906
rect 10576 21198 10634 21552
rect 10576 20906 10588 21198
rect 10622 20906 10634 21198
rect 10576 20552 10634 20906
rect 11634 21198 11692 21552
rect 11634 20906 11646 21198
rect 11680 20906 11692 21198
rect 11634 20552 11692 20906
rect 12692 21198 12750 21552
rect 12692 20906 12704 21198
rect 12738 20906 12750 21198
rect 12692 20552 12750 20906
rect 13750 21198 13808 21552
rect 13750 20906 13762 21198
rect 13796 20906 13808 21198
rect 13750 20552 13808 20906
rect 14966 21206 15024 21560
rect 14966 20914 14978 21206
rect 15012 20914 15024 21206
rect 14966 20560 15024 20914
rect 16024 21206 16082 21560
rect 16024 20914 16036 21206
rect 16070 20914 16082 21206
rect 16024 20560 16082 20914
rect 17082 21206 17140 21560
rect 17082 20914 17094 21206
rect 17128 20914 17140 21206
rect 17082 20560 17140 20914
rect 18140 21206 18198 21560
rect 18140 20914 18152 21206
rect 18186 20914 18198 21206
rect 18140 20560 18198 20914
rect 19198 21206 19256 21560
rect 19198 20914 19210 21206
rect 19244 20914 19256 21206
rect 19198 20560 19256 20914
rect 20256 21206 20314 21560
rect 20256 20914 20268 21206
rect 20302 20914 20314 21206
rect 20256 20560 20314 20914
rect 21456 21190 21514 21544
rect 21456 20898 21468 21190
rect 21502 20898 21514 21190
rect 21456 20544 21514 20898
rect 22514 21190 22572 21544
rect 22514 20898 22526 21190
rect 22560 20898 22572 21190
rect 22514 20544 22572 20898
rect 23572 21190 23630 21544
rect 23572 20898 23584 21190
rect 23618 20898 23630 21190
rect 23572 20544 23630 20898
rect 24630 21190 24688 21544
rect 24630 20898 24642 21190
rect 24676 20898 24688 21190
rect 24630 20544 24688 20898
rect 25688 21190 25746 21544
rect 25688 20898 25700 21190
rect 25734 20898 25746 21190
rect 25688 20544 25746 20898
rect 26746 21190 26804 21544
rect 26746 20898 26758 21190
rect 26792 20898 26804 21190
rect 26746 20544 26804 20898
rect 27978 21206 28036 21560
rect 27978 20914 27990 21206
rect 28024 20914 28036 21206
rect 27978 20560 28036 20914
rect 29036 21206 29094 21560
rect 29036 20914 29048 21206
rect 29082 20914 29094 21206
rect 29036 20560 29094 20914
rect 30094 21206 30152 21560
rect 30094 20914 30106 21206
rect 30140 20914 30152 21206
rect 30094 20560 30152 20914
rect 31152 21206 31210 21560
rect 31152 20914 31164 21206
rect 31198 20914 31210 21206
rect 31152 20560 31210 20914
rect 32210 21206 32268 21560
rect 32210 20914 32222 21206
rect 32256 20914 32268 21206
rect 32210 20560 32268 20914
rect 33268 21206 33326 21560
rect 33268 20914 33280 21206
rect 33314 20914 33326 21206
rect 33268 20560 33326 20914
rect 34488 21212 34546 21566
rect 34488 20920 34500 21212
rect 34534 20920 34546 21212
rect 34488 20566 34546 20920
rect 35546 21212 35604 21566
rect 35546 20920 35558 21212
rect 35592 20920 35604 21212
rect 35546 20566 35604 20920
rect 36604 21212 36662 21566
rect 36604 20920 36616 21212
rect 36650 20920 36662 21212
rect 36604 20566 36662 20920
rect 37662 21212 37720 21566
rect 37662 20920 37674 21212
rect 37708 20920 37720 21212
rect 37662 20566 37720 20920
rect 38720 21212 38778 21566
rect 38720 20920 38732 21212
rect 38766 20920 38778 21212
rect 38720 20566 38778 20920
rect 39778 21212 39836 21566
rect 39778 20920 39790 21212
rect 39824 20920 39836 21212
rect 39778 20566 39836 20920
rect 40978 21212 41036 21566
rect 40978 20920 40990 21212
rect 41024 20920 41036 21212
rect 40978 20566 41036 20920
rect 42036 21212 42094 21566
rect 42036 20920 42048 21212
rect 42082 20920 42094 21212
rect 42036 20566 42094 20920
rect 43094 21212 43152 21566
rect 43094 20920 43106 21212
rect 43140 20920 43152 21212
rect 43094 20566 43152 20920
rect 44152 21212 44210 21566
rect 44152 20920 44164 21212
rect 44198 20920 44210 21212
rect 44152 20566 44210 20920
rect 45210 21212 45268 21566
rect 45210 20920 45222 21212
rect 45256 20920 45268 21212
rect 45210 20566 45268 20920
rect 46268 21212 46326 21566
rect 46268 20920 46280 21212
rect 46314 20920 46326 21212
rect 46268 20566 46326 20920
rect 47566 21234 47624 21588
rect 47566 20942 47578 21234
rect 47612 20942 47624 21234
rect 47566 20588 47624 20942
rect 48624 21234 48682 21588
rect 48624 20942 48636 21234
rect 48670 20942 48682 21234
rect 48624 20588 48682 20942
rect 49682 21234 49740 21588
rect 49682 20942 49694 21234
rect 49728 20942 49740 21234
rect 49682 20588 49740 20942
rect 50740 21234 50798 21588
rect 50740 20942 50752 21234
rect 50786 20942 50798 21234
rect 50740 20588 50798 20942
rect 51798 21234 51856 21588
rect 51798 20942 51810 21234
rect 51844 20942 51856 21234
rect 51798 20588 51856 20942
rect 52856 21234 52914 21588
rect 52856 20942 52868 21234
rect 52902 20942 52914 21234
rect 52856 20588 52914 20942
rect 54080 21248 54138 21602
rect 54080 20956 54092 21248
rect 54126 20956 54138 21248
rect 54080 20602 54138 20956
rect 55138 21248 55196 21602
rect 55138 20956 55150 21248
rect 55184 20956 55196 21248
rect 55138 20602 55196 20956
rect 56196 21248 56254 21602
rect 56196 20956 56208 21248
rect 56242 20956 56254 21248
rect 56196 20602 56254 20956
rect 57254 21248 57312 21602
rect 57254 20956 57266 21248
rect 57300 20956 57312 21248
rect 57254 20602 57312 20956
rect 58312 21248 58370 21602
rect 58312 20956 58324 21248
rect 58358 20956 58370 21248
rect 58312 20602 58370 20956
rect 59370 21248 59428 21602
rect 59370 20956 59382 21248
rect 59416 20956 59428 21248
rect 59370 20602 59428 20956
rect 1946 19702 2004 20056
rect 1946 19410 1958 19702
rect 1992 19410 2004 19702
rect 1946 19056 2004 19410
rect 3004 19702 3062 20056
rect 3004 19410 3016 19702
rect 3050 19410 3062 19702
rect 3004 19056 3062 19410
rect 4062 19702 4120 20056
rect 4062 19410 4074 19702
rect 4108 19410 4120 19702
rect 4062 19056 4120 19410
rect 5120 19702 5178 20056
rect 5120 19410 5132 19702
rect 5166 19410 5178 19702
rect 5120 19056 5178 19410
rect 6178 19702 6236 20056
rect 6178 19410 6190 19702
rect 6224 19410 6236 19702
rect 6178 19056 6236 19410
rect 7236 19702 7294 20056
rect 7236 19410 7248 19702
rect 7282 19410 7294 19702
rect 7236 19056 7294 19410
rect 8460 19710 8518 20064
rect 8460 19418 8472 19710
rect 8506 19418 8518 19710
rect 8460 19064 8518 19418
rect 9518 19710 9576 20064
rect 9518 19418 9530 19710
rect 9564 19418 9576 19710
rect 9518 19064 9576 19418
rect 10576 19710 10634 20064
rect 10576 19418 10588 19710
rect 10622 19418 10634 19710
rect 10576 19064 10634 19418
rect 11634 19710 11692 20064
rect 11634 19418 11646 19710
rect 11680 19418 11692 19710
rect 11634 19064 11692 19418
rect 12692 19710 12750 20064
rect 12692 19418 12704 19710
rect 12738 19418 12750 19710
rect 12692 19064 12750 19418
rect 13750 19710 13808 20064
rect 13750 19418 13762 19710
rect 13796 19418 13808 19710
rect 13750 19064 13808 19418
rect 14966 19718 15024 20072
rect 14966 19426 14978 19718
rect 15012 19426 15024 19718
rect 14966 19072 15024 19426
rect 16024 19718 16082 20072
rect 16024 19426 16036 19718
rect 16070 19426 16082 19718
rect 16024 19072 16082 19426
rect 17082 19718 17140 20072
rect 17082 19426 17094 19718
rect 17128 19426 17140 19718
rect 17082 19072 17140 19426
rect 18140 19718 18198 20072
rect 18140 19426 18152 19718
rect 18186 19426 18198 19718
rect 18140 19072 18198 19426
rect 19198 19718 19256 20072
rect 19198 19426 19210 19718
rect 19244 19426 19256 19718
rect 19198 19072 19256 19426
rect 20256 19718 20314 20072
rect 20256 19426 20268 19718
rect 20302 19426 20314 19718
rect 20256 19072 20314 19426
rect 21456 19702 21514 20056
rect 21456 19410 21468 19702
rect 21502 19410 21514 19702
rect 21456 19056 21514 19410
rect 22514 19702 22572 20056
rect 22514 19410 22526 19702
rect 22560 19410 22572 19702
rect 22514 19056 22572 19410
rect 23572 19702 23630 20056
rect 23572 19410 23584 19702
rect 23618 19410 23630 19702
rect 23572 19056 23630 19410
rect 24630 19702 24688 20056
rect 24630 19410 24642 19702
rect 24676 19410 24688 19702
rect 24630 19056 24688 19410
rect 25688 19702 25746 20056
rect 25688 19410 25700 19702
rect 25734 19410 25746 19702
rect 25688 19056 25746 19410
rect 26746 19702 26804 20056
rect 26746 19410 26758 19702
rect 26792 19410 26804 19702
rect 26746 19056 26804 19410
rect 27978 19718 28036 20072
rect 27978 19426 27990 19718
rect 28024 19426 28036 19718
rect 27978 19072 28036 19426
rect 29036 19718 29094 20072
rect 29036 19426 29048 19718
rect 29082 19426 29094 19718
rect 29036 19072 29094 19426
rect 30094 19718 30152 20072
rect 30094 19426 30106 19718
rect 30140 19426 30152 19718
rect 30094 19072 30152 19426
rect 31152 19718 31210 20072
rect 31152 19426 31164 19718
rect 31198 19426 31210 19718
rect 31152 19072 31210 19426
rect 32210 19718 32268 20072
rect 32210 19426 32222 19718
rect 32256 19426 32268 19718
rect 32210 19072 32268 19426
rect 33268 19718 33326 20072
rect 33268 19426 33280 19718
rect 33314 19426 33326 19718
rect 33268 19072 33326 19426
rect 34488 19724 34546 20078
rect 34488 19432 34500 19724
rect 34534 19432 34546 19724
rect 34488 19078 34546 19432
rect 35546 19724 35604 20078
rect 35546 19432 35558 19724
rect 35592 19432 35604 19724
rect 35546 19078 35604 19432
rect 36604 19724 36662 20078
rect 36604 19432 36616 19724
rect 36650 19432 36662 19724
rect 36604 19078 36662 19432
rect 37662 19724 37720 20078
rect 37662 19432 37674 19724
rect 37708 19432 37720 19724
rect 37662 19078 37720 19432
rect 38720 19724 38778 20078
rect 38720 19432 38732 19724
rect 38766 19432 38778 19724
rect 38720 19078 38778 19432
rect 39778 19724 39836 20078
rect 39778 19432 39790 19724
rect 39824 19432 39836 19724
rect 39778 19078 39836 19432
rect 40978 19724 41036 20078
rect 40978 19432 40990 19724
rect 41024 19432 41036 19724
rect 40978 19078 41036 19432
rect 42036 19724 42094 20078
rect 42036 19432 42048 19724
rect 42082 19432 42094 19724
rect 42036 19078 42094 19432
rect 43094 19724 43152 20078
rect 43094 19432 43106 19724
rect 43140 19432 43152 19724
rect 43094 19078 43152 19432
rect 44152 19724 44210 20078
rect 44152 19432 44164 19724
rect 44198 19432 44210 19724
rect 44152 19078 44210 19432
rect 45210 19724 45268 20078
rect 45210 19432 45222 19724
rect 45256 19432 45268 19724
rect 45210 19078 45268 19432
rect 46268 19724 46326 20078
rect 46268 19432 46280 19724
rect 46314 19432 46326 19724
rect 46268 19078 46326 19432
rect 47566 19746 47624 20100
rect 47566 19454 47578 19746
rect 47612 19454 47624 19746
rect 47566 19100 47624 19454
rect 48624 19746 48682 20100
rect 48624 19454 48636 19746
rect 48670 19454 48682 19746
rect 48624 19100 48682 19454
rect 49682 19746 49740 20100
rect 49682 19454 49694 19746
rect 49728 19454 49740 19746
rect 49682 19100 49740 19454
rect 50740 19746 50798 20100
rect 50740 19454 50752 19746
rect 50786 19454 50798 19746
rect 50740 19100 50798 19454
rect 51798 19746 51856 20100
rect 51798 19454 51810 19746
rect 51844 19454 51856 19746
rect 51798 19100 51856 19454
rect 52856 19746 52914 20100
rect 52856 19454 52868 19746
rect 52902 19454 52914 19746
rect 52856 19100 52914 19454
rect 54080 19760 54138 20114
rect 54080 19468 54092 19760
rect 54126 19468 54138 19760
rect 54080 19114 54138 19468
rect 55138 19760 55196 20114
rect 55138 19468 55150 19760
rect 55184 19468 55196 19760
rect 55138 19114 55196 19468
rect 56196 19760 56254 20114
rect 56196 19468 56208 19760
rect 56242 19468 56254 19760
rect 56196 19114 56254 19468
rect 57254 19760 57312 20114
rect 57254 19468 57266 19760
rect 57300 19468 57312 19760
rect 57254 19114 57312 19468
rect 58312 19760 58370 20114
rect 58312 19468 58324 19760
rect 58358 19468 58370 19760
rect 58312 19114 58370 19468
rect 59370 19760 59428 20114
rect 59370 19468 59382 19760
rect 59416 19468 59428 19760
rect 59370 19114 59428 19468
rect 1946 18608 2004 18962
rect 1946 18316 1958 18608
rect 1992 18316 2004 18608
rect 1946 17962 2004 18316
rect 3004 18608 3062 18962
rect 3004 18316 3016 18608
rect 3050 18316 3062 18608
rect 3004 17962 3062 18316
rect 4062 18608 4120 18962
rect 4062 18316 4074 18608
rect 4108 18316 4120 18608
rect 4062 17962 4120 18316
rect 5120 18608 5178 18962
rect 5120 18316 5132 18608
rect 5166 18316 5178 18608
rect 5120 17962 5178 18316
rect 6178 18608 6236 18962
rect 6178 18316 6190 18608
rect 6224 18316 6236 18608
rect 6178 17962 6236 18316
rect 7236 18608 7294 18962
rect 7236 18316 7248 18608
rect 7282 18316 7294 18608
rect 8460 18616 8518 18970
rect 7236 17962 7294 18316
rect 1946 17514 2004 17868
rect 1946 17222 1958 17514
rect 1992 17222 2004 17514
rect 1946 16868 2004 17222
rect 3004 17514 3062 17868
rect 3004 17222 3016 17514
rect 3050 17222 3062 17514
rect 3004 16868 3062 17222
rect 4062 17514 4120 17868
rect 4062 17222 4074 17514
rect 4108 17222 4120 17514
rect 4062 16868 4120 17222
rect 5120 17514 5178 17868
rect 5120 17222 5132 17514
rect 5166 17222 5178 17514
rect 5120 16868 5178 17222
rect 6178 17514 6236 17868
rect 6178 17222 6190 17514
rect 6224 17222 6236 17514
rect 6178 16868 6236 17222
rect 7236 17514 7294 17868
rect 7236 17222 7248 17514
rect 7282 17222 7294 17514
rect 7236 16868 7294 17222
rect 8460 18324 8472 18616
rect 8506 18324 8518 18616
rect 8460 17970 8518 18324
rect 9518 18616 9576 18970
rect 9518 18324 9530 18616
rect 9564 18324 9576 18616
rect 9518 17970 9576 18324
rect 10576 18616 10634 18970
rect 10576 18324 10588 18616
rect 10622 18324 10634 18616
rect 10576 17970 10634 18324
rect 11634 18616 11692 18970
rect 11634 18324 11646 18616
rect 11680 18324 11692 18616
rect 11634 17970 11692 18324
rect 12692 18616 12750 18970
rect 12692 18324 12704 18616
rect 12738 18324 12750 18616
rect 12692 17970 12750 18324
rect 13750 18616 13808 18970
rect 13750 18324 13762 18616
rect 13796 18324 13808 18616
rect 14966 18624 15024 18978
rect 13750 17970 13808 18324
rect 1946 16420 2004 16774
rect 1946 16128 1958 16420
rect 1992 16128 2004 16420
rect 1946 15774 2004 16128
rect 3004 16420 3062 16774
rect 3004 16128 3016 16420
rect 3050 16128 3062 16420
rect 3004 15774 3062 16128
rect 4062 16420 4120 16774
rect 4062 16128 4074 16420
rect 4108 16128 4120 16420
rect 4062 15774 4120 16128
rect 5120 16420 5178 16774
rect 5120 16128 5132 16420
rect 5166 16128 5178 16420
rect 5120 15774 5178 16128
rect 6178 16420 6236 16774
rect 6178 16128 6190 16420
rect 6224 16128 6236 16420
rect 6178 15774 6236 16128
rect 7236 16420 7294 16774
rect 8460 17522 8518 17876
rect 8460 17230 8472 17522
rect 8506 17230 8518 17522
rect 8460 16876 8518 17230
rect 9518 17522 9576 17876
rect 9518 17230 9530 17522
rect 9564 17230 9576 17522
rect 9518 16876 9576 17230
rect 10576 17522 10634 17876
rect 10576 17230 10588 17522
rect 10622 17230 10634 17522
rect 10576 16876 10634 17230
rect 11634 17522 11692 17876
rect 11634 17230 11646 17522
rect 11680 17230 11692 17522
rect 11634 16876 11692 17230
rect 12692 17522 12750 17876
rect 12692 17230 12704 17522
rect 12738 17230 12750 17522
rect 12692 16876 12750 17230
rect 13750 17522 13808 17876
rect 13750 17230 13762 17522
rect 13796 17230 13808 17522
rect 13750 16876 13808 17230
rect 14966 18332 14978 18624
rect 15012 18332 15024 18624
rect 14966 17978 15024 18332
rect 16024 18624 16082 18978
rect 16024 18332 16036 18624
rect 16070 18332 16082 18624
rect 16024 17978 16082 18332
rect 17082 18624 17140 18978
rect 17082 18332 17094 18624
rect 17128 18332 17140 18624
rect 17082 17978 17140 18332
rect 18140 18624 18198 18978
rect 18140 18332 18152 18624
rect 18186 18332 18198 18624
rect 18140 17978 18198 18332
rect 19198 18624 19256 18978
rect 19198 18332 19210 18624
rect 19244 18332 19256 18624
rect 19198 17978 19256 18332
rect 20256 18624 20314 18978
rect 20256 18332 20268 18624
rect 20302 18332 20314 18624
rect 20256 17978 20314 18332
rect 21456 18608 21514 18962
rect 7236 16128 7248 16420
rect 7282 16128 7294 16420
rect 7236 15774 7294 16128
rect 8460 16428 8518 16782
rect 8460 16136 8472 16428
rect 8506 16136 8518 16428
rect 8460 15782 8518 16136
rect 9518 16428 9576 16782
rect 9518 16136 9530 16428
rect 9564 16136 9576 16428
rect 9518 15782 9576 16136
rect 10576 16428 10634 16782
rect 10576 16136 10588 16428
rect 10622 16136 10634 16428
rect 10576 15782 10634 16136
rect 11634 16428 11692 16782
rect 11634 16136 11646 16428
rect 11680 16136 11692 16428
rect 11634 15782 11692 16136
rect 12692 16428 12750 16782
rect 12692 16136 12704 16428
rect 12738 16136 12750 16428
rect 12692 15782 12750 16136
rect 13750 16428 13808 16782
rect 14966 17530 15024 17884
rect 14966 17238 14978 17530
rect 15012 17238 15024 17530
rect 14966 16884 15024 17238
rect 16024 17530 16082 17884
rect 16024 17238 16036 17530
rect 16070 17238 16082 17530
rect 16024 16884 16082 17238
rect 17082 17530 17140 17884
rect 17082 17238 17094 17530
rect 17128 17238 17140 17530
rect 17082 16884 17140 17238
rect 18140 17530 18198 17884
rect 18140 17238 18152 17530
rect 18186 17238 18198 17530
rect 18140 16884 18198 17238
rect 19198 17530 19256 17884
rect 19198 17238 19210 17530
rect 19244 17238 19256 17530
rect 19198 16884 19256 17238
rect 20256 17530 20314 17884
rect 20256 17238 20268 17530
rect 20302 17238 20314 17530
rect 20256 16884 20314 17238
rect 21456 18316 21468 18608
rect 21502 18316 21514 18608
rect 21456 17962 21514 18316
rect 22514 18608 22572 18962
rect 22514 18316 22526 18608
rect 22560 18316 22572 18608
rect 22514 17962 22572 18316
rect 23572 18608 23630 18962
rect 23572 18316 23584 18608
rect 23618 18316 23630 18608
rect 23572 17962 23630 18316
rect 24630 18608 24688 18962
rect 24630 18316 24642 18608
rect 24676 18316 24688 18608
rect 24630 17962 24688 18316
rect 25688 18608 25746 18962
rect 25688 18316 25700 18608
rect 25734 18316 25746 18608
rect 25688 17962 25746 18316
rect 26746 18608 26804 18962
rect 26746 18316 26758 18608
rect 26792 18316 26804 18608
rect 27978 18624 28036 18978
rect 26746 17962 26804 18316
rect 13750 16136 13762 16428
rect 13796 16136 13808 16428
rect 13750 15782 13808 16136
rect 14966 16436 15024 16790
rect 14966 16144 14978 16436
rect 15012 16144 15024 16436
rect 14966 15790 15024 16144
rect 16024 16436 16082 16790
rect 16024 16144 16036 16436
rect 16070 16144 16082 16436
rect 16024 15790 16082 16144
rect 17082 16436 17140 16790
rect 17082 16144 17094 16436
rect 17128 16144 17140 16436
rect 17082 15790 17140 16144
rect 18140 16436 18198 16790
rect 18140 16144 18152 16436
rect 18186 16144 18198 16436
rect 18140 15790 18198 16144
rect 19198 16436 19256 16790
rect 19198 16144 19210 16436
rect 19244 16144 19256 16436
rect 19198 15790 19256 16144
rect 20256 16436 20314 16790
rect 21456 17514 21514 17868
rect 21456 17222 21468 17514
rect 21502 17222 21514 17514
rect 21456 16868 21514 17222
rect 22514 17514 22572 17868
rect 22514 17222 22526 17514
rect 22560 17222 22572 17514
rect 22514 16868 22572 17222
rect 23572 17514 23630 17868
rect 23572 17222 23584 17514
rect 23618 17222 23630 17514
rect 23572 16868 23630 17222
rect 24630 17514 24688 17868
rect 24630 17222 24642 17514
rect 24676 17222 24688 17514
rect 24630 16868 24688 17222
rect 25688 17514 25746 17868
rect 25688 17222 25700 17514
rect 25734 17222 25746 17514
rect 25688 16868 25746 17222
rect 26746 17514 26804 17868
rect 26746 17222 26758 17514
rect 26792 17222 26804 17514
rect 26746 16868 26804 17222
rect 27978 18332 27990 18624
rect 28024 18332 28036 18624
rect 27978 17978 28036 18332
rect 29036 18624 29094 18978
rect 29036 18332 29048 18624
rect 29082 18332 29094 18624
rect 29036 17978 29094 18332
rect 30094 18624 30152 18978
rect 30094 18332 30106 18624
rect 30140 18332 30152 18624
rect 30094 17978 30152 18332
rect 31152 18624 31210 18978
rect 31152 18332 31164 18624
rect 31198 18332 31210 18624
rect 31152 17978 31210 18332
rect 32210 18624 32268 18978
rect 32210 18332 32222 18624
rect 32256 18332 32268 18624
rect 32210 17978 32268 18332
rect 33268 18624 33326 18978
rect 33268 18332 33280 18624
rect 33314 18332 33326 18624
rect 34488 18630 34546 18984
rect 33268 17978 33326 18332
rect 20256 16144 20268 16436
rect 20302 16144 20314 16436
rect 20256 15790 20314 16144
rect 21456 16420 21514 16774
rect 21456 16128 21468 16420
rect 21502 16128 21514 16420
rect 21456 15774 21514 16128
rect 22514 16420 22572 16774
rect 22514 16128 22526 16420
rect 22560 16128 22572 16420
rect 22514 15774 22572 16128
rect 23572 16420 23630 16774
rect 23572 16128 23584 16420
rect 23618 16128 23630 16420
rect 23572 15774 23630 16128
rect 24630 16420 24688 16774
rect 24630 16128 24642 16420
rect 24676 16128 24688 16420
rect 24630 15774 24688 16128
rect 25688 16420 25746 16774
rect 25688 16128 25700 16420
rect 25734 16128 25746 16420
rect 25688 15774 25746 16128
rect 26746 16420 26804 16774
rect 27978 17530 28036 17884
rect 27978 17238 27990 17530
rect 28024 17238 28036 17530
rect 27978 16884 28036 17238
rect 29036 17530 29094 17884
rect 29036 17238 29048 17530
rect 29082 17238 29094 17530
rect 29036 16884 29094 17238
rect 30094 17530 30152 17884
rect 30094 17238 30106 17530
rect 30140 17238 30152 17530
rect 30094 16884 30152 17238
rect 31152 17530 31210 17884
rect 31152 17238 31164 17530
rect 31198 17238 31210 17530
rect 31152 16884 31210 17238
rect 32210 17530 32268 17884
rect 32210 17238 32222 17530
rect 32256 17238 32268 17530
rect 32210 16884 32268 17238
rect 33268 17530 33326 17884
rect 33268 17238 33280 17530
rect 33314 17238 33326 17530
rect 33268 16884 33326 17238
rect 34488 18338 34500 18630
rect 34534 18338 34546 18630
rect 34488 17984 34546 18338
rect 35546 18630 35604 18984
rect 35546 18338 35558 18630
rect 35592 18338 35604 18630
rect 35546 17984 35604 18338
rect 36604 18630 36662 18984
rect 36604 18338 36616 18630
rect 36650 18338 36662 18630
rect 36604 17984 36662 18338
rect 37662 18630 37720 18984
rect 37662 18338 37674 18630
rect 37708 18338 37720 18630
rect 37662 17984 37720 18338
rect 38720 18630 38778 18984
rect 38720 18338 38732 18630
rect 38766 18338 38778 18630
rect 38720 17984 38778 18338
rect 39778 18630 39836 18984
rect 39778 18338 39790 18630
rect 39824 18338 39836 18630
rect 40978 18630 41036 18984
rect 39778 17984 39836 18338
rect 26746 16128 26758 16420
rect 26792 16128 26804 16420
rect 26746 15774 26804 16128
rect 27978 16436 28036 16790
rect 27978 16144 27990 16436
rect 28024 16144 28036 16436
rect 27978 15790 28036 16144
rect 29036 16436 29094 16790
rect 29036 16144 29048 16436
rect 29082 16144 29094 16436
rect 29036 15790 29094 16144
rect 30094 16436 30152 16790
rect 30094 16144 30106 16436
rect 30140 16144 30152 16436
rect 30094 15790 30152 16144
rect 31152 16436 31210 16790
rect 31152 16144 31164 16436
rect 31198 16144 31210 16436
rect 31152 15790 31210 16144
rect 32210 16436 32268 16790
rect 32210 16144 32222 16436
rect 32256 16144 32268 16436
rect 32210 15790 32268 16144
rect 33268 16436 33326 16790
rect 34488 17536 34546 17890
rect 34488 17244 34500 17536
rect 34534 17244 34546 17536
rect 34488 16890 34546 17244
rect 35546 17536 35604 17890
rect 35546 17244 35558 17536
rect 35592 17244 35604 17536
rect 35546 16890 35604 17244
rect 36604 17536 36662 17890
rect 36604 17244 36616 17536
rect 36650 17244 36662 17536
rect 36604 16890 36662 17244
rect 37662 17536 37720 17890
rect 37662 17244 37674 17536
rect 37708 17244 37720 17536
rect 37662 16890 37720 17244
rect 38720 17536 38778 17890
rect 38720 17244 38732 17536
rect 38766 17244 38778 17536
rect 38720 16890 38778 17244
rect 39778 17536 39836 17890
rect 39778 17244 39790 17536
rect 39824 17244 39836 17536
rect 39778 16890 39836 17244
rect 40978 18338 40990 18630
rect 41024 18338 41036 18630
rect 40978 17984 41036 18338
rect 42036 18630 42094 18984
rect 42036 18338 42048 18630
rect 42082 18338 42094 18630
rect 42036 17984 42094 18338
rect 43094 18630 43152 18984
rect 43094 18338 43106 18630
rect 43140 18338 43152 18630
rect 43094 17984 43152 18338
rect 44152 18630 44210 18984
rect 44152 18338 44164 18630
rect 44198 18338 44210 18630
rect 44152 17984 44210 18338
rect 45210 18630 45268 18984
rect 45210 18338 45222 18630
rect 45256 18338 45268 18630
rect 45210 17984 45268 18338
rect 46268 18630 46326 18984
rect 46268 18338 46280 18630
rect 46314 18338 46326 18630
rect 47566 18652 47624 19006
rect 46268 17984 46326 18338
rect 33268 16144 33280 16436
rect 33314 16144 33326 16436
rect 33268 15790 33326 16144
rect 34488 16442 34546 16796
rect 34488 16150 34500 16442
rect 34534 16150 34546 16442
rect 34488 15796 34546 16150
rect 35546 16442 35604 16796
rect 35546 16150 35558 16442
rect 35592 16150 35604 16442
rect 35546 15796 35604 16150
rect 36604 16442 36662 16796
rect 36604 16150 36616 16442
rect 36650 16150 36662 16442
rect 36604 15796 36662 16150
rect 37662 16442 37720 16796
rect 37662 16150 37674 16442
rect 37708 16150 37720 16442
rect 37662 15796 37720 16150
rect 38720 16442 38778 16796
rect 38720 16150 38732 16442
rect 38766 16150 38778 16442
rect 38720 15796 38778 16150
rect 39778 16442 39836 16796
rect 40978 17536 41036 17890
rect 40978 17244 40990 17536
rect 41024 17244 41036 17536
rect 40978 16890 41036 17244
rect 42036 17536 42094 17890
rect 42036 17244 42048 17536
rect 42082 17244 42094 17536
rect 42036 16890 42094 17244
rect 43094 17536 43152 17890
rect 43094 17244 43106 17536
rect 43140 17244 43152 17536
rect 43094 16890 43152 17244
rect 44152 17536 44210 17890
rect 44152 17244 44164 17536
rect 44198 17244 44210 17536
rect 44152 16890 44210 17244
rect 45210 17536 45268 17890
rect 45210 17244 45222 17536
rect 45256 17244 45268 17536
rect 45210 16890 45268 17244
rect 46268 17536 46326 17890
rect 46268 17244 46280 17536
rect 46314 17244 46326 17536
rect 46268 16890 46326 17244
rect 47566 18360 47578 18652
rect 47612 18360 47624 18652
rect 47566 18006 47624 18360
rect 48624 18652 48682 19006
rect 48624 18360 48636 18652
rect 48670 18360 48682 18652
rect 48624 18006 48682 18360
rect 49682 18652 49740 19006
rect 49682 18360 49694 18652
rect 49728 18360 49740 18652
rect 49682 18006 49740 18360
rect 50740 18652 50798 19006
rect 50740 18360 50752 18652
rect 50786 18360 50798 18652
rect 50740 18006 50798 18360
rect 51798 18652 51856 19006
rect 51798 18360 51810 18652
rect 51844 18360 51856 18652
rect 51798 18006 51856 18360
rect 52856 18652 52914 19006
rect 52856 18360 52868 18652
rect 52902 18360 52914 18652
rect 54080 18666 54138 19020
rect 52856 18006 52914 18360
rect 39778 16150 39790 16442
rect 39824 16150 39836 16442
rect 39778 15796 39836 16150
rect 40978 16442 41036 16796
rect 40978 16150 40990 16442
rect 41024 16150 41036 16442
rect 40978 15796 41036 16150
rect 42036 16442 42094 16796
rect 42036 16150 42048 16442
rect 42082 16150 42094 16442
rect 42036 15796 42094 16150
rect 43094 16442 43152 16796
rect 43094 16150 43106 16442
rect 43140 16150 43152 16442
rect 43094 15796 43152 16150
rect 44152 16442 44210 16796
rect 44152 16150 44164 16442
rect 44198 16150 44210 16442
rect 44152 15796 44210 16150
rect 45210 16442 45268 16796
rect 45210 16150 45222 16442
rect 45256 16150 45268 16442
rect 45210 15796 45268 16150
rect 46268 16442 46326 16796
rect 47566 17558 47624 17912
rect 47566 17266 47578 17558
rect 47612 17266 47624 17558
rect 47566 16912 47624 17266
rect 48624 17558 48682 17912
rect 48624 17266 48636 17558
rect 48670 17266 48682 17558
rect 48624 16912 48682 17266
rect 49682 17558 49740 17912
rect 49682 17266 49694 17558
rect 49728 17266 49740 17558
rect 49682 16912 49740 17266
rect 50740 17558 50798 17912
rect 50740 17266 50752 17558
rect 50786 17266 50798 17558
rect 50740 16912 50798 17266
rect 51798 17558 51856 17912
rect 51798 17266 51810 17558
rect 51844 17266 51856 17558
rect 51798 16912 51856 17266
rect 52856 17558 52914 17912
rect 52856 17266 52868 17558
rect 52902 17266 52914 17558
rect 52856 16912 52914 17266
rect 54080 18374 54092 18666
rect 54126 18374 54138 18666
rect 54080 18020 54138 18374
rect 55138 18666 55196 19020
rect 55138 18374 55150 18666
rect 55184 18374 55196 18666
rect 55138 18020 55196 18374
rect 56196 18666 56254 19020
rect 56196 18374 56208 18666
rect 56242 18374 56254 18666
rect 56196 18020 56254 18374
rect 57254 18666 57312 19020
rect 57254 18374 57266 18666
rect 57300 18374 57312 18666
rect 57254 18020 57312 18374
rect 58312 18666 58370 19020
rect 58312 18374 58324 18666
rect 58358 18374 58370 18666
rect 58312 18020 58370 18374
rect 59370 18666 59428 19020
rect 59370 18374 59382 18666
rect 59416 18374 59428 18666
rect 59370 18020 59428 18374
rect 46268 16150 46280 16442
rect 46314 16150 46326 16442
rect 46268 15796 46326 16150
rect 47566 16464 47624 16818
rect 47566 16172 47578 16464
rect 47612 16172 47624 16464
rect 47566 15818 47624 16172
rect 48624 16464 48682 16818
rect 48624 16172 48636 16464
rect 48670 16172 48682 16464
rect 48624 15818 48682 16172
rect 49682 16464 49740 16818
rect 49682 16172 49694 16464
rect 49728 16172 49740 16464
rect 49682 15818 49740 16172
rect 50740 16464 50798 16818
rect 50740 16172 50752 16464
rect 50786 16172 50798 16464
rect 50740 15818 50798 16172
rect 51798 16464 51856 16818
rect 51798 16172 51810 16464
rect 51844 16172 51856 16464
rect 51798 15818 51856 16172
rect 52856 16464 52914 16818
rect 54080 17572 54138 17926
rect 54080 17280 54092 17572
rect 54126 17280 54138 17572
rect 54080 16926 54138 17280
rect 55138 17572 55196 17926
rect 55138 17280 55150 17572
rect 55184 17280 55196 17572
rect 55138 16926 55196 17280
rect 56196 17572 56254 17926
rect 56196 17280 56208 17572
rect 56242 17280 56254 17572
rect 56196 16926 56254 17280
rect 57254 17572 57312 17926
rect 57254 17280 57266 17572
rect 57300 17280 57312 17572
rect 57254 16926 57312 17280
rect 58312 17572 58370 17926
rect 58312 17280 58324 17572
rect 58358 17280 58370 17572
rect 58312 16926 58370 17280
rect 59370 17572 59428 17926
rect 59370 17280 59382 17572
rect 59416 17280 59428 17572
rect 59370 16926 59428 17280
rect 52856 16172 52868 16464
rect 52902 16172 52914 16464
rect 52856 15818 52914 16172
rect 54080 16478 54138 16832
rect 54080 16186 54092 16478
rect 54126 16186 54138 16478
rect 54080 15832 54138 16186
rect 55138 16478 55196 16832
rect 55138 16186 55150 16478
rect 55184 16186 55196 16478
rect 55138 15832 55196 16186
rect 56196 16478 56254 16832
rect 56196 16186 56208 16478
rect 56242 16186 56254 16478
rect 56196 15832 56254 16186
rect 57254 16478 57312 16832
rect 57254 16186 57266 16478
rect 57300 16186 57312 16478
rect 57254 15832 57312 16186
rect 58312 16478 58370 16832
rect 58312 16186 58324 16478
rect 58358 16186 58370 16478
rect 58312 15832 58370 16186
rect 59370 16478 59428 16832
rect 59370 16186 59382 16478
rect 59416 16186 59428 16478
rect 59370 15832 59428 16186
rect 1946 15326 2004 15680
rect 1946 15034 1958 15326
rect 1992 15034 2004 15326
rect 1946 14680 2004 15034
rect 3004 15326 3062 15680
rect 3004 15034 3016 15326
rect 3050 15034 3062 15326
rect 3004 14680 3062 15034
rect 4062 15326 4120 15680
rect 4062 15034 4074 15326
rect 4108 15034 4120 15326
rect 4062 14680 4120 15034
rect 5120 15326 5178 15680
rect 5120 15034 5132 15326
rect 5166 15034 5178 15326
rect 5120 14680 5178 15034
rect 6178 15326 6236 15680
rect 6178 15034 6190 15326
rect 6224 15034 6236 15326
rect 6178 14680 6236 15034
rect 7236 15326 7294 15680
rect 7236 15034 7248 15326
rect 7282 15034 7294 15326
rect 7236 14680 7294 15034
rect 8460 15334 8518 15688
rect 8460 15042 8472 15334
rect 8506 15042 8518 15334
rect 8460 14688 8518 15042
rect 9518 15334 9576 15688
rect 9518 15042 9530 15334
rect 9564 15042 9576 15334
rect 9518 14688 9576 15042
rect 10576 15334 10634 15688
rect 10576 15042 10588 15334
rect 10622 15042 10634 15334
rect 10576 14688 10634 15042
rect 11634 15334 11692 15688
rect 11634 15042 11646 15334
rect 11680 15042 11692 15334
rect 11634 14688 11692 15042
rect 12692 15334 12750 15688
rect 12692 15042 12704 15334
rect 12738 15042 12750 15334
rect 12692 14688 12750 15042
rect 13750 15334 13808 15688
rect 13750 15042 13762 15334
rect 13796 15042 13808 15334
rect 13750 14688 13808 15042
rect 14966 15342 15024 15696
rect 14966 15050 14978 15342
rect 15012 15050 15024 15342
rect 14966 14696 15024 15050
rect 16024 15342 16082 15696
rect 16024 15050 16036 15342
rect 16070 15050 16082 15342
rect 16024 14696 16082 15050
rect 17082 15342 17140 15696
rect 17082 15050 17094 15342
rect 17128 15050 17140 15342
rect 17082 14696 17140 15050
rect 18140 15342 18198 15696
rect 18140 15050 18152 15342
rect 18186 15050 18198 15342
rect 18140 14696 18198 15050
rect 19198 15342 19256 15696
rect 19198 15050 19210 15342
rect 19244 15050 19256 15342
rect 19198 14696 19256 15050
rect 20256 15342 20314 15696
rect 20256 15050 20268 15342
rect 20302 15050 20314 15342
rect 20256 14696 20314 15050
rect 21456 15326 21514 15680
rect 21456 15034 21468 15326
rect 21502 15034 21514 15326
rect 21456 14680 21514 15034
rect 22514 15326 22572 15680
rect 22514 15034 22526 15326
rect 22560 15034 22572 15326
rect 22514 14680 22572 15034
rect 23572 15326 23630 15680
rect 23572 15034 23584 15326
rect 23618 15034 23630 15326
rect 23572 14680 23630 15034
rect 24630 15326 24688 15680
rect 24630 15034 24642 15326
rect 24676 15034 24688 15326
rect 24630 14680 24688 15034
rect 25688 15326 25746 15680
rect 25688 15034 25700 15326
rect 25734 15034 25746 15326
rect 25688 14680 25746 15034
rect 26746 15326 26804 15680
rect 26746 15034 26758 15326
rect 26792 15034 26804 15326
rect 26746 14680 26804 15034
rect 27978 15342 28036 15696
rect 27978 15050 27990 15342
rect 28024 15050 28036 15342
rect 27978 14696 28036 15050
rect 29036 15342 29094 15696
rect 29036 15050 29048 15342
rect 29082 15050 29094 15342
rect 29036 14696 29094 15050
rect 30094 15342 30152 15696
rect 30094 15050 30106 15342
rect 30140 15050 30152 15342
rect 30094 14696 30152 15050
rect 31152 15342 31210 15696
rect 31152 15050 31164 15342
rect 31198 15050 31210 15342
rect 31152 14696 31210 15050
rect 32210 15342 32268 15696
rect 32210 15050 32222 15342
rect 32256 15050 32268 15342
rect 32210 14696 32268 15050
rect 33268 15342 33326 15696
rect 33268 15050 33280 15342
rect 33314 15050 33326 15342
rect 33268 14696 33326 15050
rect 34488 15348 34546 15702
rect 34488 15056 34500 15348
rect 34534 15056 34546 15348
rect 34488 14702 34546 15056
rect 35546 15348 35604 15702
rect 35546 15056 35558 15348
rect 35592 15056 35604 15348
rect 35546 14702 35604 15056
rect 36604 15348 36662 15702
rect 36604 15056 36616 15348
rect 36650 15056 36662 15348
rect 36604 14702 36662 15056
rect 37662 15348 37720 15702
rect 37662 15056 37674 15348
rect 37708 15056 37720 15348
rect 37662 14702 37720 15056
rect 38720 15348 38778 15702
rect 38720 15056 38732 15348
rect 38766 15056 38778 15348
rect 38720 14702 38778 15056
rect 39778 15348 39836 15702
rect 39778 15056 39790 15348
rect 39824 15056 39836 15348
rect 39778 14702 39836 15056
rect 40978 15348 41036 15702
rect 40978 15056 40990 15348
rect 41024 15056 41036 15348
rect 40978 14702 41036 15056
rect 42036 15348 42094 15702
rect 42036 15056 42048 15348
rect 42082 15056 42094 15348
rect 42036 14702 42094 15056
rect 43094 15348 43152 15702
rect 43094 15056 43106 15348
rect 43140 15056 43152 15348
rect 43094 14702 43152 15056
rect 44152 15348 44210 15702
rect 44152 15056 44164 15348
rect 44198 15056 44210 15348
rect 44152 14702 44210 15056
rect 45210 15348 45268 15702
rect 45210 15056 45222 15348
rect 45256 15056 45268 15348
rect 45210 14702 45268 15056
rect 46268 15348 46326 15702
rect 46268 15056 46280 15348
rect 46314 15056 46326 15348
rect 46268 14702 46326 15056
rect 47566 15370 47624 15724
rect 47566 15078 47578 15370
rect 47612 15078 47624 15370
rect 47566 14724 47624 15078
rect 48624 15370 48682 15724
rect 48624 15078 48636 15370
rect 48670 15078 48682 15370
rect 48624 14724 48682 15078
rect 49682 15370 49740 15724
rect 49682 15078 49694 15370
rect 49728 15078 49740 15370
rect 49682 14724 49740 15078
rect 50740 15370 50798 15724
rect 50740 15078 50752 15370
rect 50786 15078 50798 15370
rect 50740 14724 50798 15078
rect 51798 15370 51856 15724
rect 51798 15078 51810 15370
rect 51844 15078 51856 15370
rect 51798 14724 51856 15078
rect 52856 15370 52914 15724
rect 52856 15078 52868 15370
rect 52902 15078 52914 15370
rect 52856 14724 52914 15078
rect 54080 15384 54138 15738
rect 54080 15092 54092 15384
rect 54126 15092 54138 15384
rect 54080 14738 54138 15092
rect 55138 15384 55196 15738
rect 55138 15092 55150 15384
rect 55184 15092 55196 15384
rect 55138 14738 55196 15092
rect 56196 15384 56254 15738
rect 56196 15092 56208 15384
rect 56242 15092 56254 15384
rect 56196 14738 56254 15092
rect 57254 15384 57312 15738
rect 57254 15092 57266 15384
rect 57300 15092 57312 15384
rect 57254 14738 57312 15092
rect 58312 15384 58370 15738
rect 58312 15092 58324 15384
rect 58358 15092 58370 15384
rect 58312 14738 58370 15092
rect 59370 15384 59428 15738
rect 59370 15092 59382 15384
rect 59416 15092 59428 15384
rect 59370 14738 59428 15092
rect 1956 13846 2014 14200
rect 1956 13554 1968 13846
rect 2002 13554 2014 13846
rect 1956 13200 2014 13554
rect 3014 13846 3072 14200
rect 3014 13554 3026 13846
rect 3060 13554 3072 13846
rect 3014 13200 3072 13554
rect 4072 13846 4130 14200
rect 4072 13554 4084 13846
rect 4118 13554 4130 13846
rect 4072 13200 4130 13554
rect 5130 13846 5188 14200
rect 5130 13554 5142 13846
rect 5176 13554 5188 13846
rect 5130 13200 5188 13554
rect 6188 13846 6246 14200
rect 6188 13554 6200 13846
rect 6234 13554 6246 13846
rect 6188 13200 6246 13554
rect 7246 13846 7304 14200
rect 7246 13554 7258 13846
rect 7292 13554 7304 13846
rect 7246 13200 7304 13554
rect 8470 13854 8528 14208
rect 8470 13562 8482 13854
rect 8516 13562 8528 13854
rect 8470 13208 8528 13562
rect 9528 13854 9586 14208
rect 9528 13562 9540 13854
rect 9574 13562 9586 13854
rect 9528 13208 9586 13562
rect 10586 13854 10644 14208
rect 10586 13562 10598 13854
rect 10632 13562 10644 13854
rect 10586 13208 10644 13562
rect 11644 13854 11702 14208
rect 11644 13562 11656 13854
rect 11690 13562 11702 13854
rect 11644 13208 11702 13562
rect 12702 13854 12760 14208
rect 12702 13562 12714 13854
rect 12748 13562 12760 13854
rect 12702 13208 12760 13562
rect 13760 13854 13818 14208
rect 13760 13562 13772 13854
rect 13806 13562 13818 13854
rect 13760 13208 13818 13562
rect 14976 13862 15034 14216
rect 14976 13570 14988 13862
rect 15022 13570 15034 13862
rect 14976 13216 15034 13570
rect 16034 13862 16092 14216
rect 16034 13570 16046 13862
rect 16080 13570 16092 13862
rect 16034 13216 16092 13570
rect 17092 13862 17150 14216
rect 17092 13570 17104 13862
rect 17138 13570 17150 13862
rect 17092 13216 17150 13570
rect 18150 13862 18208 14216
rect 18150 13570 18162 13862
rect 18196 13570 18208 13862
rect 18150 13216 18208 13570
rect 19208 13862 19266 14216
rect 19208 13570 19220 13862
rect 19254 13570 19266 13862
rect 19208 13216 19266 13570
rect 20266 13862 20324 14216
rect 20266 13570 20278 13862
rect 20312 13570 20324 13862
rect 20266 13216 20324 13570
rect 21466 13846 21524 14200
rect 21466 13554 21478 13846
rect 21512 13554 21524 13846
rect 21466 13200 21524 13554
rect 22524 13846 22582 14200
rect 22524 13554 22536 13846
rect 22570 13554 22582 13846
rect 22524 13200 22582 13554
rect 23582 13846 23640 14200
rect 23582 13554 23594 13846
rect 23628 13554 23640 13846
rect 23582 13200 23640 13554
rect 24640 13846 24698 14200
rect 24640 13554 24652 13846
rect 24686 13554 24698 13846
rect 24640 13200 24698 13554
rect 25698 13846 25756 14200
rect 25698 13554 25710 13846
rect 25744 13554 25756 13846
rect 25698 13200 25756 13554
rect 26756 13846 26814 14200
rect 26756 13554 26768 13846
rect 26802 13554 26814 13846
rect 26756 13200 26814 13554
rect 27988 13862 28046 14216
rect 27988 13570 28000 13862
rect 28034 13570 28046 13862
rect 27988 13216 28046 13570
rect 29046 13862 29104 14216
rect 29046 13570 29058 13862
rect 29092 13570 29104 13862
rect 29046 13216 29104 13570
rect 30104 13862 30162 14216
rect 30104 13570 30116 13862
rect 30150 13570 30162 13862
rect 30104 13216 30162 13570
rect 31162 13862 31220 14216
rect 31162 13570 31174 13862
rect 31208 13570 31220 13862
rect 31162 13216 31220 13570
rect 32220 13862 32278 14216
rect 32220 13570 32232 13862
rect 32266 13570 32278 13862
rect 32220 13216 32278 13570
rect 33278 13862 33336 14216
rect 33278 13570 33290 13862
rect 33324 13570 33336 13862
rect 33278 13216 33336 13570
rect 34498 13868 34556 14222
rect 34498 13576 34510 13868
rect 34544 13576 34556 13868
rect 34498 13222 34556 13576
rect 35556 13868 35614 14222
rect 35556 13576 35568 13868
rect 35602 13576 35614 13868
rect 35556 13222 35614 13576
rect 36614 13868 36672 14222
rect 36614 13576 36626 13868
rect 36660 13576 36672 13868
rect 36614 13222 36672 13576
rect 37672 13868 37730 14222
rect 37672 13576 37684 13868
rect 37718 13576 37730 13868
rect 37672 13222 37730 13576
rect 38730 13868 38788 14222
rect 38730 13576 38742 13868
rect 38776 13576 38788 13868
rect 38730 13222 38788 13576
rect 39788 13868 39846 14222
rect 39788 13576 39800 13868
rect 39834 13576 39846 13868
rect 39788 13222 39846 13576
rect 40988 13868 41046 14222
rect 40988 13576 41000 13868
rect 41034 13576 41046 13868
rect 40988 13222 41046 13576
rect 42046 13868 42104 14222
rect 42046 13576 42058 13868
rect 42092 13576 42104 13868
rect 42046 13222 42104 13576
rect 43104 13868 43162 14222
rect 43104 13576 43116 13868
rect 43150 13576 43162 13868
rect 43104 13222 43162 13576
rect 44162 13868 44220 14222
rect 44162 13576 44174 13868
rect 44208 13576 44220 13868
rect 44162 13222 44220 13576
rect 45220 13868 45278 14222
rect 45220 13576 45232 13868
rect 45266 13576 45278 13868
rect 45220 13222 45278 13576
rect 46278 13868 46336 14222
rect 46278 13576 46290 13868
rect 46324 13576 46336 13868
rect 46278 13222 46336 13576
rect 47576 13890 47634 14244
rect 47576 13598 47588 13890
rect 47622 13598 47634 13890
rect 47576 13244 47634 13598
rect 48634 13890 48692 14244
rect 48634 13598 48646 13890
rect 48680 13598 48692 13890
rect 48634 13244 48692 13598
rect 49692 13890 49750 14244
rect 49692 13598 49704 13890
rect 49738 13598 49750 13890
rect 49692 13244 49750 13598
rect 50750 13890 50808 14244
rect 50750 13598 50762 13890
rect 50796 13598 50808 13890
rect 50750 13244 50808 13598
rect 51808 13890 51866 14244
rect 51808 13598 51820 13890
rect 51854 13598 51866 13890
rect 51808 13244 51866 13598
rect 52866 13890 52924 14244
rect 52866 13598 52878 13890
rect 52912 13598 52924 13890
rect 52866 13244 52924 13598
rect 54090 13904 54148 14258
rect 54090 13612 54102 13904
rect 54136 13612 54148 13904
rect 54090 13258 54148 13612
rect 55148 13904 55206 14258
rect 55148 13612 55160 13904
rect 55194 13612 55206 13904
rect 55148 13258 55206 13612
rect 56206 13904 56264 14258
rect 56206 13612 56218 13904
rect 56252 13612 56264 13904
rect 56206 13258 56264 13612
rect 57264 13904 57322 14258
rect 57264 13612 57276 13904
rect 57310 13612 57322 13904
rect 57264 13258 57322 13612
rect 58322 13904 58380 14258
rect 58322 13612 58334 13904
rect 58368 13612 58380 13904
rect 58322 13258 58380 13612
rect 59380 13904 59438 14258
rect 59380 13612 59392 13904
rect 59426 13612 59438 13904
rect 59380 13258 59438 13612
rect 1956 12752 2014 13106
rect 1956 12460 1968 12752
rect 2002 12460 2014 12752
rect 1956 12106 2014 12460
rect 3014 12752 3072 13106
rect 3014 12460 3026 12752
rect 3060 12460 3072 12752
rect 3014 12106 3072 12460
rect 4072 12752 4130 13106
rect 4072 12460 4084 12752
rect 4118 12460 4130 12752
rect 4072 12106 4130 12460
rect 5130 12752 5188 13106
rect 5130 12460 5142 12752
rect 5176 12460 5188 12752
rect 5130 12106 5188 12460
rect 6188 12752 6246 13106
rect 6188 12460 6200 12752
rect 6234 12460 6246 12752
rect 6188 12106 6246 12460
rect 7246 12752 7304 13106
rect 7246 12460 7258 12752
rect 7292 12460 7304 12752
rect 8470 12760 8528 13114
rect 7246 12106 7304 12460
rect 1956 11658 2014 12012
rect 1956 11366 1968 11658
rect 2002 11366 2014 11658
rect 1956 11012 2014 11366
rect 3014 11658 3072 12012
rect 3014 11366 3026 11658
rect 3060 11366 3072 11658
rect 3014 11012 3072 11366
rect 4072 11658 4130 12012
rect 4072 11366 4084 11658
rect 4118 11366 4130 11658
rect 4072 11012 4130 11366
rect 5130 11658 5188 12012
rect 5130 11366 5142 11658
rect 5176 11366 5188 11658
rect 5130 11012 5188 11366
rect 6188 11658 6246 12012
rect 6188 11366 6200 11658
rect 6234 11366 6246 11658
rect 6188 11012 6246 11366
rect 7246 11658 7304 12012
rect 7246 11366 7258 11658
rect 7292 11366 7304 11658
rect 7246 11012 7304 11366
rect 8470 12468 8482 12760
rect 8516 12468 8528 12760
rect 8470 12114 8528 12468
rect 9528 12760 9586 13114
rect 9528 12468 9540 12760
rect 9574 12468 9586 12760
rect 9528 12114 9586 12468
rect 10586 12760 10644 13114
rect 10586 12468 10598 12760
rect 10632 12468 10644 12760
rect 10586 12114 10644 12468
rect 11644 12760 11702 13114
rect 11644 12468 11656 12760
rect 11690 12468 11702 12760
rect 11644 12114 11702 12468
rect 12702 12760 12760 13114
rect 12702 12468 12714 12760
rect 12748 12468 12760 12760
rect 12702 12114 12760 12468
rect 13760 12760 13818 13114
rect 13760 12468 13772 12760
rect 13806 12468 13818 12760
rect 14976 12768 15034 13122
rect 13760 12114 13818 12468
rect 1956 10564 2014 10918
rect 1956 10272 1968 10564
rect 2002 10272 2014 10564
rect 1956 9918 2014 10272
rect 3014 10564 3072 10918
rect 3014 10272 3026 10564
rect 3060 10272 3072 10564
rect 3014 9918 3072 10272
rect 4072 10564 4130 10918
rect 4072 10272 4084 10564
rect 4118 10272 4130 10564
rect 4072 9918 4130 10272
rect 5130 10564 5188 10918
rect 5130 10272 5142 10564
rect 5176 10272 5188 10564
rect 5130 9918 5188 10272
rect 6188 10564 6246 10918
rect 6188 10272 6200 10564
rect 6234 10272 6246 10564
rect 6188 9918 6246 10272
rect 7246 10564 7304 10918
rect 8470 11666 8528 12020
rect 8470 11374 8482 11666
rect 8516 11374 8528 11666
rect 8470 11020 8528 11374
rect 9528 11666 9586 12020
rect 9528 11374 9540 11666
rect 9574 11374 9586 11666
rect 9528 11020 9586 11374
rect 10586 11666 10644 12020
rect 10586 11374 10598 11666
rect 10632 11374 10644 11666
rect 10586 11020 10644 11374
rect 11644 11666 11702 12020
rect 11644 11374 11656 11666
rect 11690 11374 11702 11666
rect 11644 11020 11702 11374
rect 12702 11666 12760 12020
rect 12702 11374 12714 11666
rect 12748 11374 12760 11666
rect 12702 11020 12760 11374
rect 13760 11666 13818 12020
rect 13760 11374 13772 11666
rect 13806 11374 13818 11666
rect 13760 11020 13818 11374
rect 14976 12476 14988 12768
rect 15022 12476 15034 12768
rect 14976 12122 15034 12476
rect 16034 12768 16092 13122
rect 16034 12476 16046 12768
rect 16080 12476 16092 12768
rect 16034 12122 16092 12476
rect 17092 12768 17150 13122
rect 17092 12476 17104 12768
rect 17138 12476 17150 12768
rect 17092 12122 17150 12476
rect 18150 12768 18208 13122
rect 18150 12476 18162 12768
rect 18196 12476 18208 12768
rect 18150 12122 18208 12476
rect 19208 12768 19266 13122
rect 19208 12476 19220 12768
rect 19254 12476 19266 12768
rect 19208 12122 19266 12476
rect 20266 12768 20324 13122
rect 20266 12476 20278 12768
rect 20312 12476 20324 12768
rect 20266 12122 20324 12476
rect 21466 12752 21524 13106
rect 7246 10272 7258 10564
rect 7292 10272 7304 10564
rect 7246 9918 7304 10272
rect 8470 10572 8528 10926
rect 8470 10280 8482 10572
rect 8516 10280 8528 10572
rect 8470 9926 8528 10280
rect 9528 10572 9586 10926
rect 9528 10280 9540 10572
rect 9574 10280 9586 10572
rect 9528 9926 9586 10280
rect 10586 10572 10644 10926
rect 10586 10280 10598 10572
rect 10632 10280 10644 10572
rect 10586 9926 10644 10280
rect 11644 10572 11702 10926
rect 11644 10280 11656 10572
rect 11690 10280 11702 10572
rect 11644 9926 11702 10280
rect 12702 10572 12760 10926
rect 12702 10280 12714 10572
rect 12748 10280 12760 10572
rect 12702 9926 12760 10280
rect 13760 10572 13818 10926
rect 14976 11674 15034 12028
rect 14976 11382 14988 11674
rect 15022 11382 15034 11674
rect 14976 11028 15034 11382
rect 16034 11674 16092 12028
rect 16034 11382 16046 11674
rect 16080 11382 16092 11674
rect 16034 11028 16092 11382
rect 17092 11674 17150 12028
rect 17092 11382 17104 11674
rect 17138 11382 17150 11674
rect 17092 11028 17150 11382
rect 18150 11674 18208 12028
rect 18150 11382 18162 11674
rect 18196 11382 18208 11674
rect 18150 11028 18208 11382
rect 19208 11674 19266 12028
rect 19208 11382 19220 11674
rect 19254 11382 19266 11674
rect 19208 11028 19266 11382
rect 20266 11674 20324 12028
rect 20266 11382 20278 11674
rect 20312 11382 20324 11674
rect 20266 11028 20324 11382
rect 21466 12460 21478 12752
rect 21512 12460 21524 12752
rect 21466 12106 21524 12460
rect 22524 12752 22582 13106
rect 22524 12460 22536 12752
rect 22570 12460 22582 12752
rect 22524 12106 22582 12460
rect 23582 12752 23640 13106
rect 23582 12460 23594 12752
rect 23628 12460 23640 12752
rect 23582 12106 23640 12460
rect 24640 12752 24698 13106
rect 24640 12460 24652 12752
rect 24686 12460 24698 12752
rect 24640 12106 24698 12460
rect 25698 12752 25756 13106
rect 25698 12460 25710 12752
rect 25744 12460 25756 12752
rect 25698 12106 25756 12460
rect 26756 12752 26814 13106
rect 26756 12460 26768 12752
rect 26802 12460 26814 12752
rect 27988 12768 28046 13122
rect 26756 12106 26814 12460
rect 13760 10280 13772 10572
rect 13806 10280 13818 10572
rect 13760 9926 13818 10280
rect 14976 10580 15034 10934
rect 14976 10288 14988 10580
rect 15022 10288 15034 10580
rect 14976 9934 15034 10288
rect 16034 10580 16092 10934
rect 16034 10288 16046 10580
rect 16080 10288 16092 10580
rect 16034 9934 16092 10288
rect 17092 10580 17150 10934
rect 17092 10288 17104 10580
rect 17138 10288 17150 10580
rect 17092 9934 17150 10288
rect 18150 10580 18208 10934
rect 18150 10288 18162 10580
rect 18196 10288 18208 10580
rect 18150 9934 18208 10288
rect 19208 10580 19266 10934
rect 19208 10288 19220 10580
rect 19254 10288 19266 10580
rect 19208 9934 19266 10288
rect 20266 10580 20324 10934
rect 21466 11658 21524 12012
rect 21466 11366 21478 11658
rect 21512 11366 21524 11658
rect 21466 11012 21524 11366
rect 22524 11658 22582 12012
rect 22524 11366 22536 11658
rect 22570 11366 22582 11658
rect 22524 11012 22582 11366
rect 23582 11658 23640 12012
rect 23582 11366 23594 11658
rect 23628 11366 23640 11658
rect 23582 11012 23640 11366
rect 24640 11658 24698 12012
rect 24640 11366 24652 11658
rect 24686 11366 24698 11658
rect 24640 11012 24698 11366
rect 25698 11658 25756 12012
rect 25698 11366 25710 11658
rect 25744 11366 25756 11658
rect 25698 11012 25756 11366
rect 26756 11658 26814 12012
rect 26756 11366 26768 11658
rect 26802 11366 26814 11658
rect 26756 11012 26814 11366
rect 27988 12476 28000 12768
rect 28034 12476 28046 12768
rect 27988 12122 28046 12476
rect 29046 12768 29104 13122
rect 29046 12476 29058 12768
rect 29092 12476 29104 12768
rect 29046 12122 29104 12476
rect 30104 12768 30162 13122
rect 30104 12476 30116 12768
rect 30150 12476 30162 12768
rect 30104 12122 30162 12476
rect 31162 12768 31220 13122
rect 31162 12476 31174 12768
rect 31208 12476 31220 12768
rect 31162 12122 31220 12476
rect 32220 12768 32278 13122
rect 32220 12476 32232 12768
rect 32266 12476 32278 12768
rect 32220 12122 32278 12476
rect 33278 12768 33336 13122
rect 33278 12476 33290 12768
rect 33324 12476 33336 12768
rect 34498 12774 34556 13128
rect 33278 12122 33336 12476
rect 20266 10288 20278 10580
rect 20312 10288 20324 10580
rect 20266 9934 20324 10288
rect 21466 10564 21524 10918
rect 21466 10272 21478 10564
rect 21512 10272 21524 10564
rect 21466 9918 21524 10272
rect 22524 10564 22582 10918
rect 22524 10272 22536 10564
rect 22570 10272 22582 10564
rect 22524 9918 22582 10272
rect 23582 10564 23640 10918
rect 23582 10272 23594 10564
rect 23628 10272 23640 10564
rect 23582 9918 23640 10272
rect 24640 10564 24698 10918
rect 24640 10272 24652 10564
rect 24686 10272 24698 10564
rect 24640 9918 24698 10272
rect 25698 10564 25756 10918
rect 25698 10272 25710 10564
rect 25744 10272 25756 10564
rect 25698 9918 25756 10272
rect 26756 10564 26814 10918
rect 27988 11674 28046 12028
rect 27988 11382 28000 11674
rect 28034 11382 28046 11674
rect 27988 11028 28046 11382
rect 29046 11674 29104 12028
rect 29046 11382 29058 11674
rect 29092 11382 29104 11674
rect 29046 11028 29104 11382
rect 30104 11674 30162 12028
rect 30104 11382 30116 11674
rect 30150 11382 30162 11674
rect 30104 11028 30162 11382
rect 31162 11674 31220 12028
rect 31162 11382 31174 11674
rect 31208 11382 31220 11674
rect 31162 11028 31220 11382
rect 32220 11674 32278 12028
rect 32220 11382 32232 11674
rect 32266 11382 32278 11674
rect 32220 11028 32278 11382
rect 33278 11674 33336 12028
rect 33278 11382 33290 11674
rect 33324 11382 33336 11674
rect 33278 11028 33336 11382
rect 34498 12482 34510 12774
rect 34544 12482 34556 12774
rect 34498 12128 34556 12482
rect 35556 12774 35614 13128
rect 35556 12482 35568 12774
rect 35602 12482 35614 12774
rect 35556 12128 35614 12482
rect 36614 12774 36672 13128
rect 36614 12482 36626 12774
rect 36660 12482 36672 12774
rect 36614 12128 36672 12482
rect 37672 12774 37730 13128
rect 37672 12482 37684 12774
rect 37718 12482 37730 12774
rect 37672 12128 37730 12482
rect 38730 12774 38788 13128
rect 38730 12482 38742 12774
rect 38776 12482 38788 12774
rect 38730 12128 38788 12482
rect 39788 12774 39846 13128
rect 39788 12482 39800 12774
rect 39834 12482 39846 12774
rect 40988 12774 41046 13128
rect 39788 12128 39846 12482
rect 26756 10272 26768 10564
rect 26802 10272 26814 10564
rect 26756 9918 26814 10272
rect 27988 10580 28046 10934
rect 27988 10288 28000 10580
rect 28034 10288 28046 10580
rect 27988 9934 28046 10288
rect 29046 10580 29104 10934
rect 29046 10288 29058 10580
rect 29092 10288 29104 10580
rect 29046 9934 29104 10288
rect 30104 10580 30162 10934
rect 30104 10288 30116 10580
rect 30150 10288 30162 10580
rect 30104 9934 30162 10288
rect 31162 10580 31220 10934
rect 31162 10288 31174 10580
rect 31208 10288 31220 10580
rect 31162 9934 31220 10288
rect 32220 10580 32278 10934
rect 32220 10288 32232 10580
rect 32266 10288 32278 10580
rect 32220 9934 32278 10288
rect 33278 10580 33336 10934
rect 34498 11680 34556 12034
rect 34498 11388 34510 11680
rect 34544 11388 34556 11680
rect 34498 11034 34556 11388
rect 35556 11680 35614 12034
rect 35556 11388 35568 11680
rect 35602 11388 35614 11680
rect 35556 11034 35614 11388
rect 36614 11680 36672 12034
rect 36614 11388 36626 11680
rect 36660 11388 36672 11680
rect 36614 11034 36672 11388
rect 37672 11680 37730 12034
rect 37672 11388 37684 11680
rect 37718 11388 37730 11680
rect 37672 11034 37730 11388
rect 38730 11680 38788 12034
rect 38730 11388 38742 11680
rect 38776 11388 38788 11680
rect 38730 11034 38788 11388
rect 39788 11680 39846 12034
rect 39788 11388 39800 11680
rect 39834 11388 39846 11680
rect 39788 11034 39846 11388
rect 40988 12482 41000 12774
rect 41034 12482 41046 12774
rect 40988 12128 41046 12482
rect 42046 12774 42104 13128
rect 42046 12482 42058 12774
rect 42092 12482 42104 12774
rect 42046 12128 42104 12482
rect 43104 12774 43162 13128
rect 43104 12482 43116 12774
rect 43150 12482 43162 12774
rect 43104 12128 43162 12482
rect 44162 12774 44220 13128
rect 44162 12482 44174 12774
rect 44208 12482 44220 12774
rect 44162 12128 44220 12482
rect 45220 12774 45278 13128
rect 45220 12482 45232 12774
rect 45266 12482 45278 12774
rect 45220 12128 45278 12482
rect 46278 12774 46336 13128
rect 46278 12482 46290 12774
rect 46324 12482 46336 12774
rect 47576 12796 47634 13150
rect 46278 12128 46336 12482
rect 33278 10288 33290 10580
rect 33324 10288 33336 10580
rect 33278 9934 33336 10288
rect 34498 10586 34556 10940
rect 34498 10294 34510 10586
rect 34544 10294 34556 10586
rect 34498 9940 34556 10294
rect 35556 10586 35614 10940
rect 35556 10294 35568 10586
rect 35602 10294 35614 10586
rect 35556 9940 35614 10294
rect 36614 10586 36672 10940
rect 36614 10294 36626 10586
rect 36660 10294 36672 10586
rect 36614 9940 36672 10294
rect 37672 10586 37730 10940
rect 37672 10294 37684 10586
rect 37718 10294 37730 10586
rect 37672 9940 37730 10294
rect 38730 10586 38788 10940
rect 38730 10294 38742 10586
rect 38776 10294 38788 10586
rect 38730 9940 38788 10294
rect 39788 10586 39846 10940
rect 40988 11680 41046 12034
rect 40988 11388 41000 11680
rect 41034 11388 41046 11680
rect 40988 11034 41046 11388
rect 42046 11680 42104 12034
rect 42046 11388 42058 11680
rect 42092 11388 42104 11680
rect 42046 11034 42104 11388
rect 43104 11680 43162 12034
rect 43104 11388 43116 11680
rect 43150 11388 43162 11680
rect 43104 11034 43162 11388
rect 44162 11680 44220 12034
rect 44162 11388 44174 11680
rect 44208 11388 44220 11680
rect 44162 11034 44220 11388
rect 45220 11680 45278 12034
rect 45220 11388 45232 11680
rect 45266 11388 45278 11680
rect 45220 11034 45278 11388
rect 46278 11680 46336 12034
rect 46278 11388 46290 11680
rect 46324 11388 46336 11680
rect 46278 11034 46336 11388
rect 47576 12504 47588 12796
rect 47622 12504 47634 12796
rect 47576 12150 47634 12504
rect 48634 12796 48692 13150
rect 48634 12504 48646 12796
rect 48680 12504 48692 12796
rect 48634 12150 48692 12504
rect 49692 12796 49750 13150
rect 49692 12504 49704 12796
rect 49738 12504 49750 12796
rect 49692 12150 49750 12504
rect 50750 12796 50808 13150
rect 50750 12504 50762 12796
rect 50796 12504 50808 12796
rect 50750 12150 50808 12504
rect 51808 12796 51866 13150
rect 51808 12504 51820 12796
rect 51854 12504 51866 12796
rect 51808 12150 51866 12504
rect 52866 12796 52924 13150
rect 52866 12504 52878 12796
rect 52912 12504 52924 12796
rect 54090 12810 54148 13164
rect 52866 12150 52924 12504
rect 39788 10294 39800 10586
rect 39834 10294 39846 10586
rect 39788 9940 39846 10294
rect 40988 10586 41046 10940
rect 40988 10294 41000 10586
rect 41034 10294 41046 10586
rect 40988 9940 41046 10294
rect 42046 10586 42104 10940
rect 42046 10294 42058 10586
rect 42092 10294 42104 10586
rect 42046 9940 42104 10294
rect 43104 10586 43162 10940
rect 43104 10294 43116 10586
rect 43150 10294 43162 10586
rect 43104 9940 43162 10294
rect 44162 10586 44220 10940
rect 44162 10294 44174 10586
rect 44208 10294 44220 10586
rect 44162 9940 44220 10294
rect 45220 10586 45278 10940
rect 45220 10294 45232 10586
rect 45266 10294 45278 10586
rect 45220 9940 45278 10294
rect 46278 10586 46336 10940
rect 47576 11702 47634 12056
rect 47576 11410 47588 11702
rect 47622 11410 47634 11702
rect 47576 11056 47634 11410
rect 48634 11702 48692 12056
rect 48634 11410 48646 11702
rect 48680 11410 48692 11702
rect 48634 11056 48692 11410
rect 49692 11702 49750 12056
rect 49692 11410 49704 11702
rect 49738 11410 49750 11702
rect 49692 11056 49750 11410
rect 50750 11702 50808 12056
rect 50750 11410 50762 11702
rect 50796 11410 50808 11702
rect 50750 11056 50808 11410
rect 51808 11702 51866 12056
rect 51808 11410 51820 11702
rect 51854 11410 51866 11702
rect 51808 11056 51866 11410
rect 52866 11702 52924 12056
rect 52866 11410 52878 11702
rect 52912 11410 52924 11702
rect 52866 11056 52924 11410
rect 54090 12518 54102 12810
rect 54136 12518 54148 12810
rect 54090 12164 54148 12518
rect 55148 12810 55206 13164
rect 55148 12518 55160 12810
rect 55194 12518 55206 12810
rect 55148 12164 55206 12518
rect 56206 12810 56264 13164
rect 56206 12518 56218 12810
rect 56252 12518 56264 12810
rect 56206 12164 56264 12518
rect 57264 12810 57322 13164
rect 57264 12518 57276 12810
rect 57310 12518 57322 12810
rect 57264 12164 57322 12518
rect 58322 12810 58380 13164
rect 58322 12518 58334 12810
rect 58368 12518 58380 12810
rect 58322 12164 58380 12518
rect 59380 12810 59438 13164
rect 59380 12518 59392 12810
rect 59426 12518 59438 12810
rect 59380 12164 59438 12518
rect 46278 10294 46290 10586
rect 46324 10294 46336 10586
rect 46278 9940 46336 10294
rect 47576 10608 47634 10962
rect 47576 10316 47588 10608
rect 47622 10316 47634 10608
rect 47576 9962 47634 10316
rect 48634 10608 48692 10962
rect 48634 10316 48646 10608
rect 48680 10316 48692 10608
rect 48634 9962 48692 10316
rect 49692 10608 49750 10962
rect 49692 10316 49704 10608
rect 49738 10316 49750 10608
rect 49692 9962 49750 10316
rect 50750 10608 50808 10962
rect 50750 10316 50762 10608
rect 50796 10316 50808 10608
rect 50750 9962 50808 10316
rect 51808 10608 51866 10962
rect 51808 10316 51820 10608
rect 51854 10316 51866 10608
rect 51808 9962 51866 10316
rect 52866 10608 52924 10962
rect 54090 11716 54148 12070
rect 54090 11424 54102 11716
rect 54136 11424 54148 11716
rect 54090 11070 54148 11424
rect 55148 11716 55206 12070
rect 55148 11424 55160 11716
rect 55194 11424 55206 11716
rect 55148 11070 55206 11424
rect 56206 11716 56264 12070
rect 56206 11424 56218 11716
rect 56252 11424 56264 11716
rect 56206 11070 56264 11424
rect 57264 11716 57322 12070
rect 57264 11424 57276 11716
rect 57310 11424 57322 11716
rect 57264 11070 57322 11424
rect 58322 11716 58380 12070
rect 58322 11424 58334 11716
rect 58368 11424 58380 11716
rect 58322 11070 58380 11424
rect 59380 11716 59438 12070
rect 59380 11424 59392 11716
rect 59426 11424 59438 11716
rect 59380 11070 59438 11424
rect 52866 10316 52878 10608
rect 52912 10316 52924 10608
rect 52866 9962 52924 10316
rect 54090 10622 54148 10976
rect 54090 10330 54102 10622
rect 54136 10330 54148 10622
rect 54090 9976 54148 10330
rect 55148 10622 55206 10976
rect 55148 10330 55160 10622
rect 55194 10330 55206 10622
rect 55148 9976 55206 10330
rect 56206 10622 56264 10976
rect 56206 10330 56218 10622
rect 56252 10330 56264 10622
rect 56206 9976 56264 10330
rect 57264 10622 57322 10976
rect 57264 10330 57276 10622
rect 57310 10330 57322 10622
rect 57264 9976 57322 10330
rect 58322 10622 58380 10976
rect 58322 10330 58334 10622
rect 58368 10330 58380 10622
rect 58322 9976 58380 10330
rect 59380 10622 59438 10976
rect 59380 10330 59392 10622
rect 59426 10330 59438 10622
rect 59380 9976 59438 10330
rect 1956 9470 2014 9824
rect 1956 9178 1968 9470
rect 2002 9178 2014 9470
rect 1956 8824 2014 9178
rect 3014 9470 3072 9824
rect 3014 9178 3026 9470
rect 3060 9178 3072 9470
rect 3014 8824 3072 9178
rect 4072 9470 4130 9824
rect 4072 9178 4084 9470
rect 4118 9178 4130 9470
rect 4072 8824 4130 9178
rect 5130 9470 5188 9824
rect 5130 9178 5142 9470
rect 5176 9178 5188 9470
rect 5130 8824 5188 9178
rect 6188 9470 6246 9824
rect 6188 9178 6200 9470
rect 6234 9178 6246 9470
rect 6188 8824 6246 9178
rect 7246 9470 7304 9824
rect 7246 9178 7258 9470
rect 7292 9178 7304 9470
rect 7246 8824 7304 9178
rect 8470 9478 8528 9832
rect 8470 9186 8482 9478
rect 8516 9186 8528 9478
rect 8470 8832 8528 9186
rect 9528 9478 9586 9832
rect 9528 9186 9540 9478
rect 9574 9186 9586 9478
rect 9528 8832 9586 9186
rect 10586 9478 10644 9832
rect 10586 9186 10598 9478
rect 10632 9186 10644 9478
rect 10586 8832 10644 9186
rect 11644 9478 11702 9832
rect 11644 9186 11656 9478
rect 11690 9186 11702 9478
rect 11644 8832 11702 9186
rect 12702 9478 12760 9832
rect 12702 9186 12714 9478
rect 12748 9186 12760 9478
rect 12702 8832 12760 9186
rect 13760 9478 13818 9832
rect 13760 9186 13772 9478
rect 13806 9186 13818 9478
rect 13760 8832 13818 9186
rect 14976 9486 15034 9840
rect 14976 9194 14988 9486
rect 15022 9194 15034 9486
rect 14976 8840 15034 9194
rect 16034 9486 16092 9840
rect 16034 9194 16046 9486
rect 16080 9194 16092 9486
rect 16034 8840 16092 9194
rect 17092 9486 17150 9840
rect 17092 9194 17104 9486
rect 17138 9194 17150 9486
rect 17092 8840 17150 9194
rect 18150 9486 18208 9840
rect 18150 9194 18162 9486
rect 18196 9194 18208 9486
rect 18150 8840 18208 9194
rect 19208 9486 19266 9840
rect 19208 9194 19220 9486
rect 19254 9194 19266 9486
rect 19208 8840 19266 9194
rect 20266 9486 20324 9840
rect 20266 9194 20278 9486
rect 20312 9194 20324 9486
rect 20266 8840 20324 9194
rect 21466 9470 21524 9824
rect 21466 9178 21478 9470
rect 21512 9178 21524 9470
rect 21466 8824 21524 9178
rect 22524 9470 22582 9824
rect 22524 9178 22536 9470
rect 22570 9178 22582 9470
rect 22524 8824 22582 9178
rect 23582 9470 23640 9824
rect 23582 9178 23594 9470
rect 23628 9178 23640 9470
rect 23582 8824 23640 9178
rect 24640 9470 24698 9824
rect 24640 9178 24652 9470
rect 24686 9178 24698 9470
rect 24640 8824 24698 9178
rect 25698 9470 25756 9824
rect 25698 9178 25710 9470
rect 25744 9178 25756 9470
rect 25698 8824 25756 9178
rect 26756 9470 26814 9824
rect 26756 9178 26768 9470
rect 26802 9178 26814 9470
rect 26756 8824 26814 9178
rect 27988 9486 28046 9840
rect 27988 9194 28000 9486
rect 28034 9194 28046 9486
rect 27988 8840 28046 9194
rect 29046 9486 29104 9840
rect 29046 9194 29058 9486
rect 29092 9194 29104 9486
rect 29046 8840 29104 9194
rect 30104 9486 30162 9840
rect 30104 9194 30116 9486
rect 30150 9194 30162 9486
rect 30104 8840 30162 9194
rect 31162 9486 31220 9840
rect 31162 9194 31174 9486
rect 31208 9194 31220 9486
rect 31162 8840 31220 9194
rect 32220 9486 32278 9840
rect 32220 9194 32232 9486
rect 32266 9194 32278 9486
rect 32220 8840 32278 9194
rect 33278 9486 33336 9840
rect 33278 9194 33290 9486
rect 33324 9194 33336 9486
rect 33278 8840 33336 9194
rect 34498 9492 34556 9846
rect 34498 9200 34510 9492
rect 34544 9200 34556 9492
rect 34498 8846 34556 9200
rect 35556 9492 35614 9846
rect 35556 9200 35568 9492
rect 35602 9200 35614 9492
rect 35556 8846 35614 9200
rect 36614 9492 36672 9846
rect 36614 9200 36626 9492
rect 36660 9200 36672 9492
rect 36614 8846 36672 9200
rect 37672 9492 37730 9846
rect 37672 9200 37684 9492
rect 37718 9200 37730 9492
rect 37672 8846 37730 9200
rect 38730 9492 38788 9846
rect 38730 9200 38742 9492
rect 38776 9200 38788 9492
rect 38730 8846 38788 9200
rect 39788 9492 39846 9846
rect 39788 9200 39800 9492
rect 39834 9200 39846 9492
rect 39788 8846 39846 9200
rect 40988 9492 41046 9846
rect 40988 9200 41000 9492
rect 41034 9200 41046 9492
rect 40988 8846 41046 9200
rect 42046 9492 42104 9846
rect 42046 9200 42058 9492
rect 42092 9200 42104 9492
rect 42046 8846 42104 9200
rect 43104 9492 43162 9846
rect 43104 9200 43116 9492
rect 43150 9200 43162 9492
rect 43104 8846 43162 9200
rect 44162 9492 44220 9846
rect 44162 9200 44174 9492
rect 44208 9200 44220 9492
rect 44162 8846 44220 9200
rect 45220 9492 45278 9846
rect 45220 9200 45232 9492
rect 45266 9200 45278 9492
rect 45220 8846 45278 9200
rect 46278 9492 46336 9846
rect 46278 9200 46290 9492
rect 46324 9200 46336 9492
rect 46278 8846 46336 9200
rect 47576 9514 47634 9868
rect 47576 9222 47588 9514
rect 47622 9222 47634 9514
rect 47576 8868 47634 9222
rect 48634 9514 48692 9868
rect 48634 9222 48646 9514
rect 48680 9222 48692 9514
rect 48634 8868 48692 9222
rect 49692 9514 49750 9868
rect 49692 9222 49704 9514
rect 49738 9222 49750 9514
rect 49692 8868 49750 9222
rect 50750 9514 50808 9868
rect 50750 9222 50762 9514
rect 50796 9222 50808 9514
rect 50750 8868 50808 9222
rect 51808 9514 51866 9868
rect 51808 9222 51820 9514
rect 51854 9222 51866 9514
rect 51808 8868 51866 9222
rect 52866 9514 52924 9868
rect 52866 9222 52878 9514
rect 52912 9222 52924 9514
rect 52866 8868 52924 9222
rect 54090 9528 54148 9882
rect 54090 9236 54102 9528
rect 54136 9236 54148 9528
rect 54090 8882 54148 9236
rect 55148 9528 55206 9882
rect 55148 9236 55160 9528
rect 55194 9236 55206 9528
rect 55148 8882 55206 9236
rect 56206 9528 56264 9882
rect 56206 9236 56218 9528
rect 56252 9236 56264 9528
rect 56206 8882 56264 9236
rect 57264 9528 57322 9882
rect 57264 9236 57276 9528
rect 57310 9236 57322 9528
rect 57264 8882 57322 9236
rect 58322 9528 58380 9882
rect 58322 9236 58334 9528
rect 58368 9236 58380 9528
rect 58322 8882 58380 9236
rect 59380 9528 59438 9882
rect 59380 9236 59392 9528
rect 59426 9236 59438 9528
rect 59380 8882 59438 9236
rect 1974 7938 2032 8292
rect 1974 7646 1986 7938
rect 2020 7646 2032 7938
rect 1974 7292 2032 7646
rect 3032 7938 3090 8292
rect 3032 7646 3044 7938
rect 3078 7646 3090 7938
rect 3032 7292 3090 7646
rect 4090 7938 4148 8292
rect 4090 7646 4102 7938
rect 4136 7646 4148 7938
rect 4090 7292 4148 7646
rect 5148 7938 5206 8292
rect 5148 7646 5160 7938
rect 5194 7646 5206 7938
rect 5148 7292 5206 7646
rect 6206 7938 6264 8292
rect 6206 7646 6218 7938
rect 6252 7646 6264 7938
rect 6206 7292 6264 7646
rect 7264 7938 7322 8292
rect 7264 7646 7276 7938
rect 7310 7646 7322 7938
rect 7264 7292 7322 7646
rect 8488 7946 8546 8300
rect 8488 7654 8500 7946
rect 8534 7654 8546 7946
rect 8488 7300 8546 7654
rect 9546 7946 9604 8300
rect 9546 7654 9558 7946
rect 9592 7654 9604 7946
rect 9546 7300 9604 7654
rect 10604 7946 10662 8300
rect 10604 7654 10616 7946
rect 10650 7654 10662 7946
rect 10604 7300 10662 7654
rect 11662 7946 11720 8300
rect 11662 7654 11674 7946
rect 11708 7654 11720 7946
rect 11662 7300 11720 7654
rect 12720 7946 12778 8300
rect 12720 7654 12732 7946
rect 12766 7654 12778 7946
rect 12720 7300 12778 7654
rect 13778 7946 13836 8300
rect 13778 7654 13790 7946
rect 13824 7654 13836 7946
rect 13778 7300 13836 7654
rect 14994 7954 15052 8308
rect 14994 7662 15006 7954
rect 15040 7662 15052 7954
rect 14994 7308 15052 7662
rect 16052 7954 16110 8308
rect 16052 7662 16064 7954
rect 16098 7662 16110 7954
rect 16052 7308 16110 7662
rect 17110 7954 17168 8308
rect 17110 7662 17122 7954
rect 17156 7662 17168 7954
rect 17110 7308 17168 7662
rect 18168 7954 18226 8308
rect 18168 7662 18180 7954
rect 18214 7662 18226 7954
rect 18168 7308 18226 7662
rect 19226 7954 19284 8308
rect 19226 7662 19238 7954
rect 19272 7662 19284 7954
rect 19226 7308 19284 7662
rect 20284 7954 20342 8308
rect 20284 7662 20296 7954
rect 20330 7662 20342 7954
rect 20284 7308 20342 7662
rect 21484 7938 21542 8292
rect 21484 7646 21496 7938
rect 21530 7646 21542 7938
rect 21484 7292 21542 7646
rect 22542 7938 22600 8292
rect 22542 7646 22554 7938
rect 22588 7646 22600 7938
rect 22542 7292 22600 7646
rect 23600 7938 23658 8292
rect 23600 7646 23612 7938
rect 23646 7646 23658 7938
rect 23600 7292 23658 7646
rect 24658 7938 24716 8292
rect 24658 7646 24670 7938
rect 24704 7646 24716 7938
rect 24658 7292 24716 7646
rect 25716 7938 25774 8292
rect 25716 7646 25728 7938
rect 25762 7646 25774 7938
rect 25716 7292 25774 7646
rect 26774 7938 26832 8292
rect 26774 7646 26786 7938
rect 26820 7646 26832 7938
rect 26774 7292 26832 7646
rect 28006 7954 28064 8308
rect 28006 7662 28018 7954
rect 28052 7662 28064 7954
rect 28006 7308 28064 7662
rect 29064 7954 29122 8308
rect 29064 7662 29076 7954
rect 29110 7662 29122 7954
rect 29064 7308 29122 7662
rect 30122 7954 30180 8308
rect 30122 7662 30134 7954
rect 30168 7662 30180 7954
rect 30122 7308 30180 7662
rect 31180 7954 31238 8308
rect 31180 7662 31192 7954
rect 31226 7662 31238 7954
rect 31180 7308 31238 7662
rect 32238 7954 32296 8308
rect 32238 7662 32250 7954
rect 32284 7662 32296 7954
rect 32238 7308 32296 7662
rect 33296 7954 33354 8308
rect 33296 7662 33308 7954
rect 33342 7662 33354 7954
rect 33296 7308 33354 7662
rect 34516 7960 34574 8314
rect 34516 7668 34528 7960
rect 34562 7668 34574 7960
rect 34516 7314 34574 7668
rect 35574 7960 35632 8314
rect 35574 7668 35586 7960
rect 35620 7668 35632 7960
rect 35574 7314 35632 7668
rect 36632 7960 36690 8314
rect 36632 7668 36644 7960
rect 36678 7668 36690 7960
rect 36632 7314 36690 7668
rect 37690 7960 37748 8314
rect 37690 7668 37702 7960
rect 37736 7668 37748 7960
rect 37690 7314 37748 7668
rect 38748 7960 38806 8314
rect 38748 7668 38760 7960
rect 38794 7668 38806 7960
rect 38748 7314 38806 7668
rect 39806 7960 39864 8314
rect 39806 7668 39818 7960
rect 39852 7668 39864 7960
rect 39806 7314 39864 7668
rect 41006 7960 41064 8314
rect 41006 7668 41018 7960
rect 41052 7668 41064 7960
rect 41006 7314 41064 7668
rect 42064 7960 42122 8314
rect 42064 7668 42076 7960
rect 42110 7668 42122 7960
rect 42064 7314 42122 7668
rect 43122 7960 43180 8314
rect 43122 7668 43134 7960
rect 43168 7668 43180 7960
rect 43122 7314 43180 7668
rect 44180 7960 44238 8314
rect 44180 7668 44192 7960
rect 44226 7668 44238 7960
rect 44180 7314 44238 7668
rect 45238 7960 45296 8314
rect 45238 7668 45250 7960
rect 45284 7668 45296 7960
rect 45238 7314 45296 7668
rect 46296 7960 46354 8314
rect 46296 7668 46308 7960
rect 46342 7668 46354 7960
rect 46296 7314 46354 7668
rect 47594 7982 47652 8336
rect 47594 7690 47606 7982
rect 47640 7690 47652 7982
rect 47594 7336 47652 7690
rect 48652 7982 48710 8336
rect 48652 7690 48664 7982
rect 48698 7690 48710 7982
rect 48652 7336 48710 7690
rect 49710 7982 49768 8336
rect 49710 7690 49722 7982
rect 49756 7690 49768 7982
rect 49710 7336 49768 7690
rect 50768 7982 50826 8336
rect 50768 7690 50780 7982
rect 50814 7690 50826 7982
rect 50768 7336 50826 7690
rect 51826 7982 51884 8336
rect 51826 7690 51838 7982
rect 51872 7690 51884 7982
rect 51826 7336 51884 7690
rect 52884 7982 52942 8336
rect 52884 7690 52896 7982
rect 52930 7690 52942 7982
rect 52884 7336 52942 7690
rect 54108 7996 54166 8350
rect 54108 7704 54120 7996
rect 54154 7704 54166 7996
rect 54108 7350 54166 7704
rect 55166 7996 55224 8350
rect 55166 7704 55178 7996
rect 55212 7704 55224 7996
rect 55166 7350 55224 7704
rect 56224 7996 56282 8350
rect 56224 7704 56236 7996
rect 56270 7704 56282 7996
rect 56224 7350 56282 7704
rect 57282 7996 57340 8350
rect 57282 7704 57294 7996
rect 57328 7704 57340 7996
rect 57282 7350 57340 7704
rect 58340 7996 58398 8350
rect 58340 7704 58352 7996
rect 58386 7704 58398 7996
rect 58340 7350 58398 7704
rect 59398 7996 59456 8350
rect 59398 7704 59410 7996
rect 59444 7704 59456 7996
rect 59398 7350 59456 7704
rect 1974 6844 2032 7198
rect 1974 6552 1986 6844
rect 2020 6552 2032 6844
rect 1974 6198 2032 6552
rect 3032 6844 3090 7198
rect 3032 6552 3044 6844
rect 3078 6552 3090 6844
rect 3032 6198 3090 6552
rect 4090 6844 4148 7198
rect 4090 6552 4102 6844
rect 4136 6552 4148 6844
rect 4090 6198 4148 6552
rect 5148 6844 5206 7198
rect 5148 6552 5160 6844
rect 5194 6552 5206 6844
rect 5148 6198 5206 6552
rect 6206 6844 6264 7198
rect 6206 6552 6218 6844
rect 6252 6552 6264 6844
rect 6206 6198 6264 6552
rect 7264 6844 7322 7198
rect 7264 6552 7276 6844
rect 7310 6552 7322 6844
rect 8488 6852 8546 7206
rect 7264 6198 7322 6552
rect 1974 5750 2032 6104
rect 1974 5458 1986 5750
rect 2020 5458 2032 5750
rect 1974 5104 2032 5458
rect 3032 5750 3090 6104
rect 3032 5458 3044 5750
rect 3078 5458 3090 5750
rect 3032 5104 3090 5458
rect 4090 5750 4148 6104
rect 4090 5458 4102 5750
rect 4136 5458 4148 5750
rect 4090 5104 4148 5458
rect 5148 5750 5206 6104
rect 5148 5458 5160 5750
rect 5194 5458 5206 5750
rect 5148 5104 5206 5458
rect 6206 5750 6264 6104
rect 6206 5458 6218 5750
rect 6252 5458 6264 5750
rect 6206 5104 6264 5458
rect 7264 5750 7322 6104
rect 7264 5458 7276 5750
rect 7310 5458 7322 5750
rect 7264 5104 7322 5458
rect 8488 6560 8500 6852
rect 8534 6560 8546 6852
rect 8488 6206 8546 6560
rect 9546 6852 9604 7206
rect 9546 6560 9558 6852
rect 9592 6560 9604 6852
rect 9546 6206 9604 6560
rect 10604 6852 10662 7206
rect 10604 6560 10616 6852
rect 10650 6560 10662 6852
rect 10604 6206 10662 6560
rect 11662 6852 11720 7206
rect 11662 6560 11674 6852
rect 11708 6560 11720 6852
rect 11662 6206 11720 6560
rect 12720 6852 12778 7206
rect 12720 6560 12732 6852
rect 12766 6560 12778 6852
rect 12720 6206 12778 6560
rect 13778 6852 13836 7206
rect 13778 6560 13790 6852
rect 13824 6560 13836 6852
rect 14994 6860 15052 7214
rect 13778 6206 13836 6560
rect 1974 4656 2032 5010
rect 1974 4364 1986 4656
rect 2020 4364 2032 4656
rect 1974 4010 2032 4364
rect 3032 4656 3090 5010
rect 3032 4364 3044 4656
rect 3078 4364 3090 4656
rect 3032 4010 3090 4364
rect 4090 4656 4148 5010
rect 4090 4364 4102 4656
rect 4136 4364 4148 4656
rect 4090 4010 4148 4364
rect 5148 4656 5206 5010
rect 5148 4364 5160 4656
rect 5194 4364 5206 4656
rect 5148 4010 5206 4364
rect 6206 4656 6264 5010
rect 6206 4364 6218 4656
rect 6252 4364 6264 4656
rect 6206 4010 6264 4364
rect 7264 4656 7322 5010
rect 8488 5758 8546 6112
rect 8488 5466 8500 5758
rect 8534 5466 8546 5758
rect 8488 5112 8546 5466
rect 9546 5758 9604 6112
rect 9546 5466 9558 5758
rect 9592 5466 9604 5758
rect 9546 5112 9604 5466
rect 10604 5758 10662 6112
rect 10604 5466 10616 5758
rect 10650 5466 10662 5758
rect 10604 5112 10662 5466
rect 11662 5758 11720 6112
rect 11662 5466 11674 5758
rect 11708 5466 11720 5758
rect 11662 5112 11720 5466
rect 12720 5758 12778 6112
rect 12720 5466 12732 5758
rect 12766 5466 12778 5758
rect 12720 5112 12778 5466
rect 13778 5758 13836 6112
rect 13778 5466 13790 5758
rect 13824 5466 13836 5758
rect 13778 5112 13836 5466
rect 14994 6568 15006 6860
rect 15040 6568 15052 6860
rect 14994 6214 15052 6568
rect 16052 6860 16110 7214
rect 16052 6568 16064 6860
rect 16098 6568 16110 6860
rect 16052 6214 16110 6568
rect 17110 6860 17168 7214
rect 17110 6568 17122 6860
rect 17156 6568 17168 6860
rect 17110 6214 17168 6568
rect 18168 6860 18226 7214
rect 18168 6568 18180 6860
rect 18214 6568 18226 6860
rect 18168 6214 18226 6568
rect 19226 6860 19284 7214
rect 19226 6568 19238 6860
rect 19272 6568 19284 6860
rect 19226 6214 19284 6568
rect 20284 6860 20342 7214
rect 20284 6568 20296 6860
rect 20330 6568 20342 6860
rect 20284 6214 20342 6568
rect 21484 6844 21542 7198
rect 7264 4364 7276 4656
rect 7310 4364 7322 4656
rect 7264 4010 7322 4364
rect 8488 4664 8546 5018
rect 8488 4372 8500 4664
rect 8534 4372 8546 4664
rect 8488 4018 8546 4372
rect 9546 4664 9604 5018
rect 9546 4372 9558 4664
rect 9592 4372 9604 4664
rect 9546 4018 9604 4372
rect 10604 4664 10662 5018
rect 10604 4372 10616 4664
rect 10650 4372 10662 4664
rect 10604 4018 10662 4372
rect 11662 4664 11720 5018
rect 11662 4372 11674 4664
rect 11708 4372 11720 4664
rect 11662 4018 11720 4372
rect 12720 4664 12778 5018
rect 12720 4372 12732 4664
rect 12766 4372 12778 4664
rect 12720 4018 12778 4372
rect 13778 4664 13836 5018
rect 14994 5766 15052 6120
rect 14994 5474 15006 5766
rect 15040 5474 15052 5766
rect 14994 5120 15052 5474
rect 16052 5766 16110 6120
rect 16052 5474 16064 5766
rect 16098 5474 16110 5766
rect 16052 5120 16110 5474
rect 17110 5766 17168 6120
rect 17110 5474 17122 5766
rect 17156 5474 17168 5766
rect 17110 5120 17168 5474
rect 18168 5766 18226 6120
rect 18168 5474 18180 5766
rect 18214 5474 18226 5766
rect 18168 5120 18226 5474
rect 19226 5766 19284 6120
rect 19226 5474 19238 5766
rect 19272 5474 19284 5766
rect 19226 5120 19284 5474
rect 20284 5766 20342 6120
rect 20284 5474 20296 5766
rect 20330 5474 20342 5766
rect 20284 5120 20342 5474
rect 21484 6552 21496 6844
rect 21530 6552 21542 6844
rect 21484 6198 21542 6552
rect 22542 6844 22600 7198
rect 22542 6552 22554 6844
rect 22588 6552 22600 6844
rect 22542 6198 22600 6552
rect 23600 6844 23658 7198
rect 23600 6552 23612 6844
rect 23646 6552 23658 6844
rect 23600 6198 23658 6552
rect 24658 6844 24716 7198
rect 24658 6552 24670 6844
rect 24704 6552 24716 6844
rect 24658 6198 24716 6552
rect 25716 6844 25774 7198
rect 25716 6552 25728 6844
rect 25762 6552 25774 6844
rect 25716 6198 25774 6552
rect 26774 6844 26832 7198
rect 26774 6552 26786 6844
rect 26820 6552 26832 6844
rect 28006 6860 28064 7214
rect 26774 6198 26832 6552
rect 13778 4372 13790 4664
rect 13824 4372 13836 4664
rect 13778 4018 13836 4372
rect 14994 4672 15052 5026
rect 14994 4380 15006 4672
rect 15040 4380 15052 4672
rect 14994 4026 15052 4380
rect 16052 4672 16110 5026
rect 16052 4380 16064 4672
rect 16098 4380 16110 4672
rect 16052 4026 16110 4380
rect 17110 4672 17168 5026
rect 17110 4380 17122 4672
rect 17156 4380 17168 4672
rect 17110 4026 17168 4380
rect 18168 4672 18226 5026
rect 18168 4380 18180 4672
rect 18214 4380 18226 4672
rect 18168 4026 18226 4380
rect 19226 4672 19284 5026
rect 19226 4380 19238 4672
rect 19272 4380 19284 4672
rect 19226 4026 19284 4380
rect 20284 4672 20342 5026
rect 21484 5750 21542 6104
rect 21484 5458 21496 5750
rect 21530 5458 21542 5750
rect 21484 5104 21542 5458
rect 22542 5750 22600 6104
rect 22542 5458 22554 5750
rect 22588 5458 22600 5750
rect 22542 5104 22600 5458
rect 23600 5750 23658 6104
rect 23600 5458 23612 5750
rect 23646 5458 23658 5750
rect 23600 5104 23658 5458
rect 24658 5750 24716 6104
rect 24658 5458 24670 5750
rect 24704 5458 24716 5750
rect 24658 5104 24716 5458
rect 25716 5750 25774 6104
rect 25716 5458 25728 5750
rect 25762 5458 25774 5750
rect 25716 5104 25774 5458
rect 26774 5750 26832 6104
rect 26774 5458 26786 5750
rect 26820 5458 26832 5750
rect 26774 5104 26832 5458
rect 28006 6568 28018 6860
rect 28052 6568 28064 6860
rect 28006 6214 28064 6568
rect 29064 6860 29122 7214
rect 29064 6568 29076 6860
rect 29110 6568 29122 6860
rect 29064 6214 29122 6568
rect 30122 6860 30180 7214
rect 30122 6568 30134 6860
rect 30168 6568 30180 6860
rect 30122 6214 30180 6568
rect 31180 6860 31238 7214
rect 31180 6568 31192 6860
rect 31226 6568 31238 6860
rect 31180 6214 31238 6568
rect 32238 6860 32296 7214
rect 32238 6568 32250 6860
rect 32284 6568 32296 6860
rect 32238 6214 32296 6568
rect 33296 6860 33354 7214
rect 33296 6568 33308 6860
rect 33342 6568 33354 6860
rect 34516 6866 34574 7220
rect 33296 6214 33354 6568
rect 20284 4380 20296 4672
rect 20330 4380 20342 4672
rect 20284 4026 20342 4380
rect 21484 4656 21542 5010
rect 21484 4364 21496 4656
rect 21530 4364 21542 4656
rect 21484 4010 21542 4364
rect 22542 4656 22600 5010
rect 22542 4364 22554 4656
rect 22588 4364 22600 4656
rect 22542 4010 22600 4364
rect 23600 4656 23658 5010
rect 23600 4364 23612 4656
rect 23646 4364 23658 4656
rect 23600 4010 23658 4364
rect 24658 4656 24716 5010
rect 24658 4364 24670 4656
rect 24704 4364 24716 4656
rect 24658 4010 24716 4364
rect 25716 4656 25774 5010
rect 25716 4364 25728 4656
rect 25762 4364 25774 4656
rect 25716 4010 25774 4364
rect 26774 4656 26832 5010
rect 28006 5766 28064 6120
rect 28006 5474 28018 5766
rect 28052 5474 28064 5766
rect 28006 5120 28064 5474
rect 29064 5766 29122 6120
rect 29064 5474 29076 5766
rect 29110 5474 29122 5766
rect 29064 5120 29122 5474
rect 30122 5766 30180 6120
rect 30122 5474 30134 5766
rect 30168 5474 30180 5766
rect 30122 5120 30180 5474
rect 31180 5766 31238 6120
rect 31180 5474 31192 5766
rect 31226 5474 31238 5766
rect 31180 5120 31238 5474
rect 32238 5766 32296 6120
rect 32238 5474 32250 5766
rect 32284 5474 32296 5766
rect 32238 5120 32296 5474
rect 33296 5766 33354 6120
rect 33296 5474 33308 5766
rect 33342 5474 33354 5766
rect 33296 5120 33354 5474
rect 34516 6574 34528 6866
rect 34562 6574 34574 6866
rect 34516 6220 34574 6574
rect 35574 6866 35632 7220
rect 35574 6574 35586 6866
rect 35620 6574 35632 6866
rect 35574 6220 35632 6574
rect 36632 6866 36690 7220
rect 36632 6574 36644 6866
rect 36678 6574 36690 6866
rect 36632 6220 36690 6574
rect 37690 6866 37748 7220
rect 37690 6574 37702 6866
rect 37736 6574 37748 6866
rect 37690 6220 37748 6574
rect 38748 6866 38806 7220
rect 38748 6574 38760 6866
rect 38794 6574 38806 6866
rect 38748 6220 38806 6574
rect 39806 6866 39864 7220
rect 39806 6574 39818 6866
rect 39852 6574 39864 6866
rect 41006 6866 41064 7220
rect 39806 6220 39864 6574
rect 26774 4364 26786 4656
rect 26820 4364 26832 4656
rect 26774 4010 26832 4364
rect 28006 4672 28064 5026
rect 28006 4380 28018 4672
rect 28052 4380 28064 4672
rect 28006 4026 28064 4380
rect 29064 4672 29122 5026
rect 29064 4380 29076 4672
rect 29110 4380 29122 4672
rect 29064 4026 29122 4380
rect 30122 4672 30180 5026
rect 30122 4380 30134 4672
rect 30168 4380 30180 4672
rect 30122 4026 30180 4380
rect 31180 4672 31238 5026
rect 31180 4380 31192 4672
rect 31226 4380 31238 4672
rect 31180 4026 31238 4380
rect 32238 4672 32296 5026
rect 32238 4380 32250 4672
rect 32284 4380 32296 4672
rect 32238 4026 32296 4380
rect 33296 4672 33354 5026
rect 34516 5772 34574 6126
rect 34516 5480 34528 5772
rect 34562 5480 34574 5772
rect 34516 5126 34574 5480
rect 35574 5772 35632 6126
rect 35574 5480 35586 5772
rect 35620 5480 35632 5772
rect 35574 5126 35632 5480
rect 36632 5772 36690 6126
rect 36632 5480 36644 5772
rect 36678 5480 36690 5772
rect 36632 5126 36690 5480
rect 37690 5772 37748 6126
rect 37690 5480 37702 5772
rect 37736 5480 37748 5772
rect 37690 5126 37748 5480
rect 38748 5772 38806 6126
rect 38748 5480 38760 5772
rect 38794 5480 38806 5772
rect 38748 5126 38806 5480
rect 39806 5772 39864 6126
rect 39806 5480 39818 5772
rect 39852 5480 39864 5772
rect 39806 5126 39864 5480
rect 41006 6574 41018 6866
rect 41052 6574 41064 6866
rect 41006 6220 41064 6574
rect 42064 6866 42122 7220
rect 42064 6574 42076 6866
rect 42110 6574 42122 6866
rect 42064 6220 42122 6574
rect 43122 6866 43180 7220
rect 43122 6574 43134 6866
rect 43168 6574 43180 6866
rect 43122 6220 43180 6574
rect 44180 6866 44238 7220
rect 44180 6574 44192 6866
rect 44226 6574 44238 6866
rect 44180 6220 44238 6574
rect 45238 6866 45296 7220
rect 45238 6574 45250 6866
rect 45284 6574 45296 6866
rect 45238 6220 45296 6574
rect 46296 6866 46354 7220
rect 46296 6574 46308 6866
rect 46342 6574 46354 6866
rect 47594 6888 47652 7242
rect 46296 6220 46354 6574
rect 33296 4380 33308 4672
rect 33342 4380 33354 4672
rect 33296 4026 33354 4380
rect 34516 4678 34574 5032
rect 34516 4386 34528 4678
rect 34562 4386 34574 4678
rect 34516 4032 34574 4386
rect 35574 4678 35632 5032
rect 35574 4386 35586 4678
rect 35620 4386 35632 4678
rect 35574 4032 35632 4386
rect 36632 4678 36690 5032
rect 36632 4386 36644 4678
rect 36678 4386 36690 4678
rect 36632 4032 36690 4386
rect 37690 4678 37748 5032
rect 37690 4386 37702 4678
rect 37736 4386 37748 4678
rect 37690 4032 37748 4386
rect 38748 4678 38806 5032
rect 38748 4386 38760 4678
rect 38794 4386 38806 4678
rect 38748 4032 38806 4386
rect 39806 4678 39864 5032
rect 41006 5772 41064 6126
rect 41006 5480 41018 5772
rect 41052 5480 41064 5772
rect 41006 5126 41064 5480
rect 42064 5772 42122 6126
rect 42064 5480 42076 5772
rect 42110 5480 42122 5772
rect 42064 5126 42122 5480
rect 43122 5772 43180 6126
rect 43122 5480 43134 5772
rect 43168 5480 43180 5772
rect 43122 5126 43180 5480
rect 44180 5772 44238 6126
rect 44180 5480 44192 5772
rect 44226 5480 44238 5772
rect 44180 5126 44238 5480
rect 45238 5772 45296 6126
rect 45238 5480 45250 5772
rect 45284 5480 45296 5772
rect 45238 5126 45296 5480
rect 46296 5772 46354 6126
rect 46296 5480 46308 5772
rect 46342 5480 46354 5772
rect 46296 5126 46354 5480
rect 47594 6596 47606 6888
rect 47640 6596 47652 6888
rect 47594 6242 47652 6596
rect 48652 6888 48710 7242
rect 48652 6596 48664 6888
rect 48698 6596 48710 6888
rect 48652 6242 48710 6596
rect 49710 6888 49768 7242
rect 49710 6596 49722 6888
rect 49756 6596 49768 6888
rect 49710 6242 49768 6596
rect 50768 6888 50826 7242
rect 50768 6596 50780 6888
rect 50814 6596 50826 6888
rect 50768 6242 50826 6596
rect 51826 6888 51884 7242
rect 51826 6596 51838 6888
rect 51872 6596 51884 6888
rect 51826 6242 51884 6596
rect 52884 6888 52942 7242
rect 52884 6596 52896 6888
rect 52930 6596 52942 6888
rect 54108 6902 54166 7256
rect 52884 6242 52942 6596
rect 39806 4386 39818 4678
rect 39852 4386 39864 4678
rect 39806 4032 39864 4386
rect 41006 4678 41064 5032
rect 41006 4386 41018 4678
rect 41052 4386 41064 4678
rect 41006 4032 41064 4386
rect 42064 4678 42122 5032
rect 42064 4386 42076 4678
rect 42110 4386 42122 4678
rect 42064 4032 42122 4386
rect 43122 4678 43180 5032
rect 43122 4386 43134 4678
rect 43168 4386 43180 4678
rect 43122 4032 43180 4386
rect 44180 4678 44238 5032
rect 44180 4386 44192 4678
rect 44226 4386 44238 4678
rect 44180 4032 44238 4386
rect 45238 4678 45296 5032
rect 45238 4386 45250 4678
rect 45284 4386 45296 4678
rect 45238 4032 45296 4386
rect 46296 4678 46354 5032
rect 47594 5794 47652 6148
rect 47594 5502 47606 5794
rect 47640 5502 47652 5794
rect 47594 5148 47652 5502
rect 48652 5794 48710 6148
rect 48652 5502 48664 5794
rect 48698 5502 48710 5794
rect 48652 5148 48710 5502
rect 49710 5794 49768 6148
rect 49710 5502 49722 5794
rect 49756 5502 49768 5794
rect 49710 5148 49768 5502
rect 50768 5794 50826 6148
rect 50768 5502 50780 5794
rect 50814 5502 50826 5794
rect 50768 5148 50826 5502
rect 51826 5794 51884 6148
rect 51826 5502 51838 5794
rect 51872 5502 51884 5794
rect 51826 5148 51884 5502
rect 52884 5794 52942 6148
rect 52884 5502 52896 5794
rect 52930 5502 52942 5794
rect 52884 5148 52942 5502
rect 54108 6610 54120 6902
rect 54154 6610 54166 6902
rect 54108 6256 54166 6610
rect 55166 6902 55224 7256
rect 55166 6610 55178 6902
rect 55212 6610 55224 6902
rect 55166 6256 55224 6610
rect 56224 6902 56282 7256
rect 56224 6610 56236 6902
rect 56270 6610 56282 6902
rect 56224 6256 56282 6610
rect 57282 6902 57340 7256
rect 57282 6610 57294 6902
rect 57328 6610 57340 6902
rect 57282 6256 57340 6610
rect 58340 6902 58398 7256
rect 58340 6610 58352 6902
rect 58386 6610 58398 6902
rect 58340 6256 58398 6610
rect 59398 6902 59456 7256
rect 59398 6610 59410 6902
rect 59444 6610 59456 6902
rect 59398 6256 59456 6610
rect 46296 4386 46308 4678
rect 46342 4386 46354 4678
rect 46296 4032 46354 4386
rect 47594 4700 47652 5054
rect 47594 4408 47606 4700
rect 47640 4408 47652 4700
rect 47594 4054 47652 4408
rect 48652 4700 48710 5054
rect 48652 4408 48664 4700
rect 48698 4408 48710 4700
rect 48652 4054 48710 4408
rect 49710 4700 49768 5054
rect 49710 4408 49722 4700
rect 49756 4408 49768 4700
rect 49710 4054 49768 4408
rect 50768 4700 50826 5054
rect 50768 4408 50780 4700
rect 50814 4408 50826 4700
rect 50768 4054 50826 4408
rect 51826 4700 51884 5054
rect 51826 4408 51838 4700
rect 51872 4408 51884 4700
rect 51826 4054 51884 4408
rect 52884 4700 52942 5054
rect 54108 5808 54166 6162
rect 54108 5516 54120 5808
rect 54154 5516 54166 5808
rect 54108 5162 54166 5516
rect 55166 5808 55224 6162
rect 55166 5516 55178 5808
rect 55212 5516 55224 5808
rect 55166 5162 55224 5516
rect 56224 5808 56282 6162
rect 56224 5516 56236 5808
rect 56270 5516 56282 5808
rect 56224 5162 56282 5516
rect 57282 5808 57340 6162
rect 57282 5516 57294 5808
rect 57328 5516 57340 5808
rect 57282 5162 57340 5516
rect 58340 5808 58398 6162
rect 58340 5516 58352 5808
rect 58386 5516 58398 5808
rect 58340 5162 58398 5516
rect 59398 5808 59456 6162
rect 59398 5516 59410 5808
rect 59444 5516 59456 5808
rect 59398 5162 59456 5516
rect 52884 4408 52896 4700
rect 52930 4408 52942 4700
rect 52884 4054 52942 4408
rect 54108 4714 54166 5068
rect 54108 4422 54120 4714
rect 54154 4422 54166 4714
rect 54108 4068 54166 4422
rect 55166 4714 55224 5068
rect 55166 4422 55178 4714
rect 55212 4422 55224 4714
rect 55166 4068 55224 4422
rect 56224 4714 56282 5068
rect 56224 4422 56236 4714
rect 56270 4422 56282 4714
rect 56224 4068 56282 4422
rect 57282 4714 57340 5068
rect 57282 4422 57294 4714
rect 57328 4422 57340 4714
rect 57282 4068 57340 4422
rect 58340 4714 58398 5068
rect 58340 4422 58352 4714
rect 58386 4422 58398 4714
rect 58340 4068 58398 4422
rect 59398 4714 59456 5068
rect 59398 4422 59410 4714
rect 59444 4422 59456 4714
rect 59398 4068 59456 4422
rect 1974 3562 2032 3916
rect 1974 3270 1986 3562
rect 2020 3270 2032 3562
rect 1974 2916 2032 3270
rect 3032 3562 3090 3916
rect 3032 3270 3044 3562
rect 3078 3270 3090 3562
rect 3032 2916 3090 3270
rect 4090 3562 4148 3916
rect 4090 3270 4102 3562
rect 4136 3270 4148 3562
rect 4090 2916 4148 3270
rect 5148 3562 5206 3916
rect 5148 3270 5160 3562
rect 5194 3270 5206 3562
rect 5148 2916 5206 3270
rect 6206 3562 6264 3916
rect 6206 3270 6218 3562
rect 6252 3270 6264 3562
rect 6206 2916 6264 3270
rect 7264 3562 7322 3916
rect 7264 3270 7276 3562
rect 7310 3270 7322 3562
rect 7264 2916 7322 3270
rect 8488 3570 8546 3924
rect 8488 3278 8500 3570
rect 8534 3278 8546 3570
rect 8488 2924 8546 3278
rect 9546 3570 9604 3924
rect 9546 3278 9558 3570
rect 9592 3278 9604 3570
rect 9546 2924 9604 3278
rect 10604 3570 10662 3924
rect 10604 3278 10616 3570
rect 10650 3278 10662 3570
rect 10604 2924 10662 3278
rect 11662 3570 11720 3924
rect 11662 3278 11674 3570
rect 11708 3278 11720 3570
rect 11662 2924 11720 3278
rect 12720 3570 12778 3924
rect 12720 3278 12732 3570
rect 12766 3278 12778 3570
rect 12720 2924 12778 3278
rect 13778 3570 13836 3924
rect 13778 3278 13790 3570
rect 13824 3278 13836 3570
rect 13778 2924 13836 3278
rect 14994 3578 15052 3932
rect 14994 3286 15006 3578
rect 15040 3286 15052 3578
rect 14994 2932 15052 3286
rect 16052 3578 16110 3932
rect 16052 3286 16064 3578
rect 16098 3286 16110 3578
rect 16052 2932 16110 3286
rect 17110 3578 17168 3932
rect 17110 3286 17122 3578
rect 17156 3286 17168 3578
rect 17110 2932 17168 3286
rect 18168 3578 18226 3932
rect 18168 3286 18180 3578
rect 18214 3286 18226 3578
rect 18168 2932 18226 3286
rect 19226 3578 19284 3932
rect 19226 3286 19238 3578
rect 19272 3286 19284 3578
rect 19226 2932 19284 3286
rect 20284 3578 20342 3932
rect 20284 3286 20296 3578
rect 20330 3286 20342 3578
rect 20284 2932 20342 3286
rect 21484 3562 21542 3916
rect 21484 3270 21496 3562
rect 21530 3270 21542 3562
rect 21484 2916 21542 3270
rect 22542 3562 22600 3916
rect 22542 3270 22554 3562
rect 22588 3270 22600 3562
rect 22542 2916 22600 3270
rect 23600 3562 23658 3916
rect 23600 3270 23612 3562
rect 23646 3270 23658 3562
rect 23600 2916 23658 3270
rect 24658 3562 24716 3916
rect 24658 3270 24670 3562
rect 24704 3270 24716 3562
rect 24658 2916 24716 3270
rect 25716 3562 25774 3916
rect 25716 3270 25728 3562
rect 25762 3270 25774 3562
rect 25716 2916 25774 3270
rect 26774 3562 26832 3916
rect 26774 3270 26786 3562
rect 26820 3270 26832 3562
rect 26774 2916 26832 3270
rect 28006 3578 28064 3932
rect 28006 3286 28018 3578
rect 28052 3286 28064 3578
rect 28006 2932 28064 3286
rect 29064 3578 29122 3932
rect 29064 3286 29076 3578
rect 29110 3286 29122 3578
rect 29064 2932 29122 3286
rect 30122 3578 30180 3932
rect 30122 3286 30134 3578
rect 30168 3286 30180 3578
rect 30122 2932 30180 3286
rect 31180 3578 31238 3932
rect 31180 3286 31192 3578
rect 31226 3286 31238 3578
rect 31180 2932 31238 3286
rect 32238 3578 32296 3932
rect 32238 3286 32250 3578
rect 32284 3286 32296 3578
rect 32238 2932 32296 3286
rect 33296 3578 33354 3932
rect 33296 3286 33308 3578
rect 33342 3286 33354 3578
rect 33296 2932 33354 3286
rect 34516 3584 34574 3938
rect 34516 3292 34528 3584
rect 34562 3292 34574 3584
rect 34516 2938 34574 3292
rect 35574 3584 35632 3938
rect 35574 3292 35586 3584
rect 35620 3292 35632 3584
rect 35574 2938 35632 3292
rect 36632 3584 36690 3938
rect 36632 3292 36644 3584
rect 36678 3292 36690 3584
rect 36632 2938 36690 3292
rect 37690 3584 37748 3938
rect 37690 3292 37702 3584
rect 37736 3292 37748 3584
rect 37690 2938 37748 3292
rect 38748 3584 38806 3938
rect 38748 3292 38760 3584
rect 38794 3292 38806 3584
rect 38748 2938 38806 3292
rect 39806 3584 39864 3938
rect 39806 3292 39818 3584
rect 39852 3292 39864 3584
rect 39806 2938 39864 3292
rect 41006 3584 41064 3938
rect 41006 3292 41018 3584
rect 41052 3292 41064 3584
rect 41006 2938 41064 3292
rect 42064 3584 42122 3938
rect 42064 3292 42076 3584
rect 42110 3292 42122 3584
rect 42064 2938 42122 3292
rect 43122 3584 43180 3938
rect 43122 3292 43134 3584
rect 43168 3292 43180 3584
rect 43122 2938 43180 3292
rect 44180 3584 44238 3938
rect 44180 3292 44192 3584
rect 44226 3292 44238 3584
rect 44180 2938 44238 3292
rect 45238 3584 45296 3938
rect 45238 3292 45250 3584
rect 45284 3292 45296 3584
rect 45238 2938 45296 3292
rect 46296 3584 46354 3938
rect 46296 3292 46308 3584
rect 46342 3292 46354 3584
rect 46296 2938 46354 3292
rect 47594 3606 47652 3960
rect 47594 3314 47606 3606
rect 47640 3314 47652 3606
rect 47594 2960 47652 3314
rect 48652 3606 48710 3960
rect 48652 3314 48664 3606
rect 48698 3314 48710 3606
rect 48652 2960 48710 3314
rect 49710 3606 49768 3960
rect 49710 3314 49722 3606
rect 49756 3314 49768 3606
rect 49710 2960 49768 3314
rect 50768 3606 50826 3960
rect 50768 3314 50780 3606
rect 50814 3314 50826 3606
rect 50768 2960 50826 3314
rect 51826 3606 51884 3960
rect 51826 3314 51838 3606
rect 51872 3314 51884 3606
rect 51826 2960 51884 3314
rect 52884 3606 52942 3960
rect 52884 3314 52896 3606
rect 52930 3314 52942 3606
rect 52884 2960 52942 3314
rect 54108 3620 54166 3974
rect 54108 3328 54120 3620
rect 54154 3328 54166 3620
rect 54108 2974 54166 3328
rect 55166 3620 55224 3974
rect 55166 3328 55178 3620
rect 55212 3328 55224 3620
rect 55166 2974 55224 3328
rect 56224 3620 56282 3974
rect 56224 3328 56236 3620
rect 56270 3328 56282 3620
rect 56224 2974 56282 3328
rect 57282 3620 57340 3974
rect 57282 3328 57294 3620
rect 57328 3328 57340 3620
rect 57282 2974 57340 3328
rect 58340 3620 58398 3974
rect 58340 3328 58352 3620
rect 58386 3328 58398 3620
rect 58340 2974 58398 3328
rect 59398 3620 59456 3974
rect 59398 3328 59410 3620
rect 59444 3328 59456 3620
rect 59398 2974 59456 3328
rect 62100 25568 62158 25922
rect 62100 25276 62112 25568
rect 62146 25276 62158 25568
rect 62100 24922 62158 25276
rect 63158 25568 63216 25922
rect 63158 25276 63170 25568
rect 63204 25276 63216 25568
rect 63158 24922 63216 25276
rect 64216 25568 64274 25922
rect 64216 25276 64228 25568
rect 64262 25276 64274 25568
rect 64216 24922 64274 25276
rect 65274 25568 65332 25922
rect 65274 25276 65286 25568
rect 65320 25276 65332 25568
rect 65274 24922 65332 25276
rect 66332 25568 66390 25922
rect 66332 25276 66344 25568
rect 66378 25276 66390 25568
rect 66332 24922 66390 25276
rect 67390 25568 67448 25922
rect 67390 25276 67402 25568
rect 67436 25276 67448 25568
rect 67390 24922 67448 25276
rect 68562 25566 68620 25920
rect 68562 25274 68574 25566
rect 68608 25274 68620 25566
rect 68562 24920 68620 25274
rect 69620 25566 69678 25920
rect 69620 25274 69632 25566
rect 69666 25274 69678 25566
rect 69620 24920 69678 25274
rect 70678 25566 70736 25920
rect 70678 25274 70690 25566
rect 70724 25274 70736 25566
rect 70678 24920 70736 25274
rect 71736 25566 71794 25920
rect 71736 25274 71748 25566
rect 71782 25274 71794 25566
rect 71736 24920 71794 25274
rect 72794 25566 72852 25920
rect 72794 25274 72806 25566
rect 72840 25274 72852 25566
rect 72794 24920 72852 25274
rect 73852 25566 73910 25920
rect 73852 25274 73864 25566
rect 73898 25274 73910 25566
rect 73852 24920 73910 25274
rect 75256 25540 75314 25894
rect 75256 25248 75268 25540
rect 75302 25248 75314 25540
rect 75256 24894 75314 25248
rect 76314 25540 76372 25894
rect 76314 25248 76326 25540
rect 76360 25248 76372 25540
rect 76314 24894 76372 25248
rect 77372 25540 77430 25894
rect 77372 25248 77384 25540
rect 77418 25248 77430 25540
rect 77372 24894 77430 25248
rect 78430 25540 78488 25894
rect 78430 25248 78442 25540
rect 78476 25248 78488 25540
rect 78430 24894 78488 25248
rect 79488 25540 79546 25894
rect 79488 25248 79500 25540
rect 79534 25248 79546 25540
rect 79488 24894 79546 25248
rect 80546 25540 80604 25894
rect 80546 25248 80558 25540
rect 80592 25248 80604 25540
rect 80546 24894 80604 25248
rect 81718 25538 81776 25892
rect 81718 25246 81730 25538
rect 81764 25246 81776 25538
rect 81718 24892 81776 25246
rect 82776 25538 82834 25892
rect 82776 25246 82788 25538
rect 82822 25246 82834 25538
rect 82776 24892 82834 25246
rect 83834 25538 83892 25892
rect 83834 25246 83846 25538
rect 83880 25246 83892 25538
rect 83834 24892 83892 25246
rect 84892 25538 84950 25892
rect 84892 25246 84904 25538
rect 84938 25246 84950 25538
rect 84892 24892 84950 25246
rect 85950 25538 86008 25892
rect 85950 25246 85962 25538
rect 85996 25246 86008 25538
rect 85950 24892 86008 25246
rect 87008 25538 87066 25892
rect 87008 25246 87020 25538
rect 87054 25246 87066 25538
rect 87008 24892 87066 25246
rect 88490 25532 88548 25886
rect 88490 25240 88502 25532
rect 88536 25240 88548 25532
rect 62100 24474 62158 24828
rect 62100 24182 62112 24474
rect 62146 24182 62158 24474
rect 62100 23828 62158 24182
rect 63158 24474 63216 24828
rect 63158 24182 63170 24474
rect 63204 24182 63216 24474
rect 63158 23828 63216 24182
rect 64216 24474 64274 24828
rect 64216 24182 64228 24474
rect 64262 24182 64274 24474
rect 64216 23828 64274 24182
rect 65274 24474 65332 24828
rect 65274 24182 65286 24474
rect 65320 24182 65332 24474
rect 65274 23828 65332 24182
rect 66332 24474 66390 24828
rect 66332 24182 66344 24474
rect 66378 24182 66390 24474
rect 66332 23828 66390 24182
rect 67390 24474 67448 24828
rect 88490 24886 88548 25240
rect 89548 25532 89606 25886
rect 89548 25240 89560 25532
rect 89594 25240 89606 25532
rect 89548 24886 89606 25240
rect 90606 25532 90664 25886
rect 90606 25240 90618 25532
rect 90652 25240 90664 25532
rect 90606 24886 90664 25240
rect 91664 25532 91722 25886
rect 91664 25240 91676 25532
rect 91710 25240 91722 25532
rect 91664 24886 91722 25240
rect 92722 25532 92780 25886
rect 92722 25240 92734 25532
rect 92768 25240 92780 25532
rect 92722 24886 92780 25240
rect 93780 25532 93838 25886
rect 93780 25240 93792 25532
rect 93826 25240 93838 25532
rect 93780 24886 93838 25240
rect 94952 25530 95010 25884
rect 94952 25238 94964 25530
rect 94998 25238 95010 25530
rect 67390 24182 67402 24474
rect 67436 24182 67448 24474
rect 68562 24472 68620 24826
rect 67390 23828 67448 24182
rect 62100 23380 62158 23734
rect 62100 23088 62112 23380
rect 62146 23088 62158 23380
rect 62100 22734 62158 23088
rect 63158 23380 63216 23734
rect 63158 23088 63170 23380
rect 63204 23088 63216 23380
rect 63158 22734 63216 23088
rect 64216 23380 64274 23734
rect 64216 23088 64228 23380
rect 64262 23088 64274 23380
rect 64216 22734 64274 23088
rect 65274 23380 65332 23734
rect 65274 23088 65286 23380
rect 65320 23088 65332 23380
rect 65274 22734 65332 23088
rect 66332 23380 66390 23734
rect 66332 23088 66344 23380
rect 66378 23088 66390 23380
rect 66332 22734 66390 23088
rect 67390 23380 67448 23734
rect 67390 23088 67402 23380
rect 67436 23088 67448 23380
rect 67390 22734 67448 23088
rect 68562 24180 68574 24472
rect 68608 24180 68620 24472
rect 68562 23826 68620 24180
rect 69620 24472 69678 24826
rect 69620 24180 69632 24472
rect 69666 24180 69678 24472
rect 69620 23826 69678 24180
rect 70678 24472 70736 24826
rect 70678 24180 70690 24472
rect 70724 24180 70736 24472
rect 70678 23826 70736 24180
rect 71736 24472 71794 24826
rect 71736 24180 71748 24472
rect 71782 24180 71794 24472
rect 71736 23826 71794 24180
rect 72794 24472 72852 24826
rect 72794 24180 72806 24472
rect 72840 24180 72852 24472
rect 72794 23826 72852 24180
rect 73852 24472 73910 24826
rect 94952 24884 95010 25238
rect 96010 25530 96068 25884
rect 96010 25238 96022 25530
rect 96056 25238 96068 25530
rect 96010 24884 96068 25238
rect 97068 25530 97126 25884
rect 97068 25238 97080 25530
rect 97114 25238 97126 25530
rect 97068 24884 97126 25238
rect 98126 25530 98184 25884
rect 98126 25238 98138 25530
rect 98172 25238 98184 25530
rect 98126 24884 98184 25238
rect 99184 25530 99242 25884
rect 99184 25238 99196 25530
rect 99230 25238 99242 25530
rect 99184 24884 99242 25238
rect 100242 25530 100300 25884
rect 100242 25238 100254 25530
rect 100288 25238 100300 25530
rect 100242 24884 100300 25238
rect 73852 24180 73864 24472
rect 73898 24180 73910 24472
rect 73852 23826 73910 24180
rect 75256 24446 75314 24800
rect 62100 22286 62158 22640
rect 62100 21994 62112 22286
rect 62146 21994 62158 22286
rect 62100 21640 62158 21994
rect 63158 22286 63216 22640
rect 63158 21994 63170 22286
rect 63204 21994 63216 22286
rect 63158 21640 63216 21994
rect 64216 22286 64274 22640
rect 64216 21994 64228 22286
rect 64262 21994 64274 22286
rect 64216 21640 64274 21994
rect 65274 22286 65332 22640
rect 65274 21994 65286 22286
rect 65320 21994 65332 22286
rect 65274 21640 65332 21994
rect 66332 22286 66390 22640
rect 66332 21994 66344 22286
rect 66378 21994 66390 22286
rect 66332 21640 66390 21994
rect 67390 22286 67448 22640
rect 68562 23378 68620 23732
rect 68562 23086 68574 23378
rect 68608 23086 68620 23378
rect 68562 22732 68620 23086
rect 69620 23378 69678 23732
rect 69620 23086 69632 23378
rect 69666 23086 69678 23378
rect 69620 22732 69678 23086
rect 70678 23378 70736 23732
rect 70678 23086 70690 23378
rect 70724 23086 70736 23378
rect 70678 22732 70736 23086
rect 71736 23378 71794 23732
rect 71736 23086 71748 23378
rect 71782 23086 71794 23378
rect 71736 22732 71794 23086
rect 72794 23378 72852 23732
rect 72794 23086 72806 23378
rect 72840 23086 72852 23378
rect 72794 22732 72852 23086
rect 73852 23378 73910 23732
rect 73852 23086 73864 23378
rect 73898 23086 73910 23378
rect 73852 22732 73910 23086
rect 75256 24154 75268 24446
rect 75302 24154 75314 24446
rect 75256 23800 75314 24154
rect 76314 24446 76372 24800
rect 76314 24154 76326 24446
rect 76360 24154 76372 24446
rect 76314 23800 76372 24154
rect 77372 24446 77430 24800
rect 77372 24154 77384 24446
rect 77418 24154 77430 24446
rect 77372 23800 77430 24154
rect 78430 24446 78488 24800
rect 78430 24154 78442 24446
rect 78476 24154 78488 24446
rect 78430 23800 78488 24154
rect 79488 24446 79546 24800
rect 79488 24154 79500 24446
rect 79534 24154 79546 24446
rect 79488 23800 79546 24154
rect 80546 24446 80604 24800
rect 80546 24154 80558 24446
rect 80592 24154 80604 24446
rect 81718 24444 81776 24798
rect 80546 23800 80604 24154
rect 67390 21994 67402 22286
rect 67436 21994 67448 22286
rect 67390 21640 67448 21994
rect 68562 22284 68620 22638
rect 68562 21992 68574 22284
rect 68608 21992 68620 22284
rect 68562 21638 68620 21992
rect 69620 22284 69678 22638
rect 69620 21992 69632 22284
rect 69666 21992 69678 22284
rect 69620 21638 69678 21992
rect 70678 22284 70736 22638
rect 70678 21992 70690 22284
rect 70724 21992 70736 22284
rect 70678 21638 70736 21992
rect 71736 22284 71794 22638
rect 71736 21992 71748 22284
rect 71782 21992 71794 22284
rect 71736 21638 71794 21992
rect 72794 22284 72852 22638
rect 72794 21992 72806 22284
rect 72840 21992 72852 22284
rect 72794 21638 72852 21992
rect 73852 22284 73910 22638
rect 75256 23352 75314 23706
rect 75256 23060 75268 23352
rect 75302 23060 75314 23352
rect 75256 22706 75314 23060
rect 76314 23352 76372 23706
rect 76314 23060 76326 23352
rect 76360 23060 76372 23352
rect 76314 22706 76372 23060
rect 77372 23352 77430 23706
rect 77372 23060 77384 23352
rect 77418 23060 77430 23352
rect 77372 22706 77430 23060
rect 78430 23352 78488 23706
rect 78430 23060 78442 23352
rect 78476 23060 78488 23352
rect 78430 22706 78488 23060
rect 79488 23352 79546 23706
rect 79488 23060 79500 23352
rect 79534 23060 79546 23352
rect 79488 22706 79546 23060
rect 80546 23352 80604 23706
rect 80546 23060 80558 23352
rect 80592 23060 80604 23352
rect 80546 22706 80604 23060
rect 81718 24152 81730 24444
rect 81764 24152 81776 24444
rect 81718 23798 81776 24152
rect 82776 24444 82834 24798
rect 82776 24152 82788 24444
rect 82822 24152 82834 24444
rect 82776 23798 82834 24152
rect 83834 24444 83892 24798
rect 83834 24152 83846 24444
rect 83880 24152 83892 24444
rect 83834 23798 83892 24152
rect 84892 24444 84950 24798
rect 84892 24152 84904 24444
rect 84938 24152 84950 24444
rect 84892 23798 84950 24152
rect 85950 24444 86008 24798
rect 85950 24152 85962 24444
rect 85996 24152 86008 24444
rect 85950 23798 86008 24152
rect 87008 24444 87066 24798
rect 87008 24152 87020 24444
rect 87054 24152 87066 24444
rect 88490 24438 88548 24792
rect 87008 23798 87066 24152
rect 73852 21992 73864 22284
rect 73898 21992 73910 22284
rect 73852 21638 73910 21992
rect 75256 22258 75314 22612
rect 75256 21966 75268 22258
rect 75302 21966 75314 22258
rect 75256 21612 75314 21966
rect 76314 22258 76372 22612
rect 76314 21966 76326 22258
rect 76360 21966 76372 22258
rect 76314 21612 76372 21966
rect 77372 22258 77430 22612
rect 77372 21966 77384 22258
rect 77418 21966 77430 22258
rect 77372 21612 77430 21966
rect 78430 22258 78488 22612
rect 78430 21966 78442 22258
rect 78476 21966 78488 22258
rect 78430 21612 78488 21966
rect 79488 22258 79546 22612
rect 79488 21966 79500 22258
rect 79534 21966 79546 22258
rect 79488 21612 79546 21966
rect 80546 22258 80604 22612
rect 81718 23350 81776 23704
rect 81718 23058 81730 23350
rect 81764 23058 81776 23350
rect 81718 22704 81776 23058
rect 82776 23350 82834 23704
rect 82776 23058 82788 23350
rect 82822 23058 82834 23350
rect 82776 22704 82834 23058
rect 83834 23350 83892 23704
rect 83834 23058 83846 23350
rect 83880 23058 83892 23350
rect 83834 22704 83892 23058
rect 84892 23350 84950 23704
rect 84892 23058 84904 23350
rect 84938 23058 84950 23350
rect 84892 22704 84950 23058
rect 85950 23350 86008 23704
rect 85950 23058 85962 23350
rect 85996 23058 86008 23350
rect 85950 22704 86008 23058
rect 87008 23350 87066 23704
rect 87008 23058 87020 23350
rect 87054 23058 87066 23350
rect 87008 22704 87066 23058
rect 88490 24146 88502 24438
rect 88536 24146 88548 24438
rect 88490 23792 88548 24146
rect 89548 24438 89606 24792
rect 89548 24146 89560 24438
rect 89594 24146 89606 24438
rect 89548 23792 89606 24146
rect 90606 24438 90664 24792
rect 90606 24146 90618 24438
rect 90652 24146 90664 24438
rect 90606 23792 90664 24146
rect 91664 24438 91722 24792
rect 91664 24146 91676 24438
rect 91710 24146 91722 24438
rect 91664 23792 91722 24146
rect 92722 24438 92780 24792
rect 92722 24146 92734 24438
rect 92768 24146 92780 24438
rect 92722 23792 92780 24146
rect 93780 24438 93838 24792
rect 93780 24146 93792 24438
rect 93826 24146 93838 24438
rect 94952 24436 95010 24790
rect 93780 23792 93838 24146
rect 80546 21966 80558 22258
rect 80592 21966 80604 22258
rect 80546 21612 80604 21966
rect 81718 22256 81776 22610
rect 81718 21964 81730 22256
rect 81764 21964 81776 22256
rect 81718 21610 81776 21964
rect 82776 22256 82834 22610
rect 82776 21964 82788 22256
rect 82822 21964 82834 22256
rect 82776 21610 82834 21964
rect 83834 22256 83892 22610
rect 83834 21964 83846 22256
rect 83880 21964 83892 22256
rect 83834 21610 83892 21964
rect 84892 22256 84950 22610
rect 84892 21964 84904 22256
rect 84938 21964 84950 22256
rect 84892 21610 84950 21964
rect 85950 22256 86008 22610
rect 85950 21964 85962 22256
rect 85996 21964 86008 22256
rect 85950 21610 86008 21964
rect 87008 22256 87066 22610
rect 88490 23344 88548 23698
rect 88490 23052 88502 23344
rect 88536 23052 88548 23344
rect 88490 22698 88548 23052
rect 89548 23344 89606 23698
rect 89548 23052 89560 23344
rect 89594 23052 89606 23344
rect 89548 22698 89606 23052
rect 90606 23344 90664 23698
rect 90606 23052 90618 23344
rect 90652 23052 90664 23344
rect 90606 22698 90664 23052
rect 91664 23344 91722 23698
rect 91664 23052 91676 23344
rect 91710 23052 91722 23344
rect 91664 22698 91722 23052
rect 92722 23344 92780 23698
rect 92722 23052 92734 23344
rect 92768 23052 92780 23344
rect 92722 22698 92780 23052
rect 93780 23344 93838 23698
rect 93780 23052 93792 23344
rect 93826 23052 93838 23344
rect 93780 22698 93838 23052
rect 94952 24144 94964 24436
rect 94998 24144 95010 24436
rect 94952 23790 95010 24144
rect 96010 24436 96068 24790
rect 96010 24144 96022 24436
rect 96056 24144 96068 24436
rect 96010 23790 96068 24144
rect 97068 24436 97126 24790
rect 97068 24144 97080 24436
rect 97114 24144 97126 24436
rect 97068 23790 97126 24144
rect 98126 24436 98184 24790
rect 98126 24144 98138 24436
rect 98172 24144 98184 24436
rect 98126 23790 98184 24144
rect 99184 24436 99242 24790
rect 99184 24144 99196 24436
rect 99230 24144 99242 24436
rect 99184 23790 99242 24144
rect 100242 24436 100300 24790
rect 100242 24144 100254 24436
rect 100288 24144 100300 24436
rect 100242 23790 100300 24144
rect 87008 21964 87020 22256
rect 87054 21964 87066 22256
rect 87008 21610 87066 21964
rect 88490 22250 88548 22604
rect 88490 21958 88502 22250
rect 88536 21958 88548 22250
rect 62100 21192 62158 21546
rect 62100 20900 62112 21192
rect 62146 20900 62158 21192
rect 62100 20546 62158 20900
rect 63158 21192 63216 21546
rect 63158 20900 63170 21192
rect 63204 20900 63216 21192
rect 63158 20546 63216 20900
rect 64216 21192 64274 21546
rect 64216 20900 64228 21192
rect 64262 20900 64274 21192
rect 64216 20546 64274 20900
rect 65274 21192 65332 21546
rect 65274 20900 65286 21192
rect 65320 20900 65332 21192
rect 65274 20546 65332 20900
rect 66332 21192 66390 21546
rect 66332 20900 66344 21192
rect 66378 20900 66390 21192
rect 66332 20546 66390 20900
rect 67390 21192 67448 21546
rect 88490 21604 88548 21958
rect 89548 22250 89606 22604
rect 89548 21958 89560 22250
rect 89594 21958 89606 22250
rect 89548 21604 89606 21958
rect 90606 22250 90664 22604
rect 90606 21958 90618 22250
rect 90652 21958 90664 22250
rect 90606 21604 90664 21958
rect 91664 22250 91722 22604
rect 91664 21958 91676 22250
rect 91710 21958 91722 22250
rect 91664 21604 91722 21958
rect 92722 22250 92780 22604
rect 92722 21958 92734 22250
rect 92768 21958 92780 22250
rect 92722 21604 92780 21958
rect 93780 22250 93838 22604
rect 94952 23342 95010 23696
rect 94952 23050 94964 23342
rect 94998 23050 95010 23342
rect 94952 22696 95010 23050
rect 96010 23342 96068 23696
rect 96010 23050 96022 23342
rect 96056 23050 96068 23342
rect 96010 22696 96068 23050
rect 97068 23342 97126 23696
rect 97068 23050 97080 23342
rect 97114 23050 97126 23342
rect 97068 22696 97126 23050
rect 98126 23342 98184 23696
rect 98126 23050 98138 23342
rect 98172 23050 98184 23342
rect 98126 22696 98184 23050
rect 99184 23342 99242 23696
rect 99184 23050 99196 23342
rect 99230 23050 99242 23342
rect 99184 22696 99242 23050
rect 100242 23342 100300 23696
rect 100242 23050 100254 23342
rect 100288 23050 100300 23342
rect 100242 22696 100300 23050
rect 93780 21958 93792 22250
rect 93826 21958 93838 22250
rect 93780 21604 93838 21958
rect 94952 22248 95010 22602
rect 94952 21956 94964 22248
rect 94998 21956 95010 22248
rect 67390 20900 67402 21192
rect 67436 20900 67448 21192
rect 67390 20546 67448 20900
rect 68562 21190 68620 21544
rect 68562 20898 68574 21190
rect 68608 20898 68620 21190
rect 68562 20544 68620 20898
rect 69620 21190 69678 21544
rect 69620 20898 69632 21190
rect 69666 20898 69678 21190
rect 69620 20544 69678 20898
rect 70678 21190 70736 21544
rect 70678 20898 70690 21190
rect 70724 20898 70736 21190
rect 70678 20544 70736 20898
rect 71736 21190 71794 21544
rect 71736 20898 71748 21190
rect 71782 20898 71794 21190
rect 71736 20544 71794 20898
rect 72794 21190 72852 21544
rect 72794 20898 72806 21190
rect 72840 20898 72852 21190
rect 72794 20544 72852 20898
rect 73852 21190 73910 21544
rect 94952 21602 95010 21956
rect 96010 22248 96068 22602
rect 96010 21956 96022 22248
rect 96056 21956 96068 22248
rect 96010 21602 96068 21956
rect 97068 22248 97126 22602
rect 97068 21956 97080 22248
rect 97114 21956 97126 22248
rect 97068 21602 97126 21956
rect 98126 22248 98184 22602
rect 98126 21956 98138 22248
rect 98172 21956 98184 22248
rect 98126 21602 98184 21956
rect 99184 22248 99242 22602
rect 99184 21956 99196 22248
rect 99230 21956 99242 22248
rect 99184 21602 99242 21956
rect 100242 22248 100300 22602
rect 100242 21956 100254 22248
rect 100288 21956 100300 22248
rect 100242 21602 100300 21956
rect 73852 20898 73864 21190
rect 73898 20898 73910 21190
rect 73852 20544 73910 20898
rect 75256 21164 75314 21518
rect 75256 20872 75268 21164
rect 75302 20872 75314 21164
rect 75256 20518 75314 20872
rect 76314 21164 76372 21518
rect 76314 20872 76326 21164
rect 76360 20872 76372 21164
rect 76314 20518 76372 20872
rect 77372 21164 77430 21518
rect 77372 20872 77384 21164
rect 77418 20872 77430 21164
rect 77372 20518 77430 20872
rect 78430 21164 78488 21518
rect 78430 20872 78442 21164
rect 78476 20872 78488 21164
rect 78430 20518 78488 20872
rect 79488 21164 79546 21518
rect 79488 20872 79500 21164
rect 79534 20872 79546 21164
rect 79488 20518 79546 20872
rect 80546 21164 80604 21518
rect 80546 20872 80558 21164
rect 80592 20872 80604 21164
rect 80546 20518 80604 20872
rect 81718 21162 81776 21516
rect 81718 20870 81730 21162
rect 81764 20870 81776 21162
rect 81718 20516 81776 20870
rect 82776 21162 82834 21516
rect 82776 20870 82788 21162
rect 82822 20870 82834 21162
rect 82776 20516 82834 20870
rect 83834 21162 83892 21516
rect 83834 20870 83846 21162
rect 83880 20870 83892 21162
rect 83834 20516 83892 20870
rect 84892 21162 84950 21516
rect 84892 20870 84904 21162
rect 84938 20870 84950 21162
rect 84892 20516 84950 20870
rect 85950 21162 86008 21516
rect 85950 20870 85962 21162
rect 85996 20870 86008 21162
rect 85950 20516 86008 20870
rect 87008 21162 87066 21516
rect 87008 20870 87020 21162
rect 87054 20870 87066 21162
rect 87008 20516 87066 20870
rect 88490 21156 88548 21510
rect 88490 20864 88502 21156
rect 88536 20864 88548 21156
rect 88490 20510 88548 20864
rect 89548 21156 89606 21510
rect 89548 20864 89560 21156
rect 89594 20864 89606 21156
rect 89548 20510 89606 20864
rect 90606 21156 90664 21510
rect 90606 20864 90618 21156
rect 90652 20864 90664 21156
rect 90606 20510 90664 20864
rect 91664 21156 91722 21510
rect 91664 20864 91676 21156
rect 91710 20864 91722 21156
rect 91664 20510 91722 20864
rect 92722 21156 92780 21510
rect 92722 20864 92734 21156
rect 92768 20864 92780 21156
rect 92722 20510 92780 20864
rect 93780 21156 93838 21510
rect 93780 20864 93792 21156
rect 93826 20864 93838 21156
rect 93780 20510 93838 20864
rect 94952 21154 95010 21508
rect 94952 20862 94964 21154
rect 94998 20862 95010 21154
rect 94952 20508 95010 20862
rect 96010 21154 96068 21508
rect 96010 20862 96022 21154
rect 96056 20862 96068 21154
rect 96010 20508 96068 20862
rect 97068 21154 97126 21508
rect 97068 20862 97080 21154
rect 97114 20862 97126 21154
rect 97068 20508 97126 20862
rect 98126 21154 98184 21508
rect 98126 20862 98138 21154
rect 98172 20862 98184 21154
rect 98126 20508 98184 20862
rect 99184 21154 99242 21508
rect 99184 20862 99196 21154
rect 99230 20862 99242 21154
rect 99184 20508 99242 20862
rect 100242 21154 100300 21508
rect 100242 20862 100254 21154
rect 100288 20862 100300 21154
rect 100242 20508 100300 20862
rect 62106 19730 62164 20084
rect 62106 19438 62118 19730
rect 62152 19438 62164 19730
rect 62106 19084 62164 19438
rect 63164 19730 63222 20084
rect 63164 19438 63176 19730
rect 63210 19438 63222 19730
rect 63164 19084 63222 19438
rect 64222 19730 64280 20084
rect 64222 19438 64234 19730
rect 64268 19438 64280 19730
rect 64222 19084 64280 19438
rect 65280 19730 65338 20084
rect 65280 19438 65292 19730
rect 65326 19438 65338 19730
rect 65280 19084 65338 19438
rect 66338 19730 66396 20084
rect 66338 19438 66350 19730
rect 66384 19438 66396 19730
rect 66338 19084 66396 19438
rect 67396 19730 67454 20084
rect 67396 19438 67408 19730
rect 67442 19438 67454 19730
rect 67396 19084 67454 19438
rect 68570 19742 68628 20096
rect 68570 19450 68582 19742
rect 68616 19450 68628 19742
rect 68570 19096 68628 19450
rect 69628 19742 69686 20096
rect 69628 19450 69640 19742
rect 69674 19450 69686 19742
rect 69628 19096 69686 19450
rect 70686 19742 70744 20096
rect 70686 19450 70698 19742
rect 70732 19450 70744 19742
rect 70686 19096 70744 19450
rect 71744 19742 71802 20096
rect 71744 19450 71756 19742
rect 71790 19450 71802 19742
rect 71744 19096 71802 19450
rect 72802 19742 72860 20096
rect 72802 19450 72814 19742
rect 72848 19450 72860 19742
rect 72802 19096 72860 19450
rect 73860 19742 73918 20096
rect 73860 19450 73872 19742
rect 73906 19450 73918 19742
rect 73860 19096 73918 19450
rect 75262 19702 75320 20056
rect 75262 19410 75274 19702
rect 75308 19410 75320 19702
rect 75262 19056 75320 19410
rect 76320 19702 76378 20056
rect 76320 19410 76332 19702
rect 76366 19410 76378 19702
rect 76320 19056 76378 19410
rect 77378 19702 77436 20056
rect 77378 19410 77390 19702
rect 77424 19410 77436 19702
rect 77378 19056 77436 19410
rect 78436 19702 78494 20056
rect 78436 19410 78448 19702
rect 78482 19410 78494 19702
rect 78436 19056 78494 19410
rect 79494 19702 79552 20056
rect 79494 19410 79506 19702
rect 79540 19410 79552 19702
rect 79494 19056 79552 19410
rect 80552 19702 80610 20056
rect 80552 19410 80564 19702
rect 80598 19410 80610 19702
rect 80552 19056 80610 19410
rect 81726 19714 81784 20068
rect 81726 19422 81738 19714
rect 81772 19422 81784 19714
rect 81726 19068 81784 19422
rect 82784 19714 82842 20068
rect 82784 19422 82796 19714
rect 82830 19422 82842 19714
rect 82784 19068 82842 19422
rect 83842 19714 83900 20068
rect 83842 19422 83854 19714
rect 83888 19422 83900 19714
rect 83842 19068 83900 19422
rect 84900 19714 84958 20068
rect 84900 19422 84912 19714
rect 84946 19422 84958 19714
rect 84900 19068 84958 19422
rect 85958 19714 86016 20068
rect 85958 19422 85970 19714
rect 86004 19422 86016 19714
rect 85958 19068 86016 19422
rect 87016 19714 87074 20068
rect 87016 19422 87028 19714
rect 87062 19422 87074 19714
rect 87016 19068 87074 19422
rect 88496 19694 88554 20048
rect 88496 19402 88508 19694
rect 88542 19402 88554 19694
rect 88496 19048 88554 19402
rect 89554 19694 89612 20048
rect 89554 19402 89566 19694
rect 89600 19402 89612 19694
rect 89554 19048 89612 19402
rect 90612 19694 90670 20048
rect 90612 19402 90624 19694
rect 90658 19402 90670 19694
rect 90612 19048 90670 19402
rect 91670 19694 91728 20048
rect 91670 19402 91682 19694
rect 91716 19402 91728 19694
rect 91670 19048 91728 19402
rect 92728 19694 92786 20048
rect 92728 19402 92740 19694
rect 92774 19402 92786 19694
rect 92728 19048 92786 19402
rect 93786 19694 93844 20048
rect 93786 19402 93798 19694
rect 93832 19402 93844 19694
rect 93786 19048 93844 19402
rect 94960 19706 95018 20060
rect 94960 19414 94972 19706
rect 95006 19414 95018 19706
rect 94960 19060 95018 19414
rect 96018 19706 96076 20060
rect 96018 19414 96030 19706
rect 96064 19414 96076 19706
rect 96018 19060 96076 19414
rect 97076 19706 97134 20060
rect 97076 19414 97088 19706
rect 97122 19414 97134 19706
rect 97076 19060 97134 19414
rect 98134 19706 98192 20060
rect 98134 19414 98146 19706
rect 98180 19414 98192 19706
rect 98134 19060 98192 19414
rect 99192 19706 99250 20060
rect 99192 19414 99204 19706
rect 99238 19414 99250 19706
rect 99192 19060 99250 19414
rect 100250 19706 100308 20060
rect 100250 19414 100262 19706
rect 100296 19414 100308 19706
rect 100250 19060 100308 19414
rect 62106 18636 62164 18990
rect 62106 18344 62118 18636
rect 62152 18344 62164 18636
rect 62106 17990 62164 18344
rect 63164 18636 63222 18990
rect 63164 18344 63176 18636
rect 63210 18344 63222 18636
rect 63164 17990 63222 18344
rect 64222 18636 64280 18990
rect 64222 18344 64234 18636
rect 64268 18344 64280 18636
rect 64222 17990 64280 18344
rect 65280 18636 65338 18990
rect 65280 18344 65292 18636
rect 65326 18344 65338 18636
rect 65280 17990 65338 18344
rect 66338 18636 66396 18990
rect 66338 18344 66350 18636
rect 66384 18344 66396 18636
rect 66338 17990 66396 18344
rect 67396 18636 67454 18990
rect 67396 18344 67408 18636
rect 67442 18344 67454 18636
rect 68570 18648 68628 19002
rect 67396 17990 67454 18344
rect 62106 17542 62164 17896
rect 62106 17250 62118 17542
rect 62152 17250 62164 17542
rect 62106 16896 62164 17250
rect 63164 17542 63222 17896
rect 63164 17250 63176 17542
rect 63210 17250 63222 17542
rect 63164 16896 63222 17250
rect 64222 17542 64280 17896
rect 64222 17250 64234 17542
rect 64268 17250 64280 17542
rect 64222 16896 64280 17250
rect 65280 17542 65338 17896
rect 65280 17250 65292 17542
rect 65326 17250 65338 17542
rect 65280 16896 65338 17250
rect 66338 17542 66396 17896
rect 66338 17250 66350 17542
rect 66384 17250 66396 17542
rect 66338 16896 66396 17250
rect 67396 17542 67454 17896
rect 67396 17250 67408 17542
rect 67442 17250 67454 17542
rect 67396 16896 67454 17250
rect 68570 18356 68582 18648
rect 68616 18356 68628 18648
rect 68570 18002 68628 18356
rect 69628 18648 69686 19002
rect 69628 18356 69640 18648
rect 69674 18356 69686 18648
rect 69628 18002 69686 18356
rect 70686 18648 70744 19002
rect 70686 18356 70698 18648
rect 70732 18356 70744 18648
rect 70686 18002 70744 18356
rect 71744 18648 71802 19002
rect 71744 18356 71756 18648
rect 71790 18356 71802 18648
rect 71744 18002 71802 18356
rect 72802 18648 72860 19002
rect 72802 18356 72814 18648
rect 72848 18356 72860 18648
rect 72802 18002 72860 18356
rect 73860 18648 73918 19002
rect 73860 18356 73872 18648
rect 73906 18356 73918 18648
rect 73860 18002 73918 18356
rect 75262 18608 75320 18962
rect 62106 16448 62164 16802
rect 62106 16156 62118 16448
rect 62152 16156 62164 16448
rect 62106 15802 62164 16156
rect 63164 16448 63222 16802
rect 63164 16156 63176 16448
rect 63210 16156 63222 16448
rect 63164 15802 63222 16156
rect 64222 16448 64280 16802
rect 64222 16156 64234 16448
rect 64268 16156 64280 16448
rect 64222 15802 64280 16156
rect 65280 16448 65338 16802
rect 65280 16156 65292 16448
rect 65326 16156 65338 16448
rect 65280 15802 65338 16156
rect 66338 16448 66396 16802
rect 66338 16156 66350 16448
rect 66384 16156 66396 16448
rect 66338 15802 66396 16156
rect 67396 16448 67454 16802
rect 68570 17554 68628 17908
rect 68570 17262 68582 17554
rect 68616 17262 68628 17554
rect 68570 16908 68628 17262
rect 69628 17554 69686 17908
rect 69628 17262 69640 17554
rect 69674 17262 69686 17554
rect 69628 16908 69686 17262
rect 70686 17554 70744 17908
rect 70686 17262 70698 17554
rect 70732 17262 70744 17554
rect 70686 16908 70744 17262
rect 71744 17554 71802 17908
rect 71744 17262 71756 17554
rect 71790 17262 71802 17554
rect 71744 16908 71802 17262
rect 72802 17554 72860 17908
rect 72802 17262 72814 17554
rect 72848 17262 72860 17554
rect 72802 16908 72860 17262
rect 73860 17554 73918 17908
rect 73860 17262 73872 17554
rect 73906 17262 73918 17554
rect 73860 16908 73918 17262
rect 75262 18316 75274 18608
rect 75308 18316 75320 18608
rect 75262 17962 75320 18316
rect 76320 18608 76378 18962
rect 76320 18316 76332 18608
rect 76366 18316 76378 18608
rect 76320 17962 76378 18316
rect 77378 18608 77436 18962
rect 77378 18316 77390 18608
rect 77424 18316 77436 18608
rect 77378 17962 77436 18316
rect 78436 18608 78494 18962
rect 78436 18316 78448 18608
rect 78482 18316 78494 18608
rect 78436 17962 78494 18316
rect 79494 18608 79552 18962
rect 79494 18316 79506 18608
rect 79540 18316 79552 18608
rect 79494 17962 79552 18316
rect 80552 18608 80610 18962
rect 80552 18316 80564 18608
rect 80598 18316 80610 18608
rect 81726 18620 81784 18974
rect 80552 17962 80610 18316
rect 67396 16156 67408 16448
rect 67442 16156 67454 16448
rect 67396 15802 67454 16156
rect 68570 16460 68628 16814
rect 68570 16168 68582 16460
rect 68616 16168 68628 16460
rect 68570 15814 68628 16168
rect 69628 16460 69686 16814
rect 69628 16168 69640 16460
rect 69674 16168 69686 16460
rect 69628 15814 69686 16168
rect 70686 16460 70744 16814
rect 70686 16168 70698 16460
rect 70732 16168 70744 16460
rect 70686 15814 70744 16168
rect 71744 16460 71802 16814
rect 71744 16168 71756 16460
rect 71790 16168 71802 16460
rect 71744 15814 71802 16168
rect 72802 16460 72860 16814
rect 72802 16168 72814 16460
rect 72848 16168 72860 16460
rect 72802 15814 72860 16168
rect 73860 16460 73918 16814
rect 75262 17514 75320 17868
rect 75262 17222 75274 17514
rect 75308 17222 75320 17514
rect 75262 16868 75320 17222
rect 76320 17514 76378 17868
rect 76320 17222 76332 17514
rect 76366 17222 76378 17514
rect 76320 16868 76378 17222
rect 77378 17514 77436 17868
rect 77378 17222 77390 17514
rect 77424 17222 77436 17514
rect 77378 16868 77436 17222
rect 78436 17514 78494 17868
rect 78436 17222 78448 17514
rect 78482 17222 78494 17514
rect 78436 16868 78494 17222
rect 79494 17514 79552 17868
rect 79494 17222 79506 17514
rect 79540 17222 79552 17514
rect 79494 16868 79552 17222
rect 80552 17514 80610 17868
rect 80552 17222 80564 17514
rect 80598 17222 80610 17514
rect 80552 16868 80610 17222
rect 81726 18328 81738 18620
rect 81772 18328 81784 18620
rect 81726 17974 81784 18328
rect 82784 18620 82842 18974
rect 82784 18328 82796 18620
rect 82830 18328 82842 18620
rect 82784 17974 82842 18328
rect 83842 18620 83900 18974
rect 83842 18328 83854 18620
rect 83888 18328 83900 18620
rect 83842 17974 83900 18328
rect 84900 18620 84958 18974
rect 84900 18328 84912 18620
rect 84946 18328 84958 18620
rect 84900 17974 84958 18328
rect 85958 18620 86016 18974
rect 85958 18328 85970 18620
rect 86004 18328 86016 18620
rect 85958 17974 86016 18328
rect 87016 18620 87074 18974
rect 87016 18328 87028 18620
rect 87062 18328 87074 18620
rect 87016 17974 87074 18328
rect 88496 18600 88554 18954
rect 73860 16168 73872 16460
rect 73906 16168 73918 16460
rect 73860 15814 73918 16168
rect 75262 16420 75320 16774
rect 75262 16128 75274 16420
rect 75308 16128 75320 16420
rect 75262 15774 75320 16128
rect 76320 16420 76378 16774
rect 76320 16128 76332 16420
rect 76366 16128 76378 16420
rect 76320 15774 76378 16128
rect 77378 16420 77436 16774
rect 77378 16128 77390 16420
rect 77424 16128 77436 16420
rect 77378 15774 77436 16128
rect 78436 16420 78494 16774
rect 78436 16128 78448 16420
rect 78482 16128 78494 16420
rect 78436 15774 78494 16128
rect 79494 16420 79552 16774
rect 79494 16128 79506 16420
rect 79540 16128 79552 16420
rect 79494 15774 79552 16128
rect 80552 16420 80610 16774
rect 81726 17526 81784 17880
rect 81726 17234 81738 17526
rect 81772 17234 81784 17526
rect 81726 16880 81784 17234
rect 82784 17526 82842 17880
rect 82784 17234 82796 17526
rect 82830 17234 82842 17526
rect 82784 16880 82842 17234
rect 83842 17526 83900 17880
rect 83842 17234 83854 17526
rect 83888 17234 83900 17526
rect 83842 16880 83900 17234
rect 84900 17526 84958 17880
rect 84900 17234 84912 17526
rect 84946 17234 84958 17526
rect 84900 16880 84958 17234
rect 85958 17526 86016 17880
rect 85958 17234 85970 17526
rect 86004 17234 86016 17526
rect 85958 16880 86016 17234
rect 87016 17526 87074 17880
rect 87016 17234 87028 17526
rect 87062 17234 87074 17526
rect 87016 16880 87074 17234
rect 88496 18308 88508 18600
rect 88542 18308 88554 18600
rect 88496 17954 88554 18308
rect 89554 18600 89612 18954
rect 89554 18308 89566 18600
rect 89600 18308 89612 18600
rect 89554 17954 89612 18308
rect 90612 18600 90670 18954
rect 90612 18308 90624 18600
rect 90658 18308 90670 18600
rect 90612 17954 90670 18308
rect 91670 18600 91728 18954
rect 91670 18308 91682 18600
rect 91716 18308 91728 18600
rect 91670 17954 91728 18308
rect 92728 18600 92786 18954
rect 92728 18308 92740 18600
rect 92774 18308 92786 18600
rect 92728 17954 92786 18308
rect 93786 18600 93844 18954
rect 93786 18308 93798 18600
rect 93832 18308 93844 18600
rect 94960 18612 95018 18966
rect 93786 17954 93844 18308
rect 80552 16128 80564 16420
rect 80598 16128 80610 16420
rect 80552 15774 80610 16128
rect 81726 16432 81784 16786
rect 81726 16140 81738 16432
rect 81772 16140 81784 16432
rect 81726 15786 81784 16140
rect 82784 16432 82842 16786
rect 82784 16140 82796 16432
rect 82830 16140 82842 16432
rect 82784 15786 82842 16140
rect 83842 16432 83900 16786
rect 83842 16140 83854 16432
rect 83888 16140 83900 16432
rect 83842 15786 83900 16140
rect 84900 16432 84958 16786
rect 84900 16140 84912 16432
rect 84946 16140 84958 16432
rect 84900 15786 84958 16140
rect 85958 16432 86016 16786
rect 85958 16140 85970 16432
rect 86004 16140 86016 16432
rect 85958 15786 86016 16140
rect 87016 16432 87074 16786
rect 88496 17506 88554 17860
rect 88496 17214 88508 17506
rect 88542 17214 88554 17506
rect 88496 16860 88554 17214
rect 89554 17506 89612 17860
rect 89554 17214 89566 17506
rect 89600 17214 89612 17506
rect 89554 16860 89612 17214
rect 90612 17506 90670 17860
rect 90612 17214 90624 17506
rect 90658 17214 90670 17506
rect 90612 16860 90670 17214
rect 91670 17506 91728 17860
rect 91670 17214 91682 17506
rect 91716 17214 91728 17506
rect 91670 16860 91728 17214
rect 92728 17506 92786 17860
rect 92728 17214 92740 17506
rect 92774 17214 92786 17506
rect 92728 16860 92786 17214
rect 93786 17506 93844 17860
rect 93786 17214 93798 17506
rect 93832 17214 93844 17506
rect 93786 16860 93844 17214
rect 94960 18320 94972 18612
rect 95006 18320 95018 18612
rect 94960 17966 95018 18320
rect 96018 18612 96076 18966
rect 96018 18320 96030 18612
rect 96064 18320 96076 18612
rect 96018 17966 96076 18320
rect 97076 18612 97134 18966
rect 97076 18320 97088 18612
rect 97122 18320 97134 18612
rect 97076 17966 97134 18320
rect 98134 18612 98192 18966
rect 98134 18320 98146 18612
rect 98180 18320 98192 18612
rect 98134 17966 98192 18320
rect 99192 18612 99250 18966
rect 99192 18320 99204 18612
rect 99238 18320 99250 18612
rect 99192 17966 99250 18320
rect 100250 18612 100308 18966
rect 100250 18320 100262 18612
rect 100296 18320 100308 18612
rect 100250 17966 100308 18320
rect 87016 16140 87028 16432
rect 87062 16140 87074 16432
rect 87016 15786 87074 16140
rect 88496 16412 88554 16766
rect 88496 16120 88508 16412
rect 88542 16120 88554 16412
rect 88496 15766 88554 16120
rect 89554 16412 89612 16766
rect 89554 16120 89566 16412
rect 89600 16120 89612 16412
rect 89554 15766 89612 16120
rect 90612 16412 90670 16766
rect 90612 16120 90624 16412
rect 90658 16120 90670 16412
rect 90612 15766 90670 16120
rect 91670 16412 91728 16766
rect 91670 16120 91682 16412
rect 91716 16120 91728 16412
rect 91670 15766 91728 16120
rect 92728 16412 92786 16766
rect 92728 16120 92740 16412
rect 92774 16120 92786 16412
rect 92728 15766 92786 16120
rect 93786 16412 93844 16766
rect 94960 17518 95018 17872
rect 94960 17226 94972 17518
rect 95006 17226 95018 17518
rect 94960 16872 95018 17226
rect 96018 17518 96076 17872
rect 96018 17226 96030 17518
rect 96064 17226 96076 17518
rect 96018 16872 96076 17226
rect 97076 17518 97134 17872
rect 97076 17226 97088 17518
rect 97122 17226 97134 17518
rect 97076 16872 97134 17226
rect 98134 17518 98192 17872
rect 98134 17226 98146 17518
rect 98180 17226 98192 17518
rect 98134 16872 98192 17226
rect 99192 17518 99250 17872
rect 99192 17226 99204 17518
rect 99238 17226 99250 17518
rect 99192 16872 99250 17226
rect 100250 17518 100308 17872
rect 100250 17226 100262 17518
rect 100296 17226 100308 17518
rect 100250 16872 100308 17226
rect 93786 16120 93798 16412
rect 93832 16120 93844 16412
rect 93786 15766 93844 16120
rect 94960 16424 95018 16778
rect 94960 16132 94972 16424
rect 95006 16132 95018 16424
rect 94960 15778 95018 16132
rect 96018 16424 96076 16778
rect 96018 16132 96030 16424
rect 96064 16132 96076 16424
rect 96018 15778 96076 16132
rect 97076 16424 97134 16778
rect 97076 16132 97088 16424
rect 97122 16132 97134 16424
rect 97076 15778 97134 16132
rect 98134 16424 98192 16778
rect 98134 16132 98146 16424
rect 98180 16132 98192 16424
rect 98134 15778 98192 16132
rect 99192 16424 99250 16778
rect 99192 16132 99204 16424
rect 99238 16132 99250 16424
rect 99192 15778 99250 16132
rect 100250 16424 100308 16778
rect 100250 16132 100262 16424
rect 100296 16132 100308 16424
rect 100250 15778 100308 16132
rect 62106 15354 62164 15708
rect 62106 15062 62118 15354
rect 62152 15062 62164 15354
rect 62106 14708 62164 15062
rect 63164 15354 63222 15708
rect 63164 15062 63176 15354
rect 63210 15062 63222 15354
rect 63164 14708 63222 15062
rect 64222 15354 64280 15708
rect 64222 15062 64234 15354
rect 64268 15062 64280 15354
rect 64222 14708 64280 15062
rect 65280 15354 65338 15708
rect 65280 15062 65292 15354
rect 65326 15062 65338 15354
rect 65280 14708 65338 15062
rect 66338 15354 66396 15708
rect 66338 15062 66350 15354
rect 66384 15062 66396 15354
rect 66338 14708 66396 15062
rect 67396 15354 67454 15708
rect 67396 15062 67408 15354
rect 67442 15062 67454 15354
rect 67396 14708 67454 15062
rect 68570 15366 68628 15720
rect 68570 15074 68582 15366
rect 68616 15074 68628 15366
rect 68570 14720 68628 15074
rect 69628 15366 69686 15720
rect 69628 15074 69640 15366
rect 69674 15074 69686 15366
rect 69628 14720 69686 15074
rect 70686 15366 70744 15720
rect 70686 15074 70698 15366
rect 70732 15074 70744 15366
rect 70686 14720 70744 15074
rect 71744 15366 71802 15720
rect 71744 15074 71756 15366
rect 71790 15074 71802 15366
rect 71744 14720 71802 15074
rect 72802 15366 72860 15720
rect 72802 15074 72814 15366
rect 72848 15074 72860 15366
rect 72802 14720 72860 15074
rect 73860 15366 73918 15720
rect 73860 15074 73872 15366
rect 73906 15074 73918 15366
rect 73860 14720 73918 15074
rect 75262 15326 75320 15680
rect 75262 15034 75274 15326
rect 75308 15034 75320 15326
rect 75262 14680 75320 15034
rect 76320 15326 76378 15680
rect 76320 15034 76332 15326
rect 76366 15034 76378 15326
rect 76320 14680 76378 15034
rect 77378 15326 77436 15680
rect 77378 15034 77390 15326
rect 77424 15034 77436 15326
rect 77378 14680 77436 15034
rect 78436 15326 78494 15680
rect 78436 15034 78448 15326
rect 78482 15034 78494 15326
rect 78436 14680 78494 15034
rect 79494 15326 79552 15680
rect 79494 15034 79506 15326
rect 79540 15034 79552 15326
rect 79494 14680 79552 15034
rect 80552 15326 80610 15680
rect 80552 15034 80564 15326
rect 80598 15034 80610 15326
rect 80552 14680 80610 15034
rect 81726 15338 81784 15692
rect 81726 15046 81738 15338
rect 81772 15046 81784 15338
rect 81726 14692 81784 15046
rect 82784 15338 82842 15692
rect 82784 15046 82796 15338
rect 82830 15046 82842 15338
rect 82784 14692 82842 15046
rect 83842 15338 83900 15692
rect 83842 15046 83854 15338
rect 83888 15046 83900 15338
rect 83842 14692 83900 15046
rect 84900 15338 84958 15692
rect 84900 15046 84912 15338
rect 84946 15046 84958 15338
rect 84900 14692 84958 15046
rect 85958 15338 86016 15692
rect 85958 15046 85970 15338
rect 86004 15046 86016 15338
rect 85958 14692 86016 15046
rect 87016 15338 87074 15692
rect 87016 15046 87028 15338
rect 87062 15046 87074 15338
rect 87016 14692 87074 15046
rect 88496 15318 88554 15672
rect 88496 15026 88508 15318
rect 88542 15026 88554 15318
rect 88496 14672 88554 15026
rect 89554 15318 89612 15672
rect 89554 15026 89566 15318
rect 89600 15026 89612 15318
rect 89554 14672 89612 15026
rect 90612 15318 90670 15672
rect 90612 15026 90624 15318
rect 90658 15026 90670 15318
rect 90612 14672 90670 15026
rect 91670 15318 91728 15672
rect 91670 15026 91682 15318
rect 91716 15026 91728 15318
rect 91670 14672 91728 15026
rect 92728 15318 92786 15672
rect 92728 15026 92740 15318
rect 92774 15026 92786 15318
rect 92728 14672 92786 15026
rect 93786 15318 93844 15672
rect 93786 15026 93798 15318
rect 93832 15026 93844 15318
rect 93786 14672 93844 15026
rect 94960 15330 95018 15684
rect 94960 15038 94972 15330
rect 95006 15038 95018 15330
rect 94960 14684 95018 15038
rect 96018 15330 96076 15684
rect 96018 15038 96030 15330
rect 96064 15038 96076 15330
rect 96018 14684 96076 15038
rect 97076 15330 97134 15684
rect 97076 15038 97088 15330
rect 97122 15038 97134 15330
rect 97076 14684 97134 15038
rect 98134 15330 98192 15684
rect 98134 15038 98146 15330
rect 98180 15038 98192 15330
rect 98134 14684 98192 15038
rect 99192 15330 99250 15684
rect 99192 15038 99204 15330
rect 99238 15038 99250 15330
rect 99192 14684 99250 15038
rect 100250 15330 100308 15684
rect 100250 15038 100262 15330
rect 100296 15038 100308 15330
rect 100250 14684 100308 15038
rect 62106 13872 62164 14226
rect 62106 13580 62118 13872
rect 62152 13580 62164 13872
rect 62106 13226 62164 13580
rect 63164 13872 63222 14226
rect 63164 13580 63176 13872
rect 63210 13580 63222 13872
rect 63164 13226 63222 13580
rect 64222 13872 64280 14226
rect 64222 13580 64234 13872
rect 64268 13580 64280 13872
rect 64222 13226 64280 13580
rect 65280 13872 65338 14226
rect 65280 13580 65292 13872
rect 65326 13580 65338 13872
rect 65280 13226 65338 13580
rect 66338 13872 66396 14226
rect 66338 13580 66350 13872
rect 66384 13580 66396 13872
rect 66338 13226 66396 13580
rect 67396 13872 67454 14226
rect 67396 13580 67408 13872
rect 67442 13580 67454 13872
rect 67396 13226 67454 13580
rect 68574 13870 68632 14224
rect 68574 13578 68586 13870
rect 68620 13578 68632 13870
rect 68574 13224 68632 13578
rect 69632 13870 69690 14224
rect 69632 13578 69644 13870
rect 69678 13578 69690 13870
rect 69632 13224 69690 13578
rect 70690 13870 70748 14224
rect 70690 13578 70702 13870
rect 70736 13578 70748 13870
rect 70690 13224 70748 13578
rect 71748 13870 71806 14224
rect 71748 13578 71760 13870
rect 71794 13578 71806 13870
rect 71748 13224 71806 13578
rect 72806 13870 72864 14224
rect 72806 13578 72818 13870
rect 72852 13578 72864 13870
rect 72806 13224 72864 13578
rect 73864 13870 73922 14224
rect 73864 13578 73876 13870
rect 73910 13578 73922 13870
rect 73864 13224 73922 13578
rect 75262 13844 75320 14198
rect 75262 13552 75274 13844
rect 75308 13552 75320 13844
rect 75262 13198 75320 13552
rect 76320 13844 76378 14198
rect 76320 13552 76332 13844
rect 76366 13552 76378 13844
rect 76320 13198 76378 13552
rect 77378 13844 77436 14198
rect 77378 13552 77390 13844
rect 77424 13552 77436 13844
rect 77378 13198 77436 13552
rect 78436 13844 78494 14198
rect 78436 13552 78448 13844
rect 78482 13552 78494 13844
rect 78436 13198 78494 13552
rect 79494 13844 79552 14198
rect 79494 13552 79506 13844
rect 79540 13552 79552 13844
rect 79494 13198 79552 13552
rect 80552 13844 80610 14198
rect 80552 13552 80564 13844
rect 80598 13552 80610 13844
rect 80552 13198 80610 13552
rect 81730 13842 81788 14196
rect 81730 13550 81742 13842
rect 81776 13550 81788 13842
rect 81730 13196 81788 13550
rect 82788 13842 82846 14196
rect 82788 13550 82800 13842
rect 82834 13550 82846 13842
rect 82788 13196 82846 13550
rect 83846 13842 83904 14196
rect 83846 13550 83858 13842
rect 83892 13550 83904 13842
rect 83846 13196 83904 13550
rect 84904 13842 84962 14196
rect 84904 13550 84916 13842
rect 84950 13550 84962 13842
rect 84904 13196 84962 13550
rect 85962 13842 86020 14196
rect 85962 13550 85974 13842
rect 86008 13550 86020 13842
rect 85962 13196 86020 13550
rect 87020 13842 87078 14196
rect 87020 13550 87032 13842
rect 87066 13550 87078 13842
rect 87020 13196 87078 13550
rect 88496 13836 88554 14190
rect 88496 13544 88508 13836
rect 88542 13544 88554 13836
rect 62106 12778 62164 13132
rect 62106 12486 62118 12778
rect 62152 12486 62164 12778
rect 62106 12132 62164 12486
rect 63164 12778 63222 13132
rect 63164 12486 63176 12778
rect 63210 12486 63222 12778
rect 63164 12132 63222 12486
rect 64222 12778 64280 13132
rect 64222 12486 64234 12778
rect 64268 12486 64280 12778
rect 64222 12132 64280 12486
rect 65280 12778 65338 13132
rect 65280 12486 65292 12778
rect 65326 12486 65338 12778
rect 65280 12132 65338 12486
rect 66338 12778 66396 13132
rect 66338 12486 66350 12778
rect 66384 12486 66396 12778
rect 66338 12132 66396 12486
rect 67396 12778 67454 13132
rect 88496 13190 88554 13544
rect 89554 13836 89612 14190
rect 89554 13544 89566 13836
rect 89600 13544 89612 13836
rect 89554 13190 89612 13544
rect 90612 13836 90670 14190
rect 90612 13544 90624 13836
rect 90658 13544 90670 13836
rect 90612 13190 90670 13544
rect 91670 13836 91728 14190
rect 91670 13544 91682 13836
rect 91716 13544 91728 13836
rect 91670 13190 91728 13544
rect 92728 13836 92786 14190
rect 92728 13544 92740 13836
rect 92774 13544 92786 13836
rect 92728 13190 92786 13544
rect 93786 13836 93844 14190
rect 93786 13544 93798 13836
rect 93832 13544 93844 13836
rect 93786 13190 93844 13544
rect 94964 13834 95022 14188
rect 94964 13542 94976 13834
rect 95010 13542 95022 13834
rect 67396 12486 67408 12778
rect 67442 12486 67454 12778
rect 68574 12776 68632 13130
rect 67396 12132 67454 12486
rect 62106 11684 62164 12038
rect 62106 11392 62118 11684
rect 62152 11392 62164 11684
rect 62106 11038 62164 11392
rect 63164 11684 63222 12038
rect 63164 11392 63176 11684
rect 63210 11392 63222 11684
rect 63164 11038 63222 11392
rect 64222 11684 64280 12038
rect 64222 11392 64234 11684
rect 64268 11392 64280 11684
rect 64222 11038 64280 11392
rect 65280 11684 65338 12038
rect 65280 11392 65292 11684
rect 65326 11392 65338 11684
rect 65280 11038 65338 11392
rect 66338 11684 66396 12038
rect 66338 11392 66350 11684
rect 66384 11392 66396 11684
rect 66338 11038 66396 11392
rect 67396 11684 67454 12038
rect 67396 11392 67408 11684
rect 67442 11392 67454 11684
rect 67396 11038 67454 11392
rect 68574 12484 68586 12776
rect 68620 12484 68632 12776
rect 68574 12130 68632 12484
rect 69632 12776 69690 13130
rect 69632 12484 69644 12776
rect 69678 12484 69690 12776
rect 69632 12130 69690 12484
rect 70690 12776 70748 13130
rect 70690 12484 70702 12776
rect 70736 12484 70748 12776
rect 70690 12130 70748 12484
rect 71748 12776 71806 13130
rect 71748 12484 71760 12776
rect 71794 12484 71806 12776
rect 71748 12130 71806 12484
rect 72806 12776 72864 13130
rect 72806 12484 72818 12776
rect 72852 12484 72864 12776
rect 72806 12130 72864 12484
rect 73864 12776 73922 13130
rect 94964 13188 95022 13542
rect 96022 13834 96080 14188
rect 96022 13542 96034 13834
rect 96068 13542 96080 13834
rect 96022 13188 96080 13542
rect 97080 13834 97138 14188
rect 97080 13542 97092 13834
rect 97126 13542 97138 13834
rect 97080 13188 97138 13542
rect 98138 13834 98196 14188
rect 98138 13542 98150 13834
rect 98184 13542 98196 13834
rect 98138 13188 98196 13542
rect 99196 13834 99254 14188
rect 99196 13542 99208 13834
rect 99242 13542 99254 13834
rect 99196 13188 99254 13542
rect 100254 13834 100312 14188
rect 100254 13542 100266 13834
rect 100300 13542 100312 13834
rect 100254 13188 100312 13542
rect 73864 12484 73876 12776
rect 73910 12484 73922 12776
rect 73864 12130 73922 12484
rect 75262 12750 75320 13104
rect 62106 10590 62164 10944
rect 62106 10298 62118 10590
rect 62152 10298 62164 10590
rect 62106 9944 62164 10298
rect 63164 10590 63222 10944
rect 63164 10298 63176 10590
rect 63210 10298 63222 10590
rect 63164 9944 63222 10298
rect 64222 10590 64280 10944
rect 64222 10298 64234 10590
rect 64268 10298 64280 10590
rect 64222 9944 64280 10298
rect 65280 10590 65338 10944
rect 65280 10298 65292 10590
rect 65326 10298 65338 10590
rect 65280 9944 65338 10298
rect 66338 10590 66396 10944
rect 66338 10298 66350 10590
rect 66384 10298 66396 10590
rect 66338 9944 66396 10298
rect 67396 10590 67454 10944
rect 68574 11682 68632 12036
rect 68574 11390 68586 11682
rect 68620 11390 68632 11682
rect 68574 11036 68632 11390
rect 69632 11682 69690 12036
rect 69632 11390 69644 11682
rect 69678 11390 69690 11682
rect 69632 11036 69690 11390
rect 70690 11682 70748 12036
rect 70690 11390 70702 11682
rect 70736 11390 70748 11682
rect 70690 11036 70748 11390
rect 71748 11682 71806 12036
rect 71748 11390 71760 11682
rect 71794 11390 71806 11682
rect 71748 11036 71806 11390
rect 72806 11682 72864 12036
rect 72806 11390 72818 11682
rect 72852 11390 72864 11682
rect 72806 11036 72864 11390
rect 73864 11682 73922 12036
rect 73864 11390 73876 11682
rect 73910 11390 73922 11682
rect 73864 11036 73922 11390
rect 75262 12458 75274 12750
rect 75308 12458 75320 12750
rect 75262 12104 75320 12458
rect 76320 12750 76378 13104
rect 76320 12458 76332 12750
rect 76366 12458 76378 12750
rect 76320 12104 76378 12458
rect 77378 12750 77436 13104
rect 77378 12458 77390 12750
rect 77424 12458 77436 12750
rect 77378 12104 77436 12458
rect 78436 12750 78494 13104
rect 78436 12458 78448 12750
rect 78482 12458 78494 12750
rect 78436 12104 78494 12458
rect 79494 12750 79552 13104
rect 79494 12458 79506 12750
rect 79540 12458 79552 12750
rect 79494 12104 79552 12458
rect 80552 12750 80610 13104
rect 80552 12458 80564 12750
rect 80598 12458 80610 12750
rect 81730 12748 81788 13102
rect 80552 12104 80610 12458
rect 67396 10298 67408 10590
rect 67442 10298 67454 10590
rect 67396 9944 67454 10298
rect 68574 10588 68632 10942
rect 68574 10296 68586 10588
rect 68620 10296 68632 10588
rect 68574 9942 68632 10296
rect 69632 10588 69690 10942
rect 69632 10296 69644 10588
rect 69678 10296 69690 10588
rect 69632 9942 69690 10296
rect 70690 10588 70748 10942
rect 70690 10296 70702 10588
rect 70736 10296 70748 10588
rect 70690 9942 70748 10296
rect 71748 10588 71806 10942
rect 71748 10296 71760 10588
rect 71794 10296 71806 10588
rect 71748 9942 71806 10296
rect 72806 10588 72864 10942
rect 72806 10296 72818 10588
rect 72852 10296 72864 10588
rect 72806 9942 72864 10296
rect 73864 10588 73922 10942
rect 75262 11656 75320 12010
rect 75262 11364 75274 11656
rect 75308 11364 75320 11656
rect 75262 11010 75320 11364
rect 76320 11656 76378 12010
rect 76320 11364 76332 11656
rect 76366 11364 76378 11656
rect 76320 11010 76378 11364
rect 77378 11656 77436 12010
rect 77378 11364 77390 11656
rect 77424 11364 77436 11656
rect 77378 11010 77436 11364
rect 78436 11656 78494 12010
rect 78436 11364 78448 11656
rect 78482 11364 78494 11656
rect 78436 11010 78494 11364
rect 79494 11656 79552 12010
rect 79494 11364 79506 11656
rect 79540 11364 79552 11656
rect 79494 11010 79552 11364
rect 80552 11656 80610 12010
rect 80552 11364 80564 11656
rect 80598 11364 80610 11656
rect 80552 11010 80610 11364
rect 81730 12456 81742 12748
rect 81776 12456 81788 12748
rect 81730 12102 81788 12456
rect 82788 12748 82846 13102
rect 82788 12456 82800 12748
rect 82834 12456 82846 12748
rect 82788 12102 82846 12456
rect 83846 12748 83904 13102
rect 83846 12456 83858 12748
rect 83892 12456 83904 12748
rect 83846 12102 83904 12456
rect 84904 12748 84962 13102
rect 84904 12456 84916 12748
rect 84950 12456 84962 12748
rect 84904 12102 84962 12456
rect 85962 12748 86020 13102
rect 85962 12456 85974 12748
rect 86008 12456 86020 12748
rect 85962 12102 86020 12456
rect 87020 12748 87078 13102
rect 87020 12456 87032 12748
rect 87066 12456 87078 12748
rect 88496 12742 88554 13096
rect 87020 12102 87078 12456
rect 73864 10296 73876 10588
rect 73910 10296 73922 10588
rect 73864 9942 73922 10296
rect 75262 10562 75320 10916
rect 75262 10270 75274 10562
rect 75308 10270 75320 10562
rect 75262 9916 75320 10270
rect 76320 10562 76378 10916
rect 76320 10270 76332 10562
rect 76366 10270 76378 10562
rect 76320 9916 76378 10270
rect 77378 10562 77436 10916
rect 77378 10270 77390 10562
rect 77424 10270 77436 10562
rect 77378 9916 77436 10270
rect 78436 10562 78494 10916
rect 78436 10270 78448 10562
rect 78482 10270 78494 10562
rect 78436 9916 78494 10270
rect 79494 10562 79552 10916
rect 79494 10270 79506 10562
rect 79540 10270 79552 10562
rect 79494 9916 79552 10270
rect 80552 10562 80610 10916
rect 81730 11654 81788 12008
rect 81730 11362 81742 11654
rect 81776 11362 81788 11654
rect 81730 11008 81788 11362
rect 82788 11654 82846 12008
rect 82788 11362 82800 11654
rect 82834 11362 82846 11654
rect 82788 11008 82846 11362
rect 83846 11654 83904 12008
rect 83846 11362 83858 11654
rect 83892 11362 83904 11654
rect 83846 11008 83904 11362
rect 84904 11654 84962 12008
rect 84904 11362 84916 11654
rect 84950 11362 84962 11654
rect 84904 11008 84962 11362
rect 85962 11654 86020 12008
rect 85962 11362 85974 11654
rect 86008 11362 86020 11654
rect 85962 11008 86020 11362
rect 87020 11654 87078 12008
rect 87020 11362 87032 11654
rect 87066 11362 87078 11654
rect 87020 11008 87078 11362
rect 88496 12450 88508 12742
rect 88542 12450 88554 12742
rect 88496 12096 88554 12450
rect 89554 12742 89612 13096
rect 89554 12450 89566 12742
rect 89600 12450 89612 12742
rect 89554 12096 89612 12450
rect 90612 12742 90670 13096
rect 90612 12450 90624 12742
rect 90658 12450 90670 12742
rect 90612 12096 90670 12450
rect 91670 12742 91728 13096
rect 91670 12450 91682 12742
rect 91716 12450 91728 12742
rect 91670 12096 91728 12450
rect 92728 12742 92786 13096
rect 92728 12450 92740 12742
rect 92774 12450 92786 12742
rect 92728 12096 92786 12450
rect 93786 12742 93844 13096
rect 93786 12450 93798 12742
rect 93832 12450 93844 12742
rect 94964 12740 95022 13094
rect 93786 12096 93844 12450
rect 80552 10270 80564 10562
rect 80598 10270 80610 10562
rect 80552 9916 80610 10270
rect 81730 10560 81788 10914
rect 81730 10268 81742 10560
rect 81776 10268 81788 10560
rect 81730 9914 81788 10268
rect 82788 10560 82846 10914
rect 82788 10268 82800 10560
rect 82834 10268 82846 10560
rect 82788 9914 82846 10268
rect 83846 10560 83904 10914
rect 83846 10268 83858 10560
rect 83892 10268 83904 10560
rect 83846 9914 83904 10268
rect 84904 10560 84962 10914
rect 84904 10268 84916 10560
rect 84950 10268 84962 10560
rect 84904 9914 84962 10268
rect 85962 10560 86020 10914
rect 85962 10268 85974 10560
rect 86008 10268 86020 10560
rect 85962 9914 86020 10268
rect 87020 10560 87078 10914
rect 88496 11648 88554 12002
rect 88496 11356 88508 11648
rect 88542 11356 88554 11648
rect 88496 11002 88554 11356
rect 89554 11648 89612 12002
rect 89554 11356 89566 11648
rect 89600 11356 89612 11648
rect 89554 11002 89612 11356
rect 90612 11648 90670 12002
rect 90612 11356 90624 11648
rect 90658 11356 90670 11648
rect 90612 11002 90670 11356
rect 91670 11648 91728 12002
rect 91670 11356 91682 11648
rect 91716 11356 91728 11648
rect 91670 11002 91728 11356
rect 92728 11648 92786 12002
rect 92728 11356 92740 11648
rect 92774 11356 92786 11648
rect 92728 11002 92786 11356
rect 93786 11648 93844 12002
rect 93786 11356 93798 11648
rect 93832 11356 93844 11648
rect 93786 11002 93844 11356
rect 94964 12448 94976 12740
rect 95010 12448 95022 12740
rect 94964 12094 95022 12448
rect 96022 12740 96080 13094
rect 96022 12448 96034 12740
rect 96068 12448 96080 12740
rect 96022 12094 96080 12448
rect 97080 12740 97138 13094
rect 97080 12448 97092 12740
rect 97126 12448 97138 12740
rect 97080 12094 97138 12448
rect 98138 12740 98196 13094
rect 98138 12448 98150 12740
rect 98184 12448 98196 12740
rect 98138 12094 98196 12448
rect 99196 12740 99254 13094
rect 99196 12448 99208 12740
rect 99242 12448 99254 12740
rect 99196 12094 99254 12448
rect 100254 12740 100312 13094
rect 100254 12448 100266 12740
rect 100300 12448 100312 12740
rect 100254 12094 100312 12448
rect 87020 10268 87032 10560
rect 87066 10268 87078 10560
rect 87020 9914 87078 10268
rect 88496 10554 88554 10908
rect 88496 10262 88508 10554
rect 88542 10262 88554 10554
rect 62106 9496 62164 9850
rect 62106 9204 62118 9496
rect 62152 9204 62164 9496
rect 62106 8850 62164 9204
rect 63164 9496 63222 9850
rect 63164 9204 63176 9496
rect 63210 9204 63222 9496
rect 63164 8850 63222 9204
rect 64222 9496 64280 9850
rect 64222 9204 64234 9496
rect 64268 9204 64280 9496
rect 64222 8850 64280 9204
rect 65280 9496 65338 9850
rect 65280 9204 65292 9496
rect 65326 9204 65338 9496
rect 65280 8850 65338 9204
rect 66338 9496 66396 9850
rect 66338 9204 66350 9496
rect 66384 9204 66396 9496
rect 66338 8850 66396 9204
rect 67396 9496 67454 9850
rect 88496 9908 88554 10262
rect 89554 10554 89612 10908
rect 89554 10262 89566 10554
rect 89600 10262 89612 10554
rect 89554 9908 89612 10262
rect 90612 10554 90670 10908
rect 90612 10262 90624 10554
rect 90658 10262 90670 10554
rect 90612 9908 90670 10262
rect 91670 10554 91728 10908
rect 91670 10262 91682 10554
rect 91716 10262 91728 10554
rect 91670 9908 91728 10262
rect 92728 10554 92786 10908
rect 92728 10262 92740 10554
rect 92774 10262 92786 10554
rect 92728 9908 92786 10262
rect 93786 10554 93844 10908
rect 94964 11646 95022 12000
rect 94964 11354 94976 11646
rect 95010 11354 95022 11646
rect 94964 11000 95022 11354
rect 96022 11646 96080 12000
rect 96022 11354 96034 11646
rect 96068 11354 96080 11646
rect 96022 11000 96080 11354
rect 97080 11646 97138 12000
rect 97080 11354 97092 11646
rect 97126 11354 97138 11646
rect 97080 11000 97138 11354
rect 98138 11646 98196 12000
rect 98138 11354 98150 11646
rect 98184 11354 98196 11646
rect 98138 11000 98196 11354
rect 99196 11646 99254 12000
rect 99196 11354 99208 11646
rect 99242 11354 99254 11646
rect 99196 11000 99254 11354
rect 100254 11646 100312 12000
rect 100254 11354 100266 11646
rect 100300 11354 100312 11646
rect 100254 11000 100312 11354
rect 93786 10262 93798 10554
rect 93832 10262 93844 10554
rect 93786 9908 93844 10262
rect 94964 10552 95022 10906
rect 94964 10260 94976 10552
rect 95010 10260 95022 10552
rect 67396 9204 67408 9496
rect 67442 9204 67454 9496
rect 67396 8850 67454 9204
rect 68574 9494 68632 9848
rect 68574 9202 68586 9494
rect 68620 9202 68632 9494
rect 68574 8848 68632 9202
rect 69632 9494 69690 9848
rect 69632 9202 69644 9494
rect 69678 9202 69690 9494
rect 69632 8848 69690 9202
rect 70690 9494 70748 9848
rect 70690 9202 70702 9494
rect 70736 9202 70748 9494
rect 70690 8848 70748 9202
rect 71748 9494 71806 9848
rect 71748 9202 71760 9494
rect 71794 9202 71806 9494
rect 71748 8848 71806 9202
rect 72806 9494 72864 9848
rect 72806 9202 72818 9494
rect 72852 9202 72864 9494
rect 72806 8848 72864 9202
rect 73864 9494 73922 9848
rect 94964 9906 95022 10260
rect 96022 10552 96080 10906
rect 96022 10260 96034 10552
rect 96068 10260 96080 10552
rect 96022 9906 96080 10260
rect 97080 10552 97138 10906
rect 97080 10260 97092 10552
rect 97126 10260 97138 10552
rect 97080 9906 97138 10260
rect 98138 10552 98196 10906
rect 98138 10260 98150 10552
rect 98184 10260 98196 10552
rect 98138 9906 98196 10260
rect 99196 10552 99254 10906
rect 99196 10260 99208 10552
rect 99242 10260 99254 10552
rect 99196 9906 99254 10260
rect 100254 10552 100312 10906
rect 100254 10260 100266 10552
rect 100300 10260 100312 10552
rect 100254 9906 100312 10260
rect 73864 9202 73876 9494
rect 73910 9202 73922 9494
rect 73864 8848 73922 9202
rect 75262 9468 75320 9822
rect 75262 9176 75274 9468
rect 75308 9176 75320 9468
rect 75262 8822 75320 9176
rect 76320 9468 76378 9822
rect 76320 9176 76332 9468
rect 76366 9176 76378 9468
rect 76320 8822 76378 9176
rect 77378 9468 77436 9822
rect 77378 9176 77390 9468
rect 77424 9176 77436 9468
rect 77378 8822 77436 9176
rect 78436 9468 78494 9822
rect 78436 9176 78448 9468
rect 78482 9176 78494 9468
rect 78436 8822 78494 9176
rect 79494 9468 79552 9822
rect 79494 9176 79506 9468
rect 79540 9176 79552 9468
rect 79494 8822 79552 9176
rect 80552 9468 80610 9822
rect 80552 9176 80564 9468
rect 80598 9176 80610 9468
rect 80552 8822 80610 9176
rect 81730 9466 81788 9820
rect 81730 9174 81742 9466
rect 81776 9174 81788 9466
rect 81730 8820 81788 9174
rect 82788 9466 82846 9820
rect 82788 9174 82800 9466
rect 82834 9174 82846 9466
rect 82788 8820 82846 9174
rect 83846 9466 83904 9820
rect 83846 9174 83858 9466
rect 83892 9174 83904 9466
rect 83846 8820 83904 9174
rect 84904 9466 84962 9820
rect 84904 9174 84916 9466
rect 84950 9174 84962 9466
rect 84904 8820 84962 9174
rect 85962 9466 86020 9820
rect 85962 9174 85974 9466
rect 86008 9174 86020 9466
rect 85962 8820 86020 9174
rect 87020 9466 87078 9820
rect 87020 9174 87032 9466
rect 87066 9174 87078 9466
rect 87020 8820 87078 9174
rect 88496 9460 88554 9814
rect 88496 9168 88508 9460
rect 88542 9168 88554 9460
rect 88496 8814 88554 9168
rect 89554 9460 89612 9814
rect 89554 9168 89566 9460
rect 89600 9168 89612 9460
rect 89554 8814 89612 9168
rect 90612 9460 90670 9814
rect 90612 9168 90624 9460
rect 90658 9168 90670 9460
rect 90612 8814 90670 9168
rect 91670 9460 91728 9814
rect 91670 9168 91682 9460
rect 91716 9168 91728 9460
rect 91670 8814 91728 9168
rect 92728 9460 92786 9814
rect 92728 9168 92740 9460
rect 92774 9168 92786 9460
rect 92728 8814 92786 9168
rect 93786 9460 93844 9814
rect 93786 9168 93798 9460
rect 93832 9168 93844 9460
rect 93786 8814 93844 9168
rect 94964 9458 95022 9812
rect 94964 9166 94976 9458
rect 95010 9166 95022 9458
rect 62106 8014 62164 8368
rect 62106 7722 62118 8014
rect 62152 7722 62164 8014
rect 62106 7368 62164 7722
rect 63164 8014 63222 8368
rect 63164 7722 63176 8014
rect 63210 7722 63222 8014
rect 63164 7368 63222 7722
rect 64222 8014 64280 8368
rect 64222 7722 64234 8014
rect 64268 7722 64280 8014
rect 64222 7368 64280 7722
rect 65280 8014 65338 8368
rect 65280 7722 65292 8014
rect 65326 7722 65338 8014
rect 65280 7368 65338 7722
rect 66338 8014 66396 8368
rect 66338 7722 66350 8014
rect 66384 7722 66396 8014
rect 66338 7368 66396 7722
rect 67396 8014 67454 8368
rect 94964 8812 95022 9166
rect 96022 9458 96080 9812
rect 96022 9166 96034 9458
rect 96068 9166 96080 9458
rect 96022 8812 96080 9166
rect 97080 9458 97138 9812
rect 97080 9166 97092 9458
rect 97126 9166 97138 9458
rect 97080 8812 97138 9166
rect 98138 9458 98196 9812
rect 98138 9166 98150 9458
rect 98184 9166 98196 9458
rect 98138 8812 98196 9166
rect 99196 9458 99254 9812
rect 99196 9166 99208 9458
rect 99242 9166 99254 9458
rect 99196 8812 99254 9166
rect 100254 9458 100312 9812
rect 100254 9166 100266 9458
rect 100300 9166 100312 9458
rect 100254 8812 100312 9166
rect 67396 7722 67408 8014
rect 67442 7722 67454 8014
rect 67396 7368 67454 7722
rect 68578 8012 68636 8366
rect 68578 7720 68590 8012
rect 68624 7720 68636 8012
rect 68578 7366 68636 7720
rect 69636 8012 69694 8366
rect 69636 7720 69648 8012
rect 69682 7720 69694 8012
rect 69636 7366 69694 7720
rect 70694 8012 70752 8366
rect 70694 7720 70706 8012
rect 70740 7720 70752 8012
rect 70694 7366 70752 7720
rect 71752 8012 71810 8366
rect 71752 7720 71764 8012
rect 71798 7720 71810 8012
rect 71752 7366 71810 7720
rect 72810 8012 72868 8366
rect 72810 7720 72822 8012
rect 72856 7720 72868 8012
rect 72810 7366 72868 7720
rect 73868 8012 73926 8366
rect 73868 7720 73880 8012
rect 73914 7720 73926 8012
rect 73868 7366 73926 7720
rect 75262 7986 75320 8340
rect 75262 7694 75274 7986
rect 75308 7694 75320 7986
rect 75262 7340 75320 7694
rect 76320 7986 76378 8340
rect 76320 7694 76332 7986
rect 76366 7694 76378 7986
rect 76320 7340 76378 7694
rect 77378 7986 77436 8340
rect 77378 7694 77390 7986
rect 77424 7694 77436 7986
rect 77378 7340 77436 7694
rect 78436 7986 78494 8340
rect 78436 7694 78448 7986
rect 78482 7694 78494 7986
rect 78436 7340 78494 7694
rect 79494 7986 79552 8340
rect 79494 7694 79506 7986
rect 79540 7694 79552 7986
rect 79494 7340 79552 7694
rect 80552 7986 80610 8340
rect 80552 7694 80564 7986
rect 80598 7694 80610 7986
rect 80552 7340 80610 7694
rect 81734 7984 81792 8338
rect 81734 7692 81746 7984
rect 81780 7692 81792 7984
rect 81734 7338 81792 7692
rect 82792 7984 82850 8338
rect 82792 7692 82804 7984
rect 82838 7692 82850 7984
rect 82792 7338 82850 7692
rect 83850 7984 83908 8338
rect 83850 7692 83862 7984
rect 83896 7692 83908 7984
rect 83850 7338 83908 7692
rect 84908 7984 84966 8338
rect 84908 7692 84920 7984
rect 84954 7692 84966 7984
rect 84908 7338 84966 7692
rect 85966 7984 86024 8338
rect 85966 7692 85978 7984
rect 86012 7692 86024 7984
rect 85966 7338 86024 7692
rect 87024 7984 87082 8338
rect 87024 7692 87036 7984
rect 87070 7692 87082 7984
rect 87024 7338 87082 7692
rect 88496 7978 88554 8332
rect 88496 7686 88508 7978
rect 88542 7686 88554 7978
rect 62106 6920 62164 7274
rect 62106 6628 62118 6920
rect 62152 6628 62164 6920
rect 62106 6274 62164 6628
rect 63164 6920 63222 7274
rect 63164 6628 63176 6920
rect 63210 6628 63222 6920
rect 63164 6274 63222 6628
rect 64222 6920 64280 7274
rect 64222 6628 64234 6920
rect 64268 6628 64280 6920
rect 64222 6274 64280 6628
rect 65280 6920 65338 7274
rect 65280 6628 65292 6920
rect 65326 6628 65338 6920
rect 65280 6274 65338 6628
rect 66338 6920 66396 7274
rect 66338 6628 66350 6920
rect 66384 6628 66396 6920
rect 66338 6274 66396 6628
rect 67396 6920 67454 7274
rect 88496 7332 88554 7686
rect 89554 7978 89612 8332
rect 89554 7686 89566 7978
rect 89600 7686 89612 7978
rect 89554 7332 89612 7686
rect 90612 7978 90670 8332
rect 90612 7686 90624 7978
rect 90658 7686 90670 7978
rect 90612 7332 90670 7686
rect 91670 7978 91728 8332
rect 91670 7686 91682 7978
rect 91716 7686 91728 7978
rect 91670 7332 91728 7686
rect 92728 7978 92786 8332
rect 92728 7686 92740 7978
rect 92774 7686 92786 7978
rect 92728 7332 92786 7686
rect 93786 7978 93844 8332
rect 93786 7686 93798 7978
rect 93832 7686 93844 7978
rect 93786 7332 93844 7686
rect 94968 7976 95026 8330
rect 94968 7684 94980 7976
rect 95014 7684 95026 7976
rect 67396 6628 67408 6920
rect 67442 6628 67454 6920
rect 68578 6918 68636 7272
rect 67396 6274 67454 6628
rect 62106 5826 62164 6180
rect 62106 5534 62118 5826
rect 62152 5534 62164 5826
rect 62106 5180 62164 5534
rect 63164 5826 63222 6180
rect 63164 5534 63176 5826
rect 63210 5534 63222 5826
rect 63164 5180 63222 5534
rect 64222 5826 64280 6180
rect 64222 5534 64234 5826
rect 64268 5534 64280 5826
rect 64222 5180 64280 5534
rect 65280 5826 65338 6180
rect 65280 5534 65292 5826
rect 65326 5534 65338 5826
rect 65280 5180 65338 5534
rect 66338 5826 66396 6180
rect 66338 5534 66350 5826
rect 66384 5534 66396 5826
rect 66338 5180 66396 5534
rect 67396 5826 67454 6180
rect 67396 5534 67408 5826
rect 67442 5534 67454 5826
rect 67396 5180 67454 5534
rect 68578 6626 68590 6918
rect 68624 6626 68636 6918
rect 68578 6272 68636 6626
rect 69636 6918 69694 7272
rect 69636 6626 69648 6918
rect 69682 6626 69694 6918
rect 69636 6272 69694 6626
rect 70694 6918 70752 7272
rect 70694 6626 70706 6918
rect 70740 6626 70752 6918
rect 70694 6272 70752 6626
rect 71752 6918 71810 7272
rect 71752 6626 71764 6918
rect 71798 6626 71810 6918
rect 71752 6272 71810 6626
rect 72810 6918 72868 7272
rect 72810 6626 72822 6918
rect 72856 6626 72868 6918
rect 72810 6272 72868 6626
rect 73868 6918 73926 7272
rect 94968 7330 95026 7684
rect 96026 7976 96084 8330
rect 96026 7684 96038 7976
rect 96072 7684 96084 7976
rect 96026 7330 96084 7684
rect 97084 7976 97142 8330
rect 97084 7684 97096 7976
rect 97130 7684 97142 7976
rect 97084 7330 97142 7684
rect 98142 7976 98200 8330
rect 98142 7684 98154 7976
rect 98188 7684 98200 7976
rect 98142 7330 98200 7684
rect 99200 7976 99258 8330
rect 99200 7684 99212 7976
rect 99246 7684 99258 7976
rect 99200 7330 99258 7684
rect 100258 7976 100316 8330
rect 100258 7684 100270 7976
rect 100304 7684 100316 7976
rect 100258 7330 100316 7684
rect 73868 6626 73880 6918
rect 73914 6626 73926 6918
rect 73868 6272 73926 6626
rect 75262 6892 75320 7246
rect 62106 4732 62164 5086
rect 62106 4440 62118 4732
rect 62152 4440 62164 4732
rect 62106 4086 62164 4440
rect 63164 4732 63222 5086
rect 63164 4440 63176 4732
rect 63210 4440 63222 4732
rect 63164 4086 63222 4440
rect 64222 4732 64280 5086
rect 64222 4440 64234 4732
rect 64268 4440 64280 4732
rect 64222 4086 64280 4440
rect 65280 4732 65338 5086
rect 65280 4440 65292 4732
rect 65326 4440 65338 4732
rect 65280 4086 65338 4440
rect 66338 4732 66396 5086
rect 66338 4440 66350 4732
rect 66384 4440 66396 4732
rect 66338 4086 66396 4440
rect 67396 4732 67454 5086
rect 68578 5824 68636 6178
rect 68578 5532 68590 5824
rect 68624 5532 68636 5824
rect 68578 5178 68636 5532
rect 69636 5824 69694 6178
rect 69636 5532 69648 5824
rect 69682 5532 69694 5824
rect 69636 5178 69694 5532
rect 70694 5824 70752 6178
rect 70694 5532 70706 5824
rect 70740 5532 70752 5824
rect 70694 5178 70752 5532
rect 71752 5824 71810 6178
rect 71752 5532 71764 5824
rect 71798 5532 71810 5824
rect 71752 5178 71810 5532
rect 72810 5824 72868 6178
rect 72810 5532 72822 5824
rect 72856 5532 72868 5824
rect 72810 5178 72868 5532
rect 73868 5824 73926 6178
rect 73868 5532 73880 5824
rect 73914 5532 73926 5824
rect 73868 5178 73926 5532
rect 75262 6600 75274 6892
rect 75308 6600 75320 6892
rect 75262 6246 75320 6600
rect 76320 6892 76378 7246
rect 76320 6600 76332 6892
rect 76366 6600 76378 6892
rect 76320 6246 76378 6600
rect 77378 6892 77436 7246
rect 77378 6600 77390 6892
rect 77424 6600 77436 6892
rect 77378 6246 77436 6600
rect 78436 6892 78494 7246
rect 78436 6600 78448 6892
rect 78482 6600 78494 6892
rect 78436 6246 78494 6600
rect 79494 6892 79552 7246
rect 79494 6600 79506 6892
rect 79540 6600 79552 6892
rect 79494 6246 79552 6600
rect 80552 6892 80610 7246
rect 80552 6600 80564 6892
rect 80598 6600 80610 6892
rect 81734 6890 81792 7244
rect 80552 6246 80610 6600
rect 67396 4440 67408 4732
rect 67442 4440 67454 4732
rect 67396 4086 67454 4440
rect 68578 4730 68636 5084
rect 68578 4438 68590 4730
rect 68624 4438 68636 4730
rect 68578 4084 68636 4438
rect 69636 4730 69694 5084
rect 69636 4438 69648 4730
rect 69682 4438 69694 4730
rect 69636 4084 69694 4438
rect 70694 4730 70752 5084
rect 70694 4438 70706 4730
rect 70740 4438 70752 4730
rect 70694 4084 70752 4438
rect 71752 4730 71810 5084
rect 71752 4438 71764 4730
rect 71798 4438 71810 4730
rect 71752 4084 71810 4438
rect 72810 4730 72868 5084
rect 72810 4438 72822 4730
rect 72856 4438 72868 4730
rect 72810 4084 72868 4438
rect 73868 4730 73926 5084
rect 75262 5798 75320 6152
rect 75262 5506 75274 5798
rect 75308 5506 75320 5798
rect 75262 5152 75320 5506
rect 76320 5798 76378 6152
rect 76320 5506 76332 5798
rect 76366 5506 76378 5798
rect 76320 5152 76378 5506
rect 77378 5798 77436 6152
rect 77378 5506 77390 5798
rect 77424 5506 77436 5798
rect 77378 5152 77436 5506
rect 78436 5798 78494 6152
rect 78436 5506 78448 5798
rect 78482 5506 78494 5798
rect 78436 5152 78494 5506
rect 79494 5798 79552 6152
rect 79494 5506 79506 5798
rect 79540 5506 79552 5798
rect 79494 5152 79552 5506
rect 80552 5798 80610 6152
rect 80552 5506 80564 5798
rect 80598 5506 80610 5798
rect 80552 5152 80610 5506
rect 81734 6598 81746 6890
rect 81780 6598 81792 6890
rect 81734 6244 81792 6598
rect 82792 6890 82850 7244
rect 82792 6598 82804 6890
rect 82838 6598 82850 6890
rect 82792 6244 82850 6598
rect 83850 6890 83908 7244
rect 83850 6598 83862 6890
rect 83896 6598 83908 6890
rect 83850 6244 83908 6598
rect 84908 6890 84966 7244
rect 84908 6598 84920 6890
rect 84954 6598 84966 6890
rect 84908 6244 84966 6598
rect 85966 6890 86024 7244
rect 85966 6598 85978 6890
rect 86012 6598 86024 6890
rect 85966 6244 86024 6598
rect 87024 6890 87082 7244
rect 87024 6598 87036 6890
rect 87070 6598 87082 6890
rect 88496 6884 88554 7238
rect 87024 6244 87082 6598
rect 73868 4438 73880 4730
rect 73914 4438 73926 4730
rect 73868 4084 73926 4438
rect 75262 4704 75320 5058
rect 75262 4412 75274 4704
rect 75308 4412 75320 4704
rect 75262 4058 75320 4412
rect 76320 4704 76378 5058
rect 76320 4412 76332 4704
rect 76366 4412 76378 4704
rect 76320 4058 76378 4412
rect 77378 4704 77436 5058
rect 77378 4412 77390 4704
rect 77424 4412 77436 4704
rect 77378 4058 77436 4412
rect 78436 4704 78494 5058
rect 78436 4412 78448 4704
rect 78482 4412 78494 4704
rect 78436 4058 78494 4412
rect 79494 4704 79552 5058
rect 79494 4412 79506 4704
rect 79540 4412 79552 4704
rect 79494 4058 79552 4412
rect 80552 4704 80610 5058
rect 81734 5796 81792 6150
rect 81734 5504 81746 5796
rect 81780 5504 81792 5796
rect 81734 5150 81792 5504
rect 82792 5796 82850 6150
rect 82792 5504 82804 5796
rect 82838 5504 82850 5796
rect 82792 5150 82850 5504
rect 83850 5796 83908 6150
rect 83850 5504 83862 5796
rect 83896 5504 83908 5796
rect 83850 5150 83908 5504
rect 84908 5796 84966 6150
rect 84908 5504 84920 5796
rect 84954 5504 84966 5796
rect 84908 5150 84966 5504
rect 85966 5796 86024 6150
rect 85966 5504 85978 5796
rect 86012 5504 86024 5796
rect 85966 5150 86024 5504
rect 87024 5796 87082 6150
rect 87024 5504 87036 5796
rect 87070 5504 87082 5796
rect 87024 5150 87082 5504
rect 88496 6592 88508 6884
rect 88542 6592 88554 6884
rect 88496 6238 88554 6592
rect 89554 6884 89612 7238
rect 89554 6592 89566 6884
rect 89600 6592 89612 6884
rect 89554 6238 89612 6592
rect 90612 6884 90670 7238
rect 90612 6592 90624 6884
rect 90658 6592 90670 6884
rect 90612 6238 90670 6592
rect 91670 6884 91728 7238
rect 91670 6592 91682 6884
rect 91716 6592 91728 6884
rect 91670 6238 91728 6592
rect 92728 6884 92786 7238
rect 92728 6592 92740 6884
rect 92774 6592 92786 6884
rect 92728 6238 92786 6592
rect 93786 6884 93844 7238
rect 93786 6592 93798 6884
rect 93832 6592 93844 6884
rect 94968 6882 95026 7236
rect 93786 6238 93844 6592
rect 80552 4412 80564 4704
rect 80598 4412 80610 4704
rect 80552 4058 80610 4412
rect 81734 4702 81792 5056
rect 81734 4410 81746 4702
rect 81780 4410 81792 4702
rect 81734 4056 81792 4410
rect 82792 4702 82850 5056
rect 82792 4410 82804 4702
rect 82838 4410 82850 4702
rect 82792 4056 82850 4410
rect 83850 4702 83908 5056
rect 83850 4410 83862 4702
rect 83896 4410 83908 4702
rect 83850 4056 83908 4410
rect 84908 4702 84966 5056
rect 84908 4410 84920 4702
rect 84954 4410 84966 4702
rect 84908 4056 84966 4410
rect 85966 4702 86024 5056
rect 85966 4410 85978 4702
rect 86012 4410 86024 4702
rect 85966 4056 86024 4410
rect 87024 4702 87082 5056
rect 88496 5790 88554 6144
rect 88496 5498 88508 5790
rect 88542 5498 88554 5790
rect 88496 5144 88554 5498
rect 89554 5790 89612 6144
rect 89554 5498 89566 5790
rect 89600 5498 89612 5790
rect 89554 5144 89612 5498
rect 90612 5790 90670 6144
rect 90612 5498 90624 5790
rect 90658 5498 90670 5790
rect 90612 5144 90670 5498
rect 91670 5790 91728 6144
rect 91670 5498 91682 5790
rect 91716 5498 91728 5790
rect 91670 5144 91728 5498
rect 92728 5790 92786 6144
rect 92728 5498 92740 5790
rect 92774 5498 92786 5790
rect 92728 5144 92786 5498
rect 93786 5790 93844 6144
rect 93786 5498 93798 5790
rect 93832 5498 93844 5790
rect 93786 5144 93844 5498
rect 94968 6590 94980 6882
rect 95014 6590 95026 6882
rect 94968 6236 95026 6590
rect 96026 6882 96084 7236
rect 96026 6590 96038 6882
rect 96072 6590 96084 6882
rect 96026 6236 96084 6590
rect 97084 6882 97142 7236
rect 97084 6590 97096 6882
rect 97130 6590 97142 6882
rect 97084 6236 97142 6590
rect 98142 6882 98200 7236
rect 98142 6590 98154 6882
rect 98188 6590 98200 6882
rect 98142 6236 98200 6590
rect 99200 6882 99258 7236
rect 99200 6590 99212 6882
rect 99246 6590 99258 6882
rect 99200 6236 99258 6590
rect 100258 6882 100316 7236
rect 100258 6590 100270 6882
rect 100304 6590 100316 6882
rect 100258 6236 100316 6590
rect 87024 4410 87036 4702
rect 87070 4410 87082 4702
rect 87024 4056 87082 4410
rect 88496 4696 88554 5050
rect 88496 4404 88508 4696
rect 88542 4404 88554 4696
rect 62106 3638 62164 3992
rect 62106 3346 62118 3638
rect 62152 3346 62164 3638
rect 62106 2992 62164 3346
rect 63164 3638 63222 3992
rect 63164 3346 63176 3638
rect 63210 3346 63222 3638
rect 63164 2992 63222 3346
rect 64222 3638 64280 3992
rect 64222 3346 64234 3638
rect 64268 3346 64280 3638
rect 64222 2992 64280 3346
rect 65280 3638 65338 3992
rect 65280 3346 65292 3638
rect 65326 3346 65338 3638
rect 65280 2992 65338 3346
rect 66338 3638 66396 3992
rect 66338 3346 66350 3638
rect 66384 3346 66396 3638
rect 66338 2992 66396 3346
rect 67396 3638 67454 3992
rect 88496 4050 88554 4404
rect 89554 4696 89612 5050
rect 89554 4404 89566 4696
rect 89600 4404 89612 4696
rect 89554 4050 89612 4404
rect 90612 4696 90670 5050
rect 90612 4404 90624 4696
rect 90658 4404 90670 4696
rect 90612 4050 90670 4404
rect 91670 4696 91728 5050
rect 91670 4404 91682 4696
rect 91716 4404 91728 4696
rect 91670 4050 91728 4404
rect 92728 4696 92786 5050
rect 92728 4404 92740 4696
rect 92774 4404 92786 4696
rect 92728 4050 92786 4404
rect 93786 4696 93844 5050
rect 94968 5788 95026 6142
rect 94968 5496 94980 5788
rect 95014 5496 95026 5788
rect 94968 5142 95026 5496
rect 96026 5788 96084 6142
rect 96026 5496 96038 5788
rect 96072 5496 96084 5788
rect 96026 5142 96084 5496
rect 97084 5788 97142 6142
rect 97084 5496 97096 5788
rect 97130 5496 97142 5788
rect 97084 5142 97142 5496
rect 98142 5788 98200 6142
rect 98142 5496 98154 5788
rect 98188 5496 98200 5788
rect 98142 5142 98200 5496
rect 99200 5788 99258 6142
rect 99200 5496 99212 5788
rect 99246 5496 99258 5788
rect 99200 5142 99258 5496
rect 100258 5788 100316 6142
rect 100258 5496 100270 5788
rect 100304 5496 100316 5788
rect 100258 5142 100316 5496
rect 93786 4404 93798 4696
rect 93832 4404 93844 4696
rect 93786 4050 93844 4404
rect 94968 4694 95026 5048
rect 94968 4402 94980 4694
rect 95014 4402 95026 4694
rect 67396 3346 67408 3638
rect 67442 3346 67454 3638
rect 67396 2992 67454 3346
rect 68578 3636 68636 3990
rect 68578 3344 68590 3636
rect 68624 3344 68636 3636
rect 68578 2990 68636 3344
rect 69636 3636 69694 3990
rect 69636 3344 69648 3636
rect 69682 3344 69694 3636
rect 69636 2990 69694 3344
rect 70694 3636 70752 3990
rect 70694 3344 70706 3636
rect 70740 3344 70752 3636
rect 70694 2990 70752 3344
rect 71752 3636 71810 3990
rect 71752 3344 71764 3636
rect 71798 3344 71810 3636
rect 71752 2990 71810 3344
rect 72810 3636 72868 3990
rect 72810 3344 72822 3636
rect 72856 3344 72868 3636
rect 72810 2990 72868 3344
rect 73868 3636 73926 3990
rect 94968 4048 95026 4402
rect 96026 4694 96084 5048
rect 96026 4402 96038 4694
rect 96072 4402 96084 4694
rect 96026 4048 96084 4402
rect 97084 4694 97142 5048
rect 97084 4402 97096 4694
rect 97130 4402 97142 4694
rect 97084 4048 97142 4402
rect 98142 4694 98200 5048
rect 98142 4402 98154 4694
rect 98188 4402 98200 4694
rect 98142 4048 98200 4402
rect 99200 4694 99258 5048
rect 99200 4402 99212 4694
rect 99246 4402 99258 4694
rect 99200 4048 99258 4402
rect 100258 4694 100316 5048
rect 100258 4402 100270 4694
rect 100304 4402 100316 4694
rect 100258 4048 100316 4402
rect 73868 3344 73880 3636
rect 73914 3344 73926 3636
rect 73868 2990 73926 3344
rect 75262 3610 75320 3964
rect 75262 3318 75274 3610
rect 75308 3318 75320 3610
rect 75262 2964 75320 3318
rect 76320 3610 76378 3964
rect 76320 3318 76332 3610
rect 76366 3318 76378 3610
rect 76320 2964 76378 3318
rect 77378 3610 77436 3964
rect 77378 3318 77390 3610
rect 77424 3318 77436 3610
rect 77378 2964 77436 3318
rect 78436 3610 78494 3964
rect 78436 3318 78448 3610
rect 78482 3318 78494 3610
rect 78436 2964 78494 3318
rect 79494 3610 79552 3964
rect 79494 3318 79506 3610
rect 79540 3318 79552 3610
rect 79494 2964 79552 3318
rect 80552 3610 80610 3964
rect 80552 3318 80564 3610
rect 80598 3318 80610 3610
rect 80552 2964 80610 3318
rect 81734 3608 81792 3962
rect 81734 3316 81746 3608
rect 81780 3316 81792 3608
rect 81734 2962 81792 3316
rect 82792 3608 82850 3962
rect 82792 3316 82804 3608
rect 82838 3316 82850 3608
rect 82792 2962 82850 3316
rect 83850 3608 83908 3962
rect 83850 3316 83862 3608
rect 83896 3316 83908 3608
rect 83850 2962 83908 3316
rect 84908 3608 84966 3962
rect 84908 3316 84920 3608
rect 84954 3316 84966 3608
rect 84908 2962 84966 3316
rect 85966 3608 86024 3962
rect 85966 3316 85978 3608
rect 86012 3316 86024 3608
rect 85966 2962 86024 3316
rect 87024 3608 87082 3962
rect 87024 3316 87036 3608
rect 87070 3316 87082 3608
rect 87024 2962 87082 3316
rect 88496 3602 88554 3956
rect 88496 3310 88508 3602
rect 88542 3310 88554 3602
rect 88496 2956 88554 3310
rect 89554 3602 89612 3956
rect 89554 3310 89566 3602
rect 89600 3310 89612 3602
rect 89554 2956 89612 3310
rect 90612 3602 90670 3956
rect 90612 3310 90624 3602
rect 90658 3310 90670 3602
rect 90612 2956 90670 3310
rect 91670 3602 91728 3956
rect 91670 3310 91682 3602
rect 91716 3310 91728 3602
rect 91670 2956 91728 3310
rect 92728 3602 92786 3956
rect 92728 3310 92740 3602
rect 92774 3310 92786 3602
rect 92728 2956 92786 3310
rect 93786 3602 93844 3956
rect 93786 3310 93798 3602
rect 93832 3310 93844 3602
rect 93786 2956 93844 3310
rect 94968 3600 95026 3954
rect 94968 3308 94980 3600
rect 95014 3308 95026 3600
rect 94968 2954 95026 3308
rect 96026 3600 96084 3954
rect 96026 3308 96038 3600
rect 96072 3308 96084 3600
rect 96026 2954 96084 3308
rect 97084 3600 97142 3954
rect 97084 3308 97096 3600
rect 97130 3308 97142 3600
rect 97084 2954 97142 3308
rect 98142 3600 98200 3954
rect 98142 3308 98154 3600
rect 98188 3308 98200 3600
rect 98142 2954 98200 3308
rect 99200 3600 99258 3954
rect 99200 3308 99212 3600
rect 99246 3308 99258 3600
rect 99200 2954 99258 3308
rect 100258 3600 100316 3954
rect 100258 3308 100270 3600
rect 100304 3308 100316 3600
rect 100258 2954 100316 3308
<< mvpdiff >>
rect 71326 74040 71384 74254
rect 42196 73228 42796 73240
rect 42196 73194 42410 73228
rect 42582 73194 42796 73228
rect 42196 73182 42796 73194
rect 42890 73228 43490 73240
rect 42890 73194 43104 73228
rect 43276 73194 43490 73228
rect 42890 73182 43490 73194
rect 43584 73228 44184 73240
rect 43584 73194 43798 73228
rect 43970 73194 44184 73228
rect 43584 73182 44184 73194
rect 44278 73228 44878 73240
rect 44278 73194 44492 73228
rect 44664 73194 44878 73228
rect 44278 73182 44878 73194
rect 44972 73228 45572 73240
rect 44972 73194 45186 73228
rect 45358 73194 45572 73228
rect 44972 73182 45572 73194
rect 46204 73226 46804 73238
rect 46204 73192 46418 73226
rect 46590 73192 46804 73226
rect 46204 73180 46804 73192
rect 46898 73226 47498 73238
rect 46898 73192 47112 73226
rect 47284 73192 47498 73226
rect 46898 73180 47498 73192
rect 47592 73226 48192 73238
rect 47592 73192 47806 73226
rect 47978 73192 48192 73226
rect 47592 73180 48192 73192
rect 48286 73226 48886 73238
rect 48286 73192 48500 73226
rect 48672 73192 48886 73226
rect 48286 73180 48886 73192
rect 48980 73226 49580 73238
rect 48980 73192 49194 73226
rect 49366 73192 49580 73226
rect 48980 73180 49580 73192
rect 50216 73226 50816 73238
rect 50216 73192 50430 73226
rect 50602 73192 50816 73226
rect 50216 73180 50816 73192
rect 50910 73226 51510 73238
rect 50910 73192 51124 73226
rect 51296 73192 51510 73226
rect 50910 73180 51510 73192
rect 51604 73226 52204 73238
rect 51604 73192 51818 73226
rect 51990 73192 52204 73226
rect 51604 73180 52204 73192
rect 52298 73226 52898 73238
rect 52298 73192 52512 73226
rect 52684 73192 52898 73226
rect 52298 73180 52898 73192
rect 52992 73226 53592 73238
rect 52992 73192 53206 73226
rect 53378 73192 53592 73226
rect 52992 73180 53592 73192
rect 54226 73226 54826 73238
rect 54226 73192 54440 73226
rect 54612 73192 54826 73226
rect 54226 73180 54826 73192
rect 54920 73226 55520 73238
rect 54920 73192 55134 73226
rect 55306 73192 55520 73226
rect 54920 73180 55520 73192
rect 55614 73226 56214 73238
rect 55614 73192 55828 73226
rect 56000 73192 56214 73226
rect 55614 73180 56214 73192
rect 56308 73226 56908 73238
rect 56308 73192 56522 73226
rect 56694 73192 56908 73226
rect 56308 73180 56908 73192
rect 57002 73226 57602 73238
rect 57002 73192 57216 73226
rect 57388 73192 57602 73226
rect 57002 73180 57602 73192
rect 42196 72570 42796 72582
rect 42196 72536 42410 72570
rect 42582 72536 42796 72570
rect 42196 72524 42796 72536
rect 42890 72570 43490 72582
rect 42890 72536 43104 72570
rect 43276 72536 43490 72570
rect 42890 72524 43490 72536
rect 43584 72570 44184 72582
rect 43584 72536 43798 72570
rect 43970 72536 44184 72570
rect 43584 72524 44184 72536
rect 44278 72570 44878 72582
rect 44278 72536 44492 72570
rect 44664 72536 44878 72570
rect 44278 72524 44878 72536
rect 44972 72570 45572 72582
rect 44972 72536 45186 72570
rect 45358 72536 45572 72570
rect 44972 72524 45572 72536
rect 71326 73868 71338 74040
rect 71372 73868 71384 74040
rect 71326 73654 71384 73868
rect 71984 74040 72042 74254
rect 71984 73868 71996 74040
rect 72030 73868 72042 74040
rect 71984 73654 72042 73868
rect 72642 74040 72700 74254
rect 72642 73868 72654 74040
rect 72688 73868 72700 74040
rect 72642 73654 72700 73868
rect 73300 74040 73358 74254
rect 73300 73868 73312 74040
rect 73346 73868 73358 74040
rect 73300 73654 73358 73868
rect 73958 74040 74016 74254
rect 73958 73868 73970 74040
rect 74004 73868 74016 74040
rect 73958 73654 74016 73868
rect 75190 74020 75248 74234
rect 75190 73848 75202 74020
rect 75236 73848 75248 74020
rect 75190 73634 75248 73848
rect 75848 74020 75906 74234
rect 75848 73848 75860 74020
rect 75894 73848 75906 74020
rect 75848 73634 75906 73848
rect 76506 74020 76564 74234
rect 76506 73848 76518 74020
rect 76552 73848 76564 74020
rect 76506 73634 76564 73848
rect 77164 74020 77222 74234
rect 77164 73848 77176 74020
rect 77210 73848 77222 74020
rect 77164 73634 77222 73848
rect 77822 74020 77880 74234
rect 77822 73848 77834 74020
rect 77868 73848 77880 74020
rect 77822 73634 77880 73848
rect 79040 74034 79098 74248
rect 79040 73862 79052 74034
rect 79086 73862 79098 74034
rect 79040 73648 79098 73862
rect 79698 74034 79756 74248
rect 79698 73862 79710 74034
rect 79744 73862 79756 74034
rect 79698 73648 79756 73862
rect 80356 74034 80414 74248
rect 80356 73862 80368 74034
rect 80402 73862 80414 74034
rect 80356 73648 80414 73862
rect 81014 74034 81072 74248
rect 81014 73862 81026 74034
rect 81060 73862 81072 74034
rect 81014 73648 81072 73862
rect 81672 74034 81730 74248
rect 81672 73862 81684 74034
rect 81718 73862 81730 74034
rect 81672 73648 81730 73862
rect 46204 72568 46804 72580
rect 46204 72534 46418 72568
rect 46590 72534 46804 72568
rect 46204 72522 46804 72534
rect 46898 72568 47498 72580
rect 46898 72534 47112 72568
rect 47284 72534 47498 72568
rect 46898 72522 47498 72534
rect 47592 72568 48192 72580
rect 47592 72534 47806 72568
rect 47978 72534 48192 72568
rect 47592 72522 48192 72534
rect 48286 72568 48886 72580
rect 48286 72534 48500 72568
rect 48672 72534 48886 72568
rect 48286 72522 48886 72534
rect 48980 72568 49580 72580
rect 48980 72534 49194 72568
rect 49366 72534 49580 72568
rect 48980 72522 49580 72534
rect 50216 72568 50816 72580
rect 50216 72534 50430 72568
rect 50602 72534 50816 72568
rect 50216 72522 50816 72534
rect 50910 72568 51510 72580
rect 50910 72534 51124 72568
rect 51296 72534 51510 72568
rect 50910 72522 51510 72534
rect 51604 72568 52204 72580
rect 51604 72534 51818 72568
rect 51990 72534 52204 72568
rect 51604 72522 52204 72534
rect 52298 72568 52898 72580
rect 52298 72534 52512 72568
rect 52684 72534 52898 72568
rect 52298 72522 52898 72534
rect 52992 72568 53592 72580
rect 52992 72534 53206 72568
rect 53378 72534 53592 72568
rect 52992 72522 53592 72534
rect 54226 72568 54826 72580
rect 54226 72534 54440 72568
rect 54612 72534 54826 72568
rect 54226 72522 54826 72534
rect 54920 72568 55520 72580
rect 54920 72534 55134 72568
rect 55306 72534 55520 72568
rect 54920 72522 55520 72534
rect 55614 72568 56214 72580
rect 55614 72534 55828 72568
rect 56000 72534 56214 72568
rect 55614 72522 56214 72534
rect 56308 72568 56908 72580
rect 56308 72534 56522 72568
rect 56694 72534 56908 72568
rect 56308 72522 56908 72534
rect 57002 72568 57602 72580
rect 57002 72534 57216 72568
rect 57388 72534 57602 72568
rect 57002 72522 57602 72534
rect 42196 71912 42796 71924
rect 42196 71878 42410 71912
rect 42582 71878 42796 71912
rect 42196 71866 42796 71878
rect 42890 71912 43490 71924
rect 42890 71878 43104 71912
rect 43276 71878 43490 71912
rect 42890 71866 43490 71878
rect 43584 71912 44184 71924
rect 43584 71878 43798 71912
rect 43970 71878 44184 71912
rect 43584 71866 44184 71878
rect 44278 71912 44878 71924
rect 44278 71878 44492 71912
rect 44664 71878 44878 71912
rect 44278 71866 44878 71878
rect 44972 71912 45572 71924
rect 44972 71878 45186 71912
rect 45358 71878 45572 71912
rect 44972 71866 45572 71878
rect 46204 71910 46804 71922
rect 46204 71876 46418 71910
rect 46590 71876 46804 71910
rect 46204 71864 46804 71876
rect 46898 71910 47498 71922
rect 46898 71876 47112 71910
rect 47284 71876 47498 71910
rect 46898 71864 47498 71876
rect 47592 71910 48192 71922
rect 47592 71876 47806 71910
rect 47978 71876 48192 71910
rect 47592 71864 48192 71876
rect 48286 71910 48886 71922
rect 48286 71876 48500 71910
rect 48672 71876 48886 71910
rect 48286 71864 48886 71876
rect 48980 71910 49580 71922
rect 48980 71876 49194 71910
rect 49366 71876 49580 71910
rect 48980 71864 49580 71876
rect 50216 71910 50816 71922
rect 50216 71876 50430 71910
rect 50602 71876 50816 71910
rect 50216 71864 50816 71876
rect 50910 71910 51510 71922
rect 50910 71876 51124 71910
rect 51296 71876 51510 71910
rect 50910 71864 51510 71876
rect 51604 71910 52204 71922
rect 51604 71876 51818 71910
rect 51990 71876 52204 71910
rect 51604 71864 52204 71876
rect 52298 71910 52898 71922
rect 52298 71876 52512 71910
rect 52684 71876 52898 71910
rect 52298 71864 52898 71876
rect 52992 71910 53592 71922
rect 52992 71876 53206 71910
rect 53378 71876 53592 71910
rect 52992 71864 53592 71876
rect 54226 71910 54826 71922
rect 54226 71876 54440 71910
rect 54612 71876 54826 71910
rect 54226 71864 54826 71876
rect 54920 71910 55520 71922
rect 54920 71876 55134 71910
rect 55306 71876 55520 71910
rect 54920 71864 55520 71876
rect 55614 71910 56214 71922
rect 55614 71876 55828 71910
rect 56000 71876 56214 71910
rect 55614 71864 56214 71876
rect 56308 71910 56908 71922
rect 56308 71876 56522 71910
rect 56694 71876 56908 71910
rect 56308 71864 56908 71876
rect 57002 71910 57602 71922
rect 57002 71876 57216 71910
rect 57388 71876 57602 71910
rect 57002 71864 57602 71876
rect 42196 71254 42796 71266
rect 42196 71220 42410 71254
rect 42582 71220 42796 71254
rect 42196 71208 42796 71220
rect 42890 71254 43490 71266
rect 42890 71220 43104 71254
rect 43276 71220 43490 71254
rect 42890 71208 43490 71220
rect 43584 71254 44184 71266
rect 43584 71220 43798 71254
rect 43970 71220 44184 71254
rect 43584 71208 44184 71220
rect 44278 71254 44878 71266
rect 44278 71220 44492 71254
rect 44664 71220 44878 71254
rect 44278 71208 44878 71220
rect 44972 71254 45572 71266
rect 44972 71220 45186 71254
rect 45358 71220 45572 71254
rect 44972 71208 45572 71220
rect 46204 71252 46804 71264
rect 46204 71218 46418 71252
rect 46590 71218 46804 71252
rect 46204 71206 46804 71218
rect 46898 71252 47498 71264
rect 46898 71218 47112 71252
rect 47284 71218 47498 71252
rect 46898 71206 47498 71218
rect 47592 71252 48192 71264
rect 47592 71218 47806 71252
rect 47978 71218 48192 71252
rect 47592 71206 48192 71218
rect 48286 71252 48886 71264
rect 48286 71218 48500 71252
rect 48672 71218 48886 71252
rect 48286 71206 48886 71218
rect 48980 71252 49580 71264
rect 48980 71218 49194 71252
rect 49366 71218 49580 71252
rect 48980 71206 49580 71218
rect 50216 71252 50816 71264
rect 50216 71218 50430 71252
rect 50602 71218 50816 71252
rect 50216 71206 50816 71218
rect 50910 71252 51510 71264
rect 50910 71218 51124 71252
rect 51296 71218 51510 71252
rect 50910 71206 51510 71218
rect 51604 71252 52204 71264
rect 51604 71218 51818 71252
rect 51990 71218 52204 71252
rect 51604 71206 52204 71218
rect 52298 71252 52898 71264
rect 52298 71218 52512 71252
rect 52684 71218 52898 71252
rect 52298 71206 52898 71218
rect 52992 71252 53592 71264
rect 52992 71218 53206 71252
rect 53378 71218 53592 71252
rect 52992 71206 53592 71218
rect 54226 71252 54826 71264
rect 54226 71218 54440 71252
rect 54612 71218 54826 71252
rect 54226 71206 54826 71218
rect 54920 71252 55520 71264
rect 54920 71218 55134 71252
rect 55306 71218 55520 71252
rect 54920 71206 55520 71218
rect 55614 71252 56214 71264
rect 55614 71218 55828 71252
rect 56000 71218 56214 71252
rect 55614 71206 56214 71218
rect 56308 71252 56908 71264
rect 56308 71218 56522 71252
rect 56694 71218 56908 71252
rect 56308 71206 56908 71218
rect 57002 71252 57602 71264
rect 57002 71218 57216 71252
rect 57388 71218 57602 71252
rect 57002 71206 57602 71218
rect 42196 70596 42796 70608
rect 42196 70562 42410 70596
rect 42582 70562 42796 70596
rect 42196 70550 42796 70562
rect 42890 70596 43490 70608
rect 42890 70562 43104 70596
rect 43276 70562 43490 70596
rect 42890 70550 43490 70562
rect 43584 70596 44184 70608
rect 43584 70562 43798 70596
rect 43970 70562 44184 70596
rect 43584 70550 44184 70562
rect 44278 70596 44878 70608
rect 44278 70562 44492 70596
rect 44664 70562 44878 70596
rect 44278 70550 44878 70562
rect 44972 70596 45572 70608
rect 44972 70562 45186 70596
rect 45358 70562 45572 70596
rect 44972 70550 45572 70562
rect 46204 70594 46804 70606
rect 46204 70560 46418 70594
rect 46590 70560 46804 70594
rect 46204 70548 46804 70560
rect 46898 70594 47498 70606
rect 46898 70560 47112 70594
rect 47284 70560 47498 70594
rect 46898 70548 47498 70560
rect 47592 70594 48192 70606
rect 47592 70560 47806 70594
rect 47978 70560 48192 70594
rect 47592 70548 48192 70560
rect 48286 70594 48886 70606
rect 48286 70560 48500 70594
rect 48672 70560 48886 70594
rect 48286 70548 48886 70560
rect 48980 70594 49580 70606
rect 48980 70560 49194 70594
rect 49366 70560 49580 70594
rect 48980 70548 49580 70560
rect 50216 70594 50816 70606
rect 50216 70560 50430 70594
rect 50602 70560 50816 70594
rect 50216 70548 50816 70560
rect 50910 70594 51510 70606
rect 50910 70560 51124 70594
rect 51296 70560 51510 70594
rect 50910 70548 51510 70560
rect 51604 70594 52204 70606
rect 51604 70560 51818 70594
rect 51990 70560 52204 70594
rect 51604 70548 52204 70560
rect 52298 70594 52898 70606
rect 52298 70560 52512 70594
rect 52684 70560 52898 70594
rect 52298 70548 52898 70560
rect 52992 70594 53592 70606
rect 52992 70560 53206 70594
rect 53378 70560 53592 70594
rect 52992 70548 53592 70560
rect 54226 70594 54826 70606
rect 54226 70560 54440 70594
rect 54612 70560 54826 70594
rect 54226 70548 54826 70560
rect 54920 70594 55520 70606
rect 54920 70560 55134 70594
rect 55306 70560 55520 70594
rect 54920 70548 55520 70560
rect 55614 70594 56214 70606
rect 55614 70560 55828 70594
rect 56000 70560 56214 70594
rect 55614 70548 56214 70560
rect 56308 70594 56908 70606
rect 56308 70560 56522 70594
rect 56694 70560 56908 70594
rect 56308 70548 56908 70560
rect 57002 70594 57602 70606
rect 57002 70560 57216 70594
rect 57388 70560 57602 70594
rect 57002 70548 57602 70560
rect 42196 69938 42796 69950
rect 42196 69904 42410 69938
rect 42582 69904 42796 69938
rect 42196 69892 42796 69904
rect 42890 69938 43490 69950
rect 42890 69904 43104 69938
rect 43276 69904 43490 69938
rect 42890 69892 43490 69904
rect 43584 69938 44184 69950
rect 43584 69904 43798 69938
rect 43970 69904 44184 69938
rect 43584 69892 44184 69904
rect 44278 69938 44878 69950
rect 44278 69904 44492 69938
rect 44664 69904 44878 69938
rect 44278 69892 44878 69904
rect 44972 69938 45572 69950
rect 44972 69904 45186 69938
rect 45358 69904 45572 69938
rect 44972 69892 45572 69904
rect 46204 69936 46804 69948
rect 46204 69902 46418 69936
rect 46590 69902 46804 69936
rect 46204 69890 46804 69902
rect 46898 69936 47498 69948
rect 46898 69902 47112 69936
rect 47284 69902 47498 69936
rect 46898 69890 47498 69902
rect 47592 69936 48192 69948
rect 47592 69902 47806 69936
rect 47978 69902 48192 69936
rect 47592 69890 48192 69902
rect 48286 69936 48886 69948
rect 48286 69902 48500 69936
rect 48672 69902 48886 69936
rect 48286 69890 48886 69902
rect 48980 69936 49580 69948
rect 48980 69902 49194 69936
rect 49366 69902 49580 69936
rect 48980 69890 49580 69902
rect 50216 69936 50816 69948
rect 50216 69902 50430 69936
rect 50602 69902 50816 69936
rect 50216 69890 50816 69902
rect 50910 69936 51510 69948
rect 50910 69902 51124 69936
rect 51296 69902 51510 69936
rect 50910 69890 51510 69902
rect 51604 69936 52204 69948
rect 51604 69902 51818 69936
rect 51990 69902 52204 69936
rect 51604 69890 52204 69902
rect 52298 69936 52898 69948
rect 52298 69902 52512 69936
rect 52684 69902 52898 69936
rect 52298 69890 52898 69902
rect 52992 69936 53592 69948
rect 52992 69902 53206 69936
rect 53378 69902 53592 69936
rect 52992 69890 53592 69902
rect 54226 69936 54826 69948
rect 54226 69902 54440 69936
rect 54612 69902 54826 69936
rect 54226 69890 54826 69902
rect 54920 69936 55520 69948
rect 54920 69902 55134 69936
rect 55306 69902 55520 69936
rect 54920 69890 55520 69902
rect 55614 69936 56214 69948
rect 55614 69902 55828 69936
rect 56000 69902 56214 69936
rect 55614 69890 56214 69902
rect 56308 69936 56908 69948
rect 56308 69902 56522 69936
rect 56694 69902 56908 69936
rect 56308 69890 56908 69902
rect 57002 69936 57602 69948
rect 57002 69902 57216 69936
rect 57388 69902 57602 69936
rect 57002 69890 57602 69902
rect 42188 69030 42788 69042
rect 42188 68996 42402 69030
rect 42574 68996 42788 69030
rect 42188 68984 42788 68996
rect 42882 69030 43482 69042
rect 42882 68996 43096 69030
rect 43268 68996 43482 69030
rect 42882 68984 43482 68996
rect 43576 69030 44176 69042
rect 43576 68996 43790 69030
rect 43962 68996 44176 69030
rect 43576 68984 44176 68996
rect 44270 69030 44870 69042
rect 44270 68996 44484 69030
rect 44656 68996 44870 69030
rect 44270 68984 44870 68996
rect 44964 69030 45564 69042
rect 44964 68996 45178 69030
rect 45350 68996 45564 69030
rect 44964 68984 45564 68996
rect 46182 69030 46782 69042
rect 46182 68996 46396 69030
rect 46568 68996 46782 69030
rect 46182 68984 46782 68996
rect 46876 69030 47476 69042
rect 46876 68996 47090 69030
rect 47262 68996 47476 69030
rect 46876 68984 47476 68996
rect 47570 69030 48170 69042
rect 47570 68996 47784 69030
rect 47956 68996 48170 69030
rect 47570 68984 48170 68996
rect 48264 69030 48864 69042
rect 48264 68996 48478 69030
rect 48650 68996 48864 69030
rect 48264 68984 48864 68996
rect 48958 69030 49558 69042
rect 48958 68996 49172 69030
rect 49344 68996 49558 69030
rect 48958 68984 49558 68996
rect 50204 69030 50804 69042
rect 50204 68996 50418 69030
rect 50590 68996 50804 69030
rect 50204 68984 50804 68996
rect 50898 69030 51498 69042
rect 50898 68996 51112 69030
rect 51284 68996 51498 69030
rect 50898 68984 51498 68996
rect 51592 69030 52192 69042
rect 51592 68996 51806 69030
rect 51978 68996 52192 69030
rect 51592 68984 52192 68996
rect 52286 69030 52886 69042
rect 52286 68996 52500 69030
rect 52672 68996 52886 69030
rect 52286 68984 52886 68996
rect 52980 69030 53580 69042
rect 52980 68996 53194 69030
rect 53366 68996 53580 69030
rect 52980 68984 53580 68996
rect 54226 69030 54826 69042
rect 54226 68996 54440 69030
rect 54612 68996 54826 69030
rect 54226 68984 54826 68996
rect 54920 69030 55520 69042
rect 54920 68996 55134 69030
rect 55306 68996 55520 69030
rect 54920 68984 55520 68996
rect 55614 69030 56214 69042
rect 55614 68996 55828 69030
rect 56000 68996 56214 69030
rect 55614 68984 56214 68996
rect 56308 69030 56908 69042
rect 56308 68996 56522 69030
rect 56694 68996 56908 69030
rect 56308 68984 56908 68996
rect 57002 69030 57602 69042
rect 57002 68996 57216 69030
rect 57388 68996 57602 69030
rect 57002 68984 57602 68996
rect 71298 73126 71356 73340
rect 71298 72954 71310 73126
rect 71344 72954 71356 73126
rect 71298 72740 71356 72954
rect 71956 73126 72014 73340
rect 71956 72954 71968 73126
rect 72002 72954 72014 73126
rect 71956 72740 72014 72954
rect 72614 73126 72672 73340
rect 72614 72954 72626 73126
rect 72660 72954 72672 73126
rect 72614 72740 72672 72954
rect 73272 73126 73330 73340
rect 73272 72954 73284 73126
rect 73318 72954 73330 73126
rect 73272 72740 73330 72954
rect 73930 73126 73988 73340
rect 73930 72954 73942 73126
rect 73976 72954 73988 73126
rect 75162 73106 75220 73320
rect 73930 72740 73988 72954
rect 71298 72432 71356 72646
rect 71298 72260 71310 72432
rect 71344 72260 71356 72432
rect 71298 72046 71356 72260
rect 71956 72432 72014 72646
rect 71956 72260 71968 72432
rect 72002 72260 72014 72432
rect 71956 72046 72014 72260
rect 72614 72432 72672 72646
rect 72614 72260 72626 72432
rect 72660 72260 72672 72432
rect 72614 72046 72672 72260
rect 73272 72432 73330 72646
rect 73272 72260 73284 72432
rect 73318 72260 73330 72432
rect 73272 72046 73330 72260
rect 73930 72432 73988 72646
rect 73930 72260 73942 72432
rect 73976 72260 73988 72432
rect 73930 72046 73988 72260
rect 71298 71738 71356 71952
rect 71298 71566 71310 71738
rect 71344 71566 71356 71738
rect 71298 71352 71356 71566
rect 71956 71738 72014 71952
rect 71956 71566 71968 71738
rect 72002 71566 72014 71738
rect 71956 71352 72014 71566
rect 72614 71738 72672 71952
rect 72614 71566 72626 71738
rect 72660 71566 72672 71738
rect 72614 71352 72672 71566
rect 73272 71738 73330 71952
rect 73272 71566 73284 71738
rect 73318 71566 73330 71738
rect 73272 71352 73330 71566
rect 73930 71738 73988 71952
rect 73930 71566 73942 71738
rect 73976 71566 73988 71738
rect 73930 71352 73988 71566
rect 71298 71044 71356 71258
rect 71298 70872 71310 71044
rect 71344 70872 71356 71044
rect 71298 70658 71356 70872
rect 71956 71044 72014 71258
rect 71956 70872 71968 71044
rect 72002 70872 72014 71044
rect 71956 70658 72014 70872
rect 72614 71044 72672 71258
rect 72614 70872 72626 71044
rect 72660 70872 72672 71044
rect 72614 70658 72672 70872
rect 73272 71044 73330 71258
rect 73272 70872 73284 71044
rect 73318 70872 73330 71044
rect 73272 70658 73330 70872
rect 73930 71044 73988 71258
rect 73930 70872 73942 71044
rect 73976 70872 73988 71044
rect 73930 70658 73988 70872
rect 71298 70350 71356 70564
rect 71298 70178 71310 70350
rect 71344 70178 71356 70350
rect 71298 69964 71356 70178
rect 71956 70350 72014 70564
rect 71956 70178 71968 70350
rect 72002 70178 72014 70350
rect 71956 69964 72014 70178
rect 72614 70350 72672 70564
rect 72614 70178 72626 70350
rect 72660 70178 72672 70350
rect 72614 69964 72672 70178
rect 73272 70350 73330 70564
rect 73272 70178 73284 70350
rect 73318 70178 73330 70350
rect 73272 69964 73330 70178
rect 73930 70350 73988 70564
rect 73930 70178 73942 70350
rect 73976 70178 73988 70350
rect 75162 72934 75174 73106
rect 75208 72934 75220 73106
rect 75162 72720 75220 72934
rect 75820 73106 75878 73320
rect 75820 72934 75832 73106
rect 75866 72934 75878 73106
rect 75820 72720 75878 72934
rect 76478 73106 76536 73320
rect 76478 72934 76490 73106
rect 76524 72934 76536 73106
rect 76478 72720 76536 72934
rect 77136 73106 77194 73320
rect 77136 72934 77148 73106
rect 77182 72934 77194 73106
rect 77136 72720 77194 72934
rect 77794 73106 77852 73320
rect 79012 73120 79070 73334
rect 77794 72934 77806 73106
rect 77840 72934 77852 73106
rect 77794 72720 77852 72934
rect 75162 72412 75220 72626
rect 75162 72240 75174 72412
rect 75208 72240 75220 72412
rect 75162 72026 75220 72240
rect 75820 72412 75878 72626
rect 75820 72240 75832 72412
rect 75866 72240 75878 72412
rect 75820 72026 75878 72240
rect 76478 72412 76536 72626
rect 76478 72240 76490 72412
rect 76524 72240 76536 72412
rect 76478 72026 76536 72240
rect 77136 72412 77194 72626
rect 77136 72240 77148 72412
rect 77182 72240 77194 72412
rect 77136 72026 77194 72240
rect 77794 72412 77852 72626
rect 77794 72240 77806 72412
rect 77840 72240 77852 72412
rect 77794 72026 77852 72240
rect 75162 71718 75220 71932
rect 75162 71546 75174 71718
rect 75208 71546 75220 71718
rect 75162 71332 75220 71546
rect 75820 71718 75878 71932
rect 75820 71546 75832 71718
rect 75866 71546 75878 71718
rect 75820 71332 75878 71546
rect 76478 71718 76536 71932
rect 76478 71546 76490 71718
rect 76524 71546 76536 71718
rect 76478 71332 76536 71546
rect 77136 71718 77194 71932
rect 77136 71546 77148 71718
rect 77182 71546 77194 71718
rect 77136 71332 77194 71546
rect 77794 71718 77852 71932
rect 77794 71546 77806 71718
rect 77840 71546 77852 71718
rect 77794 71332 77852 71546
rect 75162 71024 75220 71238
rect 75162 70852 75174 71024
rect 75208 70852 75220 71024
rect 75162 70638 75220 70852
rect 75820 71024 75878 71238
rect 75820 70852 75832 71024
rect 75866 70852 75878 71024
rect 75820 70638 75878 70852
rect 76478 71024 76536 71238
rect 76478 70852 76490 71024
rect 76524 70852 76536 71024
rect 76478 70638 76536 70852
rect 77136 71024 77194 71238
rect 77136 70852 77148 71024
rect 77182 70852 77194 71024
rect 77136 70638 77194 70852
rect 77794 71024 77852 71238
rect 77794 70852 77806 71024
rect 77840 70852 77852 71024
rect 77794 70638 77852 70852
rect 75162 70330 75220 70544
rect 73930 69964 73988 70178
rect 75162 70158 75174 70330
rect 75208 70158 75220 70330
rect 75162 69944 75220 70158
rect 75820 70330 75878 70544
rect 75820 70158 75832 70330
rect 75866 70158 75878 70330
rect 75820 69944 75878 70158
rect 76478 70330 76536 70544
rect 76478 70158 76490 70330
rect 76524 70158 76536 70330
rect 76478 69944 76536 70158
rect 77136 70330 77194 70544
rect 77136 70158 77148 70330
rect 77182 70158 77194 70330
rect 77136 69944 77194 70158
rect 77794 70330 77852 70544
rect 77794 70158 77806 70330
rect 77840 70158 77852 70330
rect 79012 72948 79024 73120
rect 79058 72948 79070 73120
rect 79012 72734 79070 72948
rect 79670 73120 79728 73334
rect 79670 72948 79682 73120
rect 79716 72948 79728 73120
rect 79670 72734 79728 72948
rect 80328 73120 80386 73334
rect 80328 72948 80340 73120
rect 80374 72948 80386 73120
rect 80328 72734 80386 72948
rect 80986 73120 81044 73334
rect 80986 72948 80998 73120
rect 81032 72948 81044 73120
rect 80986 72734 81044 72948
rect 81644 73120 81702 73334
rect 81644 72948 81656 73120
rect 81690 72948 81702 73120
rect 81644 72734 81702 72948
rect 79012 72426 79070 72640
rect 79012 72254 79024 72426
rect 79058 72254 79070 72426
rect 79012 72040 79070 72254
rect 79670 72426 79728 72640
rect 79670 72254 79682 72426
rect 79716 72254 79728 72426
rect 79670 72040 79728 72254
rect 80328 72426 80386 72640
rect 80328 72254 80340 72426
rect 80374 72254 80386 72426
rect 80328 72040 80386 72254
rect 80986 72426 81044 72640
rect 80986 72254 80998 72426
rect 81032 72254 81044 72426
rect 80986 72040 81044 72254
rect 81644 72426 81702 72640
rect 81644 72254 81656 72426
rect 81690 72254 81702 72426
rect 81644 72040 81702 72254
rect 79012 71732 79070 71946
rect 79012 71560 79024 71732
rect 79058 71560 79070 71732
rect 79012 71346 79070 71560
rect 79670 71732 79728 71946
rect 79670 71560 79682 71732
rect 79716 71560 79728 71732
rect 79670 71346 79728 71560
rect 80328 71732 80386 71946
rect 80328 71560 80340 71732
rect 80374 71560 80386 71732
rect 80328 71346 80386 71560
rect 80986 71732 81044 71946
rect 80986 71560 80998 71732
rect 81032 71560 81044 71732
rect 80986 71346 81044 71560
rect 81644 71732 81702 71946
rect 81644 71560 81656 71732
rect 81690 71560 81702 71732
rect 81644 71346 81702 71560
rect 79012 71038 79070 71252
rect 79012 70866 79024 71038
rect 79058 70866 79070 71038
rect 79012 70652 79070 70866
rect 79670 71038 79728 71252
rect 79670 70866 79682 71038
rect 79716 70866 79728 71038
rect 79670 70652 79728 70866
rect 80328 71038 80386 71252
rect 80328 70866 80340 71038
rect 80374 70866 80386 71038
rect 80328 70652 80386 70866
rect 80986 71038 81044 71252
rect 80986 70866 80998 71038
rect 81032 70866 81044 71038
rect 80986 70652 81044 70866
rect 81644 71038 81702 71252
rect 81644 70866 81656 71038
rect 81690 70866 81702 71038
rect 81644 70652 81702 70866
rect 79012 70344 79070 70558
rect 77794 69944 77852 70158
rect 79012 70172 79024 70344
rect 79058 70172 79070 70344
rect 79012 69958 79070 70172
rect 79670 70344 79728 70558
rect 79670 70172 79682 70344
rect 79716 70172 79728 70344
rect 79670 69958 79728 70172
rect 80328 70344 80386 70558
rect 80328 70172 80340 70344
rect 80374 70172 80386 70344
rect 80328 69958 80386 70172
rect 80986 70344 81044 70558
rect 80986 70172 80998 70344
rect 81032 70172 81044 70344
rect 80986 69958 81044 70172
rect 81644 70344 81702 70558
rect 81644 70172 81656 70344
rect 81690 70172 81702 70344
rect 81644 69958 81702 70172
rect 71294 69350 71352 69564
rect 42188 68372 42788 68384
rect 42188 68338 42402 68372
rect 42574 68338 42788 68372
rect 42188 68326 42788 68338
rect 42882 68372 43482 68384
rect 42882 68338 43096 68372
rect 43268 68338 43482 68372
rect 42882 68326 43482 68338
rect 43576 68372 44176 68384
rect 43576 68338 43790 68372
rect 43962 68338 44176 68372
rect 43576 68326 44176 68338
rect 44270 68372 44870 68384
rect 44270 68338 44484 68372
rect 44656 68338 44870 68372
rect 44270 68326 44870 68338
rect 44964 68372 45564 68384
rect 44964 68338 45178 68372
rect 45350 68338 45564 68372
rect 44964 68326 45564 68338
rect 46182 68372 46782 68384
rect 46182 68338 46396 68372
rect 46568 68338 46782 68372
rect 46182 68326 46782 68338
rect 46876 68372 47476 68384
rect 46876 68338 47090 68372
rect 47262 68338 47476 68372
rect 46876 68326 47476 68338
rect 47570 68372 48170 68384
rect 47570 68338 47784 68372
rect 47956 68338 48170 68372
rect 47570 68326 48170 68338
rect 48264 68372 48864 68384
rect 48264 68338 48478 68372
rect 48650 68338 48864 68372
rect 48264 68326 48864 68338
rect 48958 68372 49558 68384
rect 48958 68338 49172 68372
rect 49344 68338 49558 68372
rect 48958 68326 49558 68338
rect 50204 68372 50804 68384
rect 50204 68338 50418 68372
rect 50590 68338 50804 68372
rect 50204 68326 50804 68338
rect 50898 68372 51498 68384
rect 50898 68338 51112 68372
rect 51284 68338 51498 68372
rect 50898 68326 51498 68338
rect 51592 68372 52192 68384
rect 51592 68338 51806 68372
rect 51978 68338 52192 68372
rect 51592 68326 52192 68338
rect 52286 68372 52886 68384
rect 52286 68338 52500 68372
rect 52672 68338 52886 68372
rect 52286 68326 52886 68338
rect 52980 68372 53580 68384
rect 52980 68338 53194 68372
rect 53366 68338 53580 68372
rect 52980 68326 53580 68338
rect 54226 68372 54826 68384
rect 54226 68338 54440 68372
rect 54612 68338 54826 68372
rect 54226 68326 54826 68338
rect 54920 68372 55520 68384
rect 54920 68338 55134 68372
rect 55306 68338 55520 68372
rect 54920 68326 55520 68338
rect 55614 68372 56214 68384
rect 55614 68338 55828 68372
rect 56000 68338 56214 68372
rect 55614 68326 56214 68338
rect 56308 68372 56908 68384
rect 56308 68338 56522 68372
rect 56694 68338 56908 68372
rect 56308 68326 56908 68338
rect 57002 68372 57602 68384
rect 57002 68338 57216 68372
rect 57388 68338 57602 68372
rect 57002 68326 57602 68338
rect 42188 67714 42788 67726
rect 42188 67680 42402 67714
rect 42574 67680 42788 67714
rect 42188 67668 42788 67680
rect 42882 67714 43482 67726
rect 42882 67680 43096 67714
rect 43268 67680 43482 67714
rect 42882 67668 43482 67680
rect 43576 67714 44176 67726
rect 43576 67680 43790 67714
rect 43962 67680 44176 67714
rect 43576 67668 44176 67680
rect 44270 67714 44870 67726
rect 44270 67680 44484 67714
rect 44656 67680 44870 67714
rect 44270 67668 44870 67680
rect 44964 67714 45564 67726
rect 44964 67680 45178 67714
rect 45350 67680 45564 67714
rect 44964 67668 45564 67680
rect 46182 67714 46782 67726
rect 46182 67680 46396 67714
rect 46568 67680 46782 67714
rect 46182 67668 46782 67680
rect 46876 67714 47476 67726
rect 46876 67680 47090 67714
rect 47262 67680 47476 67714
rect 46876 67668 47476 67680
rect 47570 67714 48170 67726
rect 47570 67680 47784 67714
rect 47956 67680 48170 67714
rect 47570 67668 48170 67680
rect 48264 67714 48864 67726
rect 48264 67680 48478 67714
rect 48650 67680 48864 67714
rect 48264 67668 48864 67680
rect 48958 67714 49558 67726
rect 48958 67680 49172 67714
rect 49344 67680 49558 67714
rect 48958 67668 49558 67680
rect 50204 67714 50804 67726
rect 50204 67680 50418 67714
rect 50590 67680 50804 67714
rect 50204 67668 50804 67680
rect 50898 67714 51498 67726
rect 50898 67680 51112 67714
rect 51284 67680 51498 67714
rect 50898 67668 51498 67680
rect 51592 67714 52192 67726
rect 51592 67680 51806 67714
rect 51978 67680 52192 67714
rect 51592 67668 52192 67680
rect 52286 67714 52886 67726
rect 52286 67680 52500 67714
rect 52672 67680 52886 67714
rect 52286 67668 52886 67680
rect 52980 67714 53580 67726
rect 52980 67680 53194 67714
rect 53366 67680 53580 67714
rect 52980 67668 53580 67680
rect 54226 67714 54826 67726
rect 54226 67680 54440 67714
rect 54612 67680 54826 67714
rect 54226 67668 54826 67680
rect 54920 67714 55520 67726
rect 54920 67680 55134 67714
rect 55306 67680 55520 67714
rect 54920 67668 55520 67680
rect 55614 67714 56214 67726
rect 55614 67680 55828 67714
rect 56000 67680 56214 67714
rect 55614 67668 56214 67680
rect 56308 67714 56908 67726
rect 56308 67680 56522 67714
rect 56694 67680 56908 67714
rect 56308 67668 56908 67680
rect 57002 67714 57602 67726
rect 57002 67680 57216 67714
rect 57388 67680 57602 67714
rect 57002 67668 57602 67680
rect 42188 67056 42788 67068
rect 42188 67022 42402 67056
rect 42574 67022 42788 67056
rect 42188 67010 42788 67022
rect 42882 67056 43482 67068
rect 42882 67022 43096 67056
rect 43268 67022 43482 67056
rect 42882 67010 43482 67022
rect 43576 67056 44176 67068
rect 43576 67022 43790 67056
rect 43962 67022 44176 67056
rect 43576 67010 44176 67022
rect 44270 67056 44870 67068
rect 44270 67022 44484 67056
rect 44656 67022 44870 67056
rect 44270 67010 44870 67022
rect 44964 67056 45564 67068
rect 44964 67022 45178 67056
rect 45350 67022 45564 67056
rect 44964 67010 45564 67022
rect 46182 67056 46782 67068
rect 46182 67022 46396 67056
rect 46568 67022 46782 67056
rect 46182 67010 46782 67022
rect 46876 67056 47476 67068
rect 46876 67022 47090 67056
rect 47262 67022 47476 67056
rect 46876 67010 47476 67022
rect 47570 67056 48170 67068
rect 47570 67022 47784 67056
rect 47956 67022 48170 67056
rect 47570 67010 48170 67022
rect 48264 67056 48864 67068
rect 48264 67022 48478 67056
rect 48650 67022 48864 67056
rect 48264 67010 48864 67022
rect 48958 67056 49558 67068
rect 48958 67022 49172 67056
rect 49344 67022 49558 67056
rect 48958 67010 49558 67022
rect 50204 67056 50804 67068
rect 50204 67022 50418 67056
rect 50590 67022 50804 67056
rect 50204 67010 50804 67022
rect 50898 67056 51498 67068
rect 50898 67022 51112 67056
rect 51284 67022 51498 67056
rect 50898 67010 51498 67022
rect 51592 67056 52192 67068
rect 51592 67022 51806 67056
rect 51978 67022 52192 67056
rect 51592 67010 52192 67022
rect 52286 67056 52886 67068
rect 52286 67022 52500 67056
rect 52672 67022 52886 67056
rect 52286 67010 52886 67022
rect 52980 67056 53580 67068
rect 52980 67022 53194 67056
rect 53366 67022 53580 67056
rect 52980 67010 53580 67022
rect 54226 67056 54826 67068
rect 54226 67022 54440 67056
rect 54612 67022 54826 67056
rect 54226 67010 54826 67022
rect 54920 67056 55520 67068
rect 54920 67022 55134 67056
rect 55306 67022 55520 67056
rect 54920 67010 55520 67022
rect 55614 67056 56214 67068
rect 55614 67022 55828 67056
rect 56000 67022 56214 67056
rect 55614 67010 56214 67022
rect 56308 67056 56908 67068
rect 56308 67022 56522 67056
rect 56694 67022 56908 67056
rect 56308 67010 56908 67022
rect 57002 67056 57602 67068
rect 57002 67022 57216 67056
rect 57388 67022 57602 67056
rect 57002 67010 57602 67022
rect 42188 66398 42788 66410
rect 42188 66364 42402 66398
rect 42574 66364 42788 66398
rect 42188 66352 42788 66364
rect 42882 66398 43482 66410
rect 42882 66364 43096 66398
rect 43268 66364 43482 66398
rect 42882 66352 43482 66364
rect 43576 66398 44176 66410
rect 43576 66364 43790 66398
rect 43962 66364 44176 66398
rect 43576 66352 44176 66364
rect 44270 66398 44870 66410
rect 44270 66364 44484 66398
rect 44656 66364 44870 66398
rect 44270 66352 44870 66364
rect 44964 66398 45564 66410
rect 44964 66364 45178 66398
rect 45350 66364 45564 66398
rect 44964 66352 45564 66364
rect 46182 66398 46782 66410
rect 46182 66364 46396 66398
rect 46568 66364 46782 66398
rect 46182 66352 46782 66364
rect 46876 66398 47476 66410
rect 46876 66364 47090 66398
rect 47262 66364 47476 66398
rect 46876 66352 47476 66364
rect 47570 66398 48170 66410
rect 47570 66364 47784 66398
rect 47956 66364 48170 66398
rect 47570 66352 48170 66364
rect 48264 66398 48864 66410
rect 48264 66364 48478 66398
rect 48650 66364 48864 66398
rect 48264 66352 48864 66364
rect 48958 66398 49558 66410
rect 48958 66364 49172 66398
rect 49344 66364 49558 66398
rect 48958 66352 49558 66364
rect 50204 66398 50804 66410
rect 50204 66364 50418 66398
rect 50590 66364 50804 66398
rect 50204 66352 50804 66364
rect 50898 66398 51498 66410
rect 50898 66364 51112 66398
rect 51284 66364 51498 66398
rect 50898 66352 51498 66364
rect 51592 66398 52192 66410
rect 51592 66364 51806 66398
rect 51978 66364 52192 66398
rect 51592 66352 52192 66364
rect 52286 66398 52886 66410
rect 52286 66364 52500 66398
rect 52672 66364 52886 66398
rect 52286 66352 52886 66364
rect 52980 66398 53580 66410
rect 52980 66364 53194 66398
rect 53366 66364 53580 66398
rect 52980 66352 53580 66364
rect 54226 66398 54826 66410
rect 54226 66364 54440 66398
rect 54612 66364 54826 66398
rect 54226 66352 54826 66364
rect 54920 66398 55520 66410
rect 54920 66364 55134 66398
rect 55306 66364 55520 66398
rect 54920 66352 55520 66364
rect 55614 66398 56214 66410
rect 55614 66364 55828 66398
rect 56000 66364 56214 66398
rect 55614 66352 56214 66364
rect 56308 66398 56908 66410
rect 56308 66364 56522 66398
rect 56694 66364 56908 66398
rect 56308 66352 56908 66364
rect 57002 66398 57602 66410
rect 57002 66364 57216 66398
rect 57388 66364 57602 66398
rect 57002 66352 57602 66364
rect 71294 69178 71306 69350
rect 71340 69178 71352 69350
rect 71294 68964 71352 69178
rect 71952 69350 72010 69564
rect 71952 69178 71964 69350
rect 71998 69178 72010 69350
rect 71952 68964 72010 69178
rect 72610 69350 72668 69564
rect 72610 69178 72622 69350
rect 72656 69178 72668 69350
rect 72610 68964 72668 69178
rect 73268 69350 73326 69564
rect 73268 69178 73280 69350
rect 73314 69178 73326 69350
rect 73268 68964 73326 69178
rect 73926 69350 73984 69564
rect 73926 69178 73938 69350
rect 73972 69178 73984 69350
rect 75158 69330 75216 69544
rect 73926 68964 73984 69178
rect 71294 68656 71352 68870
rect 71294 68484 71306 68656
rect 71340 68484 71352 68656
rect 71294 68270 71352 68484
rect 71952 68656 72010 68870
rect 71952 68484 71964 68656
rect 71998 68484 72010 68656
rect 71952 68270 72010 68484
rect 72610 68656 72668 68870
rect 72610 68484 72622 68656
rect 72656 68484 72668 68656
rect 72610 68270 72668 68484
rect 73268 68656 73326 68870
rect 73268 68484 73280 68656
rect 73314 68484 73326 68656
rect 73268 68270 73326 68484
rect 73926 68656 73984 68870
rect 73926 68484 73938 68656
rect 73972 68484 73984 68656
rect 73926 68270 73984 68484
rect 71294 67962 71352 68176
rect 71294 67790 71306 67962
rect 71340 67790 71352 67962
rect 71294 67576 71352 67790
rect 71952 67962 72010 68176
rect 71952 67790 71964 67962
rect 71998 67790 72010 67962
rect 71952 67576 72010 67790
rect 72610 67962 72668 68176
rect 72610 67790 72622 67962
rect 72656 67790 72668 67962
rect 72610 67576 72668 67790
rect 73268 67962 73326 68176
rect 73268 67790 73280 67962
rect 73314 67790 73326 67962
rect 73268 67576 73326 67790
rect 73926 67962 73984 68176
rect 73926 67790 73938 67962
rect 73972 67790 73984 67962
rect 73926 67576 73984 67790
rect 71294 67268 71352 67482
rect 71294 67096 71306 67268
rect 71340 67096 71352 67268
rect 71294 66882 71352 67096
rect 71952 67268 72010 67482
rect 71952 67096 71964 67268
rect 71998 67096 72010 67268
rect 71952 66882 72010 67096
rect 72610 67268 72668 67482
rect 72610 67096 72622 67268
rect 72656 67096 72668 67268
rect 72610 66882 72668 67096
rect 73268 67268 73326 67482
rect 73268 67096 73280 67268
rect 73314 67096 73326 67268
rect 73268 66882 73326 67096
rect 73926 67268 73984 67482
rect 73926 67096 73938 67268
rect 73972 67096 73984 67268
rect 73926 66882 73984 67096
rect 71294 66574 71352 66788
rect 19358 65620 19958 65632
rect 752 65570 1352 65582
rect 752 65536 966 65570
rect 1138 65536 1352 65570
rect 752 65524 1352 65536
rect 1446 65570 2046 65582
rect 1446 65536 1660 65570
rect 1832 65536 2046 65570
rect 1446 65524 2046 65536
rect 2140 65570 2740 65582
rect 2140 65536 2354 65570
rect 2526 65536 2740 65570
rect 2140 65524 2740 65536
rect 3420 65566 4020 65578
rect 3420 65532 3634 65566
rect 3806 65532 4020 65566
rect 3420 65520 4020 65532
rect 4114 65566 4714 65578
rect 4114 65532 4328 65566
rect 4500 65532 4714 65566
rect 4114 65520 4714 65532
rect 4808 65566 5408 65578
rect 4808 65532 5022 65566
rect 5194 65532 5408 65566
rect 4808 65520 5408 65532
rect 6094 65572 6694 65584
rect 6094 65538 6308 65572
rect 6480 65538 6694 65572
rect 6094 65526 6694 65538
rect 6788 65572 7388 65584
rect 6788 65538 7002 65572
rect 7174 65538 7388 65572
rect 6788 65526 7388 65538
rect 7482 65572 8082 65584
rect 7482 65538 7696 65572
rect 7868 65538 8082 65572
rect 7482 65526 8082 65538
rect 8740 65572 9340 65584
rect 8740 65538 8954 65572
rect 9126 65538 9340 65572
rect 8740 65526 9340 65538
rect 9434 65572 10034 65584
rect 9434 65538 9648 65572
rect 9820 65538 10034 65572
rect 9434 65526 10034 65538
rect 10128 65572 10728 65584
rect 10128 65538 10342 65572
rect 10514 65538 10728 65572
rect 10128 65526 10728 65538
rect 11394 65566 11994 65578
rect 11394 65532 11608 65566
rect 11780 65532 11994 65566
rect 752 64912 1352 64924
rect 752 64878 966 64912
rect 1138 64878 1352 64912
rect 752 64866 1352 64878
rect 1446 64912 2046 64924
rect 1446 64878 1660 64912
rect 1832 64878 2046 64912
rect 1446 64866 2046 64878
rect 2140 64912 2740 64924
rect 2140 64878 2354 64912
rect 2526 64878 2740 64912
rect 2140 64866 2740 64878
rect 11394 65520 11994 65532
rect 12088 65566 12688 65578
rect 12088 65532 12302 65566
rect 12474 65532 12688 65566
rect 12088 65520 12688 65532
rect 12782 65566 13382 65578
rect 12782 65532 12996 65566
rect 13168 65532 13382 65566
rect 12782 65520 13382 65532
rect 14048 65572 14648 65584
rect 14048 65538 14262 65572
rect 14434 65538 14648 65572
rect 14048 65526 14648 65538
rect 14742 65572 15342 65584
rect 14742 65538 14956 65572
rect 15128 65538 15342 65572
rect 14742 65526 15342 65538
rect 15436 65572 16036 65584
rect 15436 65538 15650 65572
rect 15822 65538 16036 65572
rect 15436 65526 16036 65538
rect 16674 65576 17274 65588
rect 16674 65542 16888 65576
rect 17060 65542 17274 65576
rect 16674 65530 17274 65542
rect 17368 65576 17968 65588
rect 17368 65542 17582 65576
rect 17754 65542 17968 65576
rect 17368 65530 17968 65542
rect 18062 65576 18662 65588
rect 18062 65542 18276 65576
rect 18448 65542 18662 65576
rect 19358 65586 19572 65620
rect 19744 65586 19958 65620
rect 19358 65574 19958 65586
rect 20052 65620 20652 65632
rect 20052 65586 20266 65620
rect 20438 65586 20652 65620
rect 20052 65574 20652 65586
rect 18062 65530 18662 65542
rect 3420 64908 4020 64920
rect 3420 64874 3634 64908
rect 3806 64874 4020 64908
rect 3420 64862 4020 64874
rect 4114 64908 4714 64920
rect 4114 64874 4328 64908
rect 4500 64874 4714 64908
rect 4114 64862 4714 64874
rect 4808 64908 5408 64920
rect 4808 64874 5022 64908
rect 5194 64874 5408 64908
rect 4808 64862 5408 64874
rect 6094 64914 6694 64926
rect 6094 64880 6308 64914
rect 6480 64880 6694 64914
rect 6094 64868 6694 64880
rect 6788 64914 7388 64926
rect 6788 64880 7002 64914
rect 7174 64880 7388 64914
rect 6788 64868 7388 64880
rect 7482 64914 8082 64926
rect 7482 64880 7696 64914
rect 7868 64880 8082 64914
rect 7482 64868 8082 64880
rect 8740 64914 9340 64926
rect 8740 64880 8954 64914
rect 9126 64880 9340 64914
rect 8740 64868 9340 64880
rect 9434 64914 10034 64926
rect 9434 64880 9648 64914
rect 9820 64880 10034 64914
rect 9434 64868 10034 64880
rect 10128 64914 10728 64926
rect 10128 64880 10342 64914
rect 10514 64880 10728 64914
rect 10128 64868 10728 64880
rect 752 64254 1352 64266
rect 752 64220 966 64254
rect 1138 64220 1352 64254
rect 752 64208 1352 64220
rect 1446 64254 2046 64266
rect 1446 64220 1660 64254
rect 1832 64220 2046 64254
rect 1446 64208 2046 64220
rect 2140 64254 2740 64266
rect 2140 64220 2354 64254
rect 2526 64220 2740 64254
rect 2140 64208 2740 64220
rect 11394 64908 11994 64920
rect 11394 64874 11608 64908
rect 11780 64874 11994 64908
rect 11394 64862 11994 64874
rect 12088 64908 12688 64920
rect 12088 64874 12302 64908
rect 12474 64874 12688 64908
rect 12088 64862 12688 64874
rect 12782 64908 13382 64920
rect 12782 64874 12996 64908
rect 13168 64874 13382 64908
rect 12782 64862 13382 64874
rect 14048 64914 14648 64926
rect 14048 64880 14262 64914
rect 14434 64880 14648 64914
rect 14048 64868 14648 64880
rect 14742 64914 15342 64926
rect 14742 64880 14956 64914
rect 15128 64880 15342 64914
rect 14742 64868 15342 64880
rect 15436 64914 16036 64926
rect 15436 64880 15650 64914
rect 15822 64880 16036 64914
rect 15436 64868 16036 64880
rect 16674 64918 17274 64930
rect 16674 64884 16888 64918
rect 17060 64884 17274 64918
rect 16674 64872 17274 64884
rect 17368 64918 17968 64930
rect 17368 64884 17582 64918
rect 17754 64884 17968 64918
rect 17368 64872 17968 64884
rect 18062 64918 18662 64930
rect 18062 64884 18276 64918
rect 18448 64884 18662 64918
rect 18062 64872 18662 64884
rect 19358 64962 19958 64974
rect 19358 64928 19572 64962
rect 19744 64928 19958 64962
rect 19358 64916 19958 64928
rect 20052 64962 20652 64974
rect 20052 64928 20266 64962
rect 20438 64928 20652 64962
rect 20052 64916 20652 64928
rect 3420 64250 4020 64262
rect 3420 64216 3634 64250
rect 3806 64216 4020 64250
rect 3420 64204 4020 64216
rect 4114 64250 4714 64262
rect 4114 64216 4328 64250
rect 4500 64216 4714 64250
rect 4114 64204 4714 64216
rect 4808 64250 5408 64262
rect 4808 64216 5022 64250
rect 5194 64216 5408 64250
rect 4808 64204 5408 64216
rect 6094 64256 6694 64268
rect 6094 64222 6308 64256
rect 6480 64222 6694 64256
rect 6094 64210 6694 64222
rect 6788 64256 7388 64268
rect 6788 64222 7002 64256
rect 7174 64222 7388 64256
rect 6788 64210 7388 64222
rect 7482 64256 8082 64268
rect 7482 64222 7696 64256
rect 7868 64222 8082 64256
rect 7482 64210 8082 64222
rect 8740 64256 9340 64268
rect 8740 64222 8954 64256
rect 9126 64222 9340 64256
rect 8740 64210 9340 64222
rect 9434 64256 10034 64268
rect 9434 64222 9648 64256
rect 9820 64222 10034 64256
rect 9434 64210 10034 64222
rect 10128 64256 10728 64268
rect 10128 64222 10342 64256
rect 10514 64222 10728 64256
rect 10128 64210 10728 64222
rect 752 63596 1352 63608
rect 752 63562 966 63596
rect 1138 63562 1352 63596
rect 752 63550 1352 63562
rect 1446 63596 2046 63608
rect 1446 63562 1660 63596
rect 1832 63562 2046 63596
rect 1446 63550 2046 63562
rect 2140 63596 2740 63608
rect 2140 63562 2354 63596
rect 2526 63562 2740 63596
rect 2140 63550 2740 63562
rect 11394 64250 11994 64262
rect 11394 64216 11608 64250
rect 11780 64216 11994 64250
rect 11394 64204 11994 64216
rect 12088 64250 12688 64262
rect 12088 64216 12302 64250
rect 12474 64216 12688 64250
rect 12088 64204 12688 64216
rect 12782 64250 13382 64262
rect 12782 64216 12996 64250
rect 13168 64216 13382 64250
rect 12782 64204 13382 64216
rect 14048 64256 14648 64268
rect 14048 64222 14262 64256
rect 14434 64222 14648 64256
rect 14048 64210 14648 64222
rect 14742 64256 15342 64268
rect 14742 64222 14956 64256
rect 15128 64222 15342 64256
rect 14742 64210 15342 64222
rect 15436 64256 16036 64268
rect 15436 64222 15650 64256
rect 15822 64222 16036 64256
rect 15436 64210 16036 64222
rect 16674 64260 17274 64272
rect 16674 64226 16888 64260
rect 17060 64226 17274 64260
rect 16674 64214 17274 64226
rect 17368 64260 17968 64272
rect 17368 64226 17582 64260
rect 17754 64226 17968 64260
rect 17368 64214 17968 64226
rect 18062 64260 18662 64272
rect 18062 64226 18276 64260
rect 18448 64226 18662 64260
rect 18062 64214 18662 64226
rect 19358 64304 19958 64316
rect 19358 64270 19572 64304
rect 19744 64270 19958 64304
rect 19358 64258 19958 64270
rect 20052 64304 20652 64316
rect 20052 64270 20266 64304
rect 20438 64270 20652 64304
rect 20052 64258 20652 64270
rect 3420 63592 4020 63604
rect 3420 63558 3634 63592
rect 3806 63558 4020 63592
rect 3420 63546 4020 63558
rect 4114 63592 4714 63604
rect 4114 63558 4328 63592
rect 4500 63558 4714 63592
rect 4114 63546 4714 63558
rect 4808 63592 5408 63604
rect 4808 63558 5022 63592
rect 5194 63558 5408 63592
rect 4808 63546 5408 63558
rect 6094 63598 6694 63610
rect 6094 63564 6308 63598
rect 6480 63564 6694 63598
rect 6094 63552 6694 63564
rect 6788 63598 7388 63610
rect 6788 63564 7002 63598
rect 7174 63564 7388 63598
rect 6788 63552 7388 63564
rect 7482 63598 8082 63610
rect 7482 63564 7696 63598
rect 7868 63564 8082 63598
rect 7482 63552 8082 63564
rect 8740 63598 9340 63610
rect 8740 63564 8954 63598
rect 9126 63564 9340 63598
rect 8740 63552 9340 63564
rect 9434 63598 10034 63610
rect 9434 63564 9648 63598
rect 9820 63564 10034 63598
rect 9434 63552 10034 63564
rect 10128 63598 10728 63610
rect 10128 63564 10342 63598
rect 10514 63564 10728 63598
rect 10128 63552 10728 63564
rect 752 62938 1352 62950
rect 752 62904 966 62938
rect 1138 62904 1352 62938
rect 752 62892 1352 62904
rect 1446 62938 2046 62950
rect 1446 62904 1660 62938
rect 1832 62904 2046 62938
rect 1446 62892 2046 62904
rect 2140 62938 2740 62950
rect 2140 62904 2354 62938
rect 2526 62904 2740 62938
rect 2140 62892 2740 62904
rect 11394 63592 11994 63604
rect 11394 63558 11608 63592
rect 11780 63558 11994 63592
rect 11394 63546 11994 63558
rect 12088 63592 12688 63604
rect 12088 63558 12302 63592
rect 12474 63558 12688 63592
rect 12088 63546 12688 63558
rect 12782 63592 13382 63604
rect 12782 63558 12996 63592
rect 13168 63558 13382 63592
rect 12782 63546 13382 63558
rect 14048 63598 14648 63610
rect 14048 63564 14262 63598
rect 14434 63564 14648 63598
rect 14048 63552 14648 63564
rect 14742 63598 15342 63610
rect 14742 63564 14956 63598
rect 15128 63564 15342 63598
rect 14742 63552 15342 63564
rect 15436 63598 16036 63610
rect 15436 63564 15650 63598
rect 15822 63564 16036 63598
rect 15436 63552 16036 63564
rect 16674 63602 17274 63614
rect 16674 63568 16888 63602
rect 17060 63568 17274 63602
rect 16674 63556 17274 63568
rect 17368 63602 17968 63614
rect 17368 63568 17582 63602
rect 17754 63568 17968 63602
rect 17368 63556 17968 63568
rect 18062 63602 18662 63614
rect 18062 63568 18276 63602
rect 18448 63568 18662 63602
rect 18062 63556 18662 63568
rect 19358 63646 19958 63658
rect 19358 63612 19572 63646
rect 19744 63612 19958 63646
rect 19358 63600 19958 63612
rect 20052 63646 20652 63658
rect 20052 63612 20266 63646
rect 20438 63612 20652 63646
rect 20052 63600 20652 63612
rect 3420 62934 4020 62946
rect 3420 62900 3634 62934
rect 3806 62900 4020 62934
rect 3420 62888 4020 62900
rect 4114 62934 4714 62946
rect 4114 62900 4328 62934
rect 4500 62900 4714 62934
rect 4114 62888 4714 62900
rect 4808 62934 5408 62946
rect 4808 62900 5022 62934
rect 5194 62900 5408 62934
rect 4808 62888 5408 62900
rect 6094 62940 6694 62952
rect 6094 62906 6308 62940
rect 6480 62906 6694 62940
rect 6094 62894 6694 62906
rect 6788 62940 7388 62952
rect 6788 62906 7002 62940
rect 7174 62906 7388 62940
rect 6788 62894 7388 62906
rect 7482 62940 8082 62952
rect 7482 62906 7696 62940
rect 7868 62906 8082 62940
rect 7482 62894 8082 62906
rect 8740 62940 9340 62952
rect 8740 62906 8954 62940
rect 9126 62906 9340 62940
rect 8740 62894 9340 62906
rect 9434 62940 10034 62952
rect 9434 62906 9648 62940
rect 9820 62906 10034 62940
rect 9434 62894 10034 62906
rect 10128 62940 10728 62952
rect 10128 62906 10342 62940
rect 10514 62906 10728 62940
rect 10128 62894 10728 62906
rect 752 62280 1352 62292
rect 752 62246 966 62280
rect 1138 62246 1352 62280
rect 752 62234 1352 62246
rect 1446 62280 2046 62292
rect 1446 62246 1660 62280
rect 1832 62246 2046 62280
rect 1446 62234 2046 62246
rect 2140 62280 2740 62292
rect 2140 62246 2354 62280
rect 2526 62246 2740 62280
rect 2140 62234 2740 62246
rect 11394 62934 11994 62946
rect 11394 62900 11608 62934
rect 11780 62900 11994 62934
rect 11394 62888 11994 62900
rect 12088 62934 12688 62946
rect 12088 62900 12302 62934
rect 12474 62900 12688 62934
rect 12088 62888 12688 62900
rect 12782 62934 13382 62946
rect 12782 62900 12996 62934
rect 13168 62900 13382 62934
rect 12782 62888 13382 62900
rect 14048 62940 14648 62952
rect 14048 62906 14262 62940
rect 14434 62906 14648 62940
rect 14048 62894 14648 62906
rect 14742 62940 15342 62952
rect 14742 62906 14956 62940
rect 15128 62906 15342 62940
rect 14742 62894 15342 62906
rect 15436 62940 16036 62952
rect 15436 62906 15650 62940
rect 15822 62906 16036 62940
rect 15436 62894 16036 62906
rect 16674 62944 17274 62956
rect 16674 62910 16888 62944
rect 17060 62910 17274 62944
rect 16674 62898 17274 62910
rect 17368 62944 17968 62956
rect 17368 62910 17582 62944
rect 17754 62910 17968 62944
rect 17368 62898 17968 62910
rect 18062 62944 18662 62956
rect 18062 62910 18276 62944
rect 18448 62910 18662 62944
rect 18062 62898 18662 62910
rect 19358 62988 19958 63000
rect 19358 62954 19572 62988
rect 19744 62954 19958 62988
rect 19358 62942 19958 62954
rect 20052 62988 20652 63000
rect 20052 62954 20266 62988
rect 20438 62954 20652 62988
rect 20052 62942 20652 62954
rect 3420 62276 4020 62288
rect 3420 62242 3634 62276
rect 3806 62242 4020 62276
rect 3420 62230 4020 62242
rect 4114 62276 4714 62288
rect 4114 62242 4328 62276
rect 4500 62242 4714 62276
rect 4114 62230 4714 62242
rect 4808 62276 5408 62288
rect 4808 62242 5022 62276
rect 5194 62242 5408 62276
rect 4808 62230 5408 62242
rect 6094 62282 6694 62294
rect 6094 62248 6308 62282
rect 6480 62248 6694 62282
rect 6094 62236 6694 62248
rect 6788 62282 7388 62294
rect 6788 62248 7002 62282
rect 7174 62248 7388 62282
rect 6788 62236 7388 62248
rect 7482 62282 8082 62294
rect 7482 62248 7696 62282
rect 7868 62248 8082 62282
rect 7482 62236 8082 62248
rect 8740 62282 9340 62294
rect 8740 62248 8954 62282
rect 9126 62248 9340 62282
rect 8740 62236 9340 62248
rect 9434 62282 10034 62294
rect 9434 62248 9648 62282
rect 9820 62248 10034 62282
rect 9434 62236 10034 62248
rect 10128 62282 10728 62294
rect 10128 62248 10342 62282
rect 10514 62248 10728 62282
rect 10128 62236 10728 62248
rect 752 61622 1352 61634
rect 752 61588 966 61622
rect 1138 61588 1352 61622
rect 752 61576 1352 61588
rect 1446 61622 2046 61634
rect 1446 61588 1660 61622
rect 1832 61588 2046 61622
rect 1446 61576 2046 61588
rect 2140 61622 2740 61634
rect 2140 61588 2354 61622
rect 2526 61588 2740 61622
rect 2140 61576 2740 61588
rect 11394 62276 11994 62288
rect 11394 62242 11608 62276
rect 11780 62242 11994 62276
rect 11394 62230 11994 62242
rect 12088 62276 12688 62288
rect 12088 62242 12302 62276
rect 12474 62242 12688 62276
rect 12088 62230 12688 62242
rect 12782 62276 13382 62288
rect 12782 62242 12996 62276
rect 13168 62242 13382 62276
rect 12782 62230 13382 62242
rect 14048 62282 14648 62294
rect 14048 62248 14262 62282
rect 14434 62248 14648 62282
rect 14048 62236 14648 62248
rect 14742 62282 15342 62294
rect 14742 62248 14956 62282
rect 15128 62248 15342 62282
rect 14742 62236 15342 62248
rect 15436 62282 16036 62294
rect 15436 62248 15650 62282
rect 15822 62248 16036 62282
rect 15436 62236 16036 62248
rect 16674 62286 17274 62298
rect 16674 62252 16888 62286
rect 17060 62252 17274 62286
rect 16674 62240 17274 62252
rect 17368 62286 17968 62298
rect 17368 62252 17582 62286
rect 17754 62252 17968 62286
rect 17368 62240 17968 62252
rect 18062 62286 18662 62298
rect 18062 62252 18276 62286
rect 18448 62252 18662 62286
rect 18062 62240 18662 62252
rect 19358 62330 19958 62342
rect 19358 62296 19572 62330
rect 19744 62296 19958 62330
rect 19358 62284 19958 62296
rect 20052 62330 20652 62342
rect 20052 62296 20266 62330
rect 20438 62296 20652 62330
rect 20052 62284 20652 62296
rect 3420 61618 4020 61630
rect 3420 61584 3634 61618
rect 3806 61584 4020 61618
rect 3420 61572 4020 61584
rect 4114 61618 4714 61630
rect 4114 61584 4328 61618
rect 4500 61584 4714 61618
rect 4114 61572 4714 61584
rect 4808 61618 5408 61630
rect 4808 61584 5022 61618
rect 5194 61584 5408 61618
rect 4808 61572 5408 61584
rect 6094 61624 6694 61636
rect 6094 61590 6308 61624
rect 6480 61590 6694 61624
rect 6094 61578 6694 61590
rect 6788 61624 7388 61636
rect 6788 61590 7002 61624
rect 7174 61590 7388 61624
rect 6788 61578 7388 61590
rect 7482 61624 8082 61636
rect 7482 61590 7696 61624
rect 7868 61590 8082 61624
rect 7482 61578 8082 61590
rect 8740 61624 9340 61636
rect 8740 61590 8954 61624
rect 9126 61590 9340 61624
rect 8740 61578 9340 61590
rect 9434 61624 10034 61636
rect 9434 61590 9648 61624
rect 9820 61590 10034 61624
rect 9434 61578 10034 61590
rect 10128 61624 10728 61636
rect 10128 61590 10342 61624
rect 10514 61590 10728 61624
rect 10128 61578 10728 61590
rect 752 60964 1352 60976
rect 752 60930 966 60964
rect 1138 60930 1352 60964
rect 752 60918 1352 60930
rect 1446 60964 2046 60976
rect 1446 60930 1660 60964
rect 1832 60930 2046 60964
rect 1446 60918 2046 60930
rect 2140 60964 2740 60976
rect 2140 60930 2354 60964
rect 2526 60930 2740 60964
rect 2140 60918 2740 60930
rect 11394 61618 11994 61630
rect 11394 61584 11608 61618
rect 11780 61584 11994 61618
rect 11394 61572 11994 61584
rect 12088 61618 12688 61630
rect 12088 61584 12302 61618
rect 12474 61584 12688 61618
rect 12088 61572 12688 61584
rect 12782 61618 13382 61630
rect 12782 61584 12996 61618
rect 13168 61584 13382 61618
rect 12782 61572 13382 61584
rect 14048 61624 14648 61636
rect 14048 61590 14262 61624
rect 14434 61590 14648 61624
rect 14048 61578 14648 61590
rect 14742 61624 15342 61636
rect 14742 61590 14956 61624
rect 15128 61590 15342 61624
rect 14742 61578 15342 61590
rect 15436 61624 16036 61636
rect 15436 61590 15650 61624
rect 15822 61590 16036 61624
rect 15436 61578 16036 61590
rect 16674 61628 17274 61640
rect 16674 61594 16888 61628
rect 17060 61594 17274 61628
rect 16674 61582 17274 61594
rect 17368 61628 17968 61640
rect 17368 61594 17582 61628
rect 17754 61594 17968 61628
rect 17368 61582 17968 61594
rect 18062 61628 18662 61640
rect 18062 61594 18276 61628
rect 18448 61594 18662 61628
rect 18062 61582 18662 61594
rect 19358 61672 19958 61684
rect 19358 61638 19572 61672
rect 19744 61638 19958 61672
rect 19358 61626 19958 61638
rect 20052 61672 20652 61684
rect 20052 61638 20266 61672
rect 20438 61638 20652 61672
rect 20052 61626 20652 61638
rect 3420 60960 4020 60972
rect 3420 60926 3634 60960
rect 3806 60926 4020 60960
rect 3420 60914 4020 60926
rect 4114 60960 4714 60972
rect 4114 60926 4328 60960
rect 4500 60926 4714 60960
rect 4114 60914 4714 60926
rect 4808 60960 5408 60972
rect 4808 60926 5022 60960
rect 5194 60926 5408 60960
rect 4808 60914 5408 60926
rect 6094 60966 6694 60978
rect 6094 60932 6308 60966
rect 6480 60932 6694 60966
rect 6094 60920 6694 60932
rect 6788 60966 7388 60978
rect 6788 60932 7002 60966
rect 7174 60932 7388 60966
rect 6788 60920 7388 60932
rect 7482 60966 8082 60978
rect 7482 60932 7696 60966
rect 7868 60932 8082 60966
rect 7482 60920 8082 60932
rect 8740 60966 9340 60978
rect 8740 60932 8954 60966
rect 9126 60932 9340 60966
rect 8740 60920 9340 60932
rect 9434 60966 10034 60978
rect 9434 60932 9648 60966
rect 9820 60932 10034 60966
rect 9434 60920 10034 60932
rect 10128 60966 10728 60978
rect 10128 60932 10342 60966
rect 10514 60932 10728 60966
rect 10128 60920 10728 60932
rect 752 60306 1352 60318
rect 752 60272 966 60306
rect 1138 60272 1352 60306
rect 752 60260 1352 60272
rect 1446 60306 2046 60318
rect 1446 60272 1660 60306
rect 1832 60272 2046 60306
rect 1446 60260 2046 60272
rect 2140 60306 2740 60318
rect 11394 60960 11994 60972
rect 11394 60926 11608 60960
rect 11780 60926 11994 60960
rect 11394 60914 11994 60926
rect 12088 60960 12688 60972
rect 12088 60926 12302 60960
rect 12474 60926 12688 60960
rect 12088 60914 12688 60926
rect 12782 60960 13382 60972
rect 12782 60926 12996 60960
rect 13168 60926 13382 60960
rect 12782 60914 13382 60926
rect 14048 60966 14648 60978
rect 14048 60932 14262 60966
rect 14434 60932 14648 60966
rect 14048 60920 14648 60932
rect 14742 60966 15342 60978
rect 14742 60932 14956 60966
rect 15128 60932 15342 60966
rect 14742 60920 15342 60932
rect 15436 60966 16036 60978
rect 15436 60932 15650 60966
rect 15822 60932 16036 60966
rect 15436 60920 16036 60932
rect 16674 60970 17274 60982
rect 16674 60936 16888 60970
rect 17060 60936 17274 60970
rect 16674 60924 17274 60936
rect 17368 60970 17968 60982
rect 17368 60936 17582 60970
rect 17754 60936 17968 60970
rect 17368 60924 17968 60936
rect 18062 60970 18662 60982
rect 18062 60936 18276 60970
rect 18448 60936 18662 60970
rect 18062 60924 18662 60936
rect 19358 61014 19958 61026
rect 19358 60980 19572 61014
rect 19744 60980 19958 61014
rect 19358 60968 19958 60980
rect 20052 61014 20652 61026
rect 20052 60980 20266 61014
rect 20438 60980 20652 61014
rect 20052 60968 20652 60980
rect 2140 60272 2354 60306
rect 2526 60272 2740 60306
rect 2140 60260 2740 60272
rect 3420 60302 4020 60314
rect 3420 60268 3634 60302
rect 3806 60268 4020 60302
rect 3420 60256 4020 60268
rect 4114 60302 4714 60314
rect 4114 60268 4328 60302
rect 4500 60268 4714 60302
rect 4114 60256 4714 60268
rect 4808 60302 5408 60314
rect 4808 60268 5022 60302
rect 5194 60268 5408 60302
rect 4808 60256 5408 60268
rect 6094 60308 6694 60320
rect 6094 60274 6308 60308
rect 6480 60274 6694 60308
rect 6094 60262 6694 60274
rect 6788 60308 7388 60320
rect 6788 60274 7002 60308
rect 7174 60274 7388 60308
rect 6788 60262 7388 60274
rect 7482 60308 8082 60320
rect 7482 60274 7696 60308
rect 7868 60274 8082 60308
rect 7482 60262 8082 60274
rect 8740 60308 9340 60320
rect 8740 60274 8954 60308
rect 9126 60274 9340 60308
rect 8740 60262 9340 60274
rect 9434 60308 10034 60320
rect 9434 60274 9648 60308
rect 9820 60274 10034 60308
rect 9434 60262 10034 60274
rect 10128 60308 10728 60320
rect 19358 60356 19958 60368
rect 10128 60274 10342 60308
rect 10514 60274 10728 60308
rect 10128 60262 10728 60274
rect 11394 60302 11994 60314
rect 11394 60268 11608 60302
rect 11780 60268 11994 60302
rect 11394 60256 11994 60268
rect 12088 60302 12688 60314
rect 12088 60268 12302 60302
rect 12474 60268 12688 60302
rect 12088 60256 12688 60268
rect 12782 60302 13382 60314
rect 12782 60268 12996 60302
rect 13168 60268 13382 60302
rect 12782 60256 13382 60268
rect 14048 60308 14648 60320
rect 14048 60274 14262 60308
rect 14434 60274 14648 60308
rect 14048 60262 14648 60274
rect 14742 60308 15342 60320
rect 14742 60274 14956 60308
rect 15128 60274 15342 60308
rect 14742 60262 15342 60274
rect 15436 60308 16036 60320
rect 15436 60274 15650 60308
rect 15822 60274 16036 60308
rect 15436 60262 16036 60274
rect 16674 60312 17274 60324
rect 16674 60278 16888 60312
rect 17060 60278 17274 60312
rect 16674 60266 17274 60278
rect 17368 60312 17968 60324
rect 17368 60278 17582 60312
rect 17754 60278 17968 60312
rect 17368 60266 17968 60278
rect 18062 60312 18662 60324
rect 18062 60278 18276 60312
rect 18448 60278 18662 60312
rect 19358 60322 19572 60356
rect 19744 60322 19958 60356
rect 19358 60310 19958 60322
rect 20052 60356 20652 60368
rect 20052 60322 20266 60356
rect 20438 60322 20652 60356
rect 20052 60310 20652 60322
rect 18062 60266 18662 60278
rect 19330 59352 19930 59364
rect 724 59302 1324 59314
rect 724 59268 938 59302
rect 1110 59268 1324 59302
rect 724 59256 1324 59268
rect 1418 59302 2018 59314
rect 1418 59268 1632 59302
rect 1804 59268 2018 59302
rect 1418 59256 2018 59268
rect 2112 59302 2712 59314
rect 2112 59268 2326 59302
rect 2498 59268 2712 59302
rect 2112 59256 2712 59268
rect 3392 59298 3992 59310
rect 3392 59264 3606 59298
rect 3778 59264 3992 59298
rect 3392 59252 3992 59264
rect 4086 59298 4686 59310
rect 4086 59264 4300 59298
rect 4472 59264 4686 59298
rect 4086 59252 4686 59264
rect 4780 59298 5380 59310
rect 4780 59264 4994 59298
rect 5166 59264 5380 59298
rect 4780 59252 5380 59264
rect 6066 59304 6666 59316
rect 6066 59270 6280 59304
rect 6452 59270 6666 59304
rect 6066 59258 6666 59270
rect 6760 59304 7360 59316
rect 6760 59270 6974 59304
rect 7146 59270 7360 59304
rect 6760 59258 7360 59270
rect 7454 59304 8054 59316
rect 7454 59270 7668 59304
rect 7840 59270 8054 59304
rect 7454 59258 8054 59270
rect 8712 59304 9312 59316
rect 8712 59270 8926 59304
rect 9098 59270 9312 59304
rect 8712 59258 9312 59270
rect 9406 59304 10006 59316
rect 9406 59270 9620 59304
rect 9792 59270 10006 59304
rect 9406 59258 10006 59270
rect 10100 59304 10700 59316
rect 10100 59270 10314 59304
rect 10486 59270 10700 59304
rect 10100 59258 10700 59270
rect 11366 59298 11966 59310
rect 11366 59264 11580 59298
rect 11752 59264 11966 59298
rect 724 58644 1324 58656
rect 724 58610 938 58644
rect 1110 58610 1324 58644
rect 724 58598 1324 58610
rect 1418 58644 2018 58656
rect 1418 58610 1632 58644
rect 1804 58610 2018 58644
rect 1418 58598 2018 58610
rect 2112 58644 2712 58656
rect 2112 58610 2326 58644
rect 2498 58610 2712 58644
rect 2112 58598 2712 58610
rect 11366 59252 11966 59264
rect 12060 59298 12660 59310
rect 12060 59264 12274 59298
rect 12446 59264 12660 59298
rect 12060 59252 12660 59264
rect 12754 59298 13354 59310
rect 12754 59264 12968 59298
rect 13140 59264 13354 59298
rect 12754 59252 13354 59264
rect 14020 59304 14620 59316
rect 14020 59270 14234 59304
rect 14406 59270 14620 59304
rect 14020 59258 14620 59270
rect 14714 59304 15314 59316
rect 14714 59270 14928 59304
rect 15100 59270 15314 59304
rect 14714 59258 15314 59270
rect 15408 59304 16008 59316
rect 15408 59270 15622 59304
rect 15794 59270 16008 59304
rect 15408 59258 16008 59270
rect 16646 59308 17246 59320
rect 16646 59274 16860 59308
rect 17032 59274 17246 59308
rect 16646 59262 17246 59274
rect 17340 59308 17940 59320
rect 17340 59274 17554 59308
rect 17726 59274 17940 59308
rect 17340 59262 17940 59274
rect 18034 59308 18634 59320
rect 18034 59274 18248 59308
rect 18420 59274 18634 59308
rect 19330 59318 19544 59352
rect 19716 59318 19930 59352
rect 19330 59306 19930 59318
rect 20024 59352 20624 59364
rect 20024 59318 20238 59352
rect 20410 59318 20624 59352
rect 20024 59306 20624 59318
rect 18034 59262 18634 59274
rect 3392 58640 3992 58652
rect 3392 58606 3606 58640
rect 3778 58606 3992 58640
rect 3392 58594 3992 58606
rect 4086 58640 4686 58652
rect 4086 58606 4300 58640
rect 4472 58606 4686 58640
rect 4086 58594 4686 58606
rect 4780 58640 5380 58652
rect 4780 58606 4994 58640
rect 5166 58606 5380 58640
rect 4780 58594 5380 58606
rect 6066 58646 6666 58658
rect 6066 58612 6280 58646
rect 6452 58612 6666 58646
rect 6066 58600 6666 58612
rect 6760 58646 7360 58658
rect 6760 58612 6974 58646
rect 7146 58612 7360 58646
rect 6760 58600 7360 58612
rect 7454 58646 8054 58658
rect 7454 58612 7668 58646
rect 7840 58612 8054 58646
rect 7454 58600 8054 58612
rect 8712 58646 9312 58658
rect 8712 58612 8926 58646
rect 9098 58612 9312 58646
rect 8712 58600 9312 58612
rect 9406 58646 10006 58658
rect 9406 58612 9620 58646
rect 9792 58612 10006 58646
rect 9406 58600 10006 58612
rect 10100 58646 10700 58658
rect 10100 58612 10314 58646
rect 10486 58612 10700 58646
rect 10100 58600 10700 58612
rect 724 57986 1324 57998
rect 724 57952 938 57986
rect 1110 57952 1324 57986
rect 724 57940 1324 57952
rect 1418 57986 2018 57998
rect 1418 57952 1632 57986
rect 1804 57952 2018 57986
rect 1418 57940 2018 57952
rect 2112 57986 2712 57998
rect 2112 57952 2326 57986
rect 2498 57952 2712 57986
rect 2112 57940 2712 57952
rect 11366 58640 11966 58652
rect 11366 58606 11580 58640
rect 11752 58606 11966 58640
rect 11366 58594 11966 58606
rect 12060 58640 12660 58652
rect 12060 58606 12274 58640
rect 12446 58606 12660 58640
rect 12060 58594 12660 58606
rect 12754 58640 13354 58652
rect 12754 58606 12968 58640
rect 13140 58606 13354 58640
rect 12754 58594 13354 58606
rect 14020 58646 14620 58658
rect 14020 58612 14234 58646
rect 14406 58612 14620 58646
rect 14020 58600 14620 58612
rect 14714 58646 15314 58658
rect 14714 58612 14928 58646
rect 15100 58612 15314 58646
rect 14714 58600 15314 58612
rect 15408 58646 16008 58658
rect 15408 58612 15622 58646
rect 15794 58612 16008 58646
rect 15408 58600 16008 58612
rect 16646 58650 17246 58662
rect 16646 58616 16860 58650
rect 17032 58616 17246 58650
rect 16646 58604 17246 58616
rect 17340 58650 17940 58662
rect 17340 58616 17554 58650
rect 17726 58616 17940 58650
rect 17340 58604 17940 58616
rect 18034 58650 18634 58662
rect 18034 58616 18248 58650
rect 18420 58616 18634 58650
rect 18034 58604 18634 58616
rect 19330 58694 19930 58706
rect 19330 58660 19544 58694
rect 19716 58660 19930 58694
rect 19330 58648 19930 58660
rect 20024 58694 20624 58706
rect 20024 58660 20238 58694
rect 20410 58660 20624 58694
rect 20024 58648 20624 58660
rect 3392 57982 3992 57994
rect 3392 57948 3606 57982
rect 3778 57948 3992 57982
rect 3392 57936 3992 57948
rect 4086 57982 4686 57994
rect 4086 57948 4300 57982
rect 4472 57948 4686 57982
rect 4086 57936 4686 57948
rect 4780 57982 5380 57994
rect 4780 57948 4994 57982
rect 5166 57948 5380 57982
rect 4780 57936 5380 57948
rect 6066 57988 6666 58000
rect 6066 57954 6280 57988
rect 6452 57954 6666 57988
rect 6066 57942 6666 57954
rect 6760 57988 7360 58000
rect 6760 57954 6974 57988
rect 7146 57954 7360 57988
rect 6760 57942 7360 57954
rect 7454 57988 8054 58000
rect 7454 57954 7668 57988
rect 7840 57954 8054 57988
rect 7454 57942 8054 57954
rect 8712 57988 9312 58000
rect 8712 57954 8926 57988
rect 9098 57954 9312 57988
rect 8712 57942 9312 57954
rect 9406 57988 10006 58000
rect 9406 57954 9620 57988
rect 9792 57954 10006 57988
rect 9406 57942 10006 57954
rect 10100 57988 10700 58000
rect 10100 57954 10314 57988
rect 10486 57954 10700 57988
rect 10100 57942 10700 57954
rect 724 57328 1324 57340
rect 724 57294 938 57328
rect 1110 57294 1324 57328
rect 724 57282 1324 57294
rect 1418 57328 2018 57340
rect 1418 57294 1632 57328
rect 1804 57294 2018 57328
rect 1418 57282 2018 57294
rect 2112 57328 2712 57340
rect 2112 57294 2326 57328
rect 2498 57294 2712 57328
rect 2112 57282 2712 57294
rect 11366 57982 11966 57994
rect 11366 57948 11580 57982
rect 11752 57948 11966 57982
rect 11366 57936 11966 57948
rect 12060 57982 12660 57994
rect 12060 57948 12274 57982
rect 12446 57948 12660 57982
rect 12060 57936 12660 57948
rect 12754 57982 13354 57994
rect 12754 57948 12968 57982
rect 13140 57948 13354 57982
rect 12754 57936 13354 57948
rect 14020 57988 14620 58000
rect 14020 57954 14234 57988
rect 14406 57954 14620 57988
rect 14020 57942 14620 57954
rect 14714 57988 15314 58000
rect 14714 57954 14928 57988
rect 15100 57954 15314 57988
rect 14714 57942 15314 57954
rect 15408 57988 16008 58000
rect 15408 57954 15622 57988
rect 15794 57954 16008 57988
rect 15408 57942 16008 57954
rect 16646 57992 17246 58004
rect 16646 57958 16860 57992
rect 17032 57958 17246 57992
rect 16646 57946 17246 57958
rect 17340 57992 17940 58004
rect 17340 57958 17554 57992
rect 17726 57958 17940 57992
rect 17340 57946 17940 57958
rect 18034 57992 18634 58004
rect 18034 57958 18248 57992
rect 18420 57958 18634 57992
rect 18034 57946 18634 57958
rect 19330 58036 19930 58048
rect 19330 58002 19544 58036
rect 19716 58002 19930 58036
rect 19330 57990 19930 58002
rect 20024 58036 20624 58048
rect 20024 58002 20238 58036
rect 20410 58002 20624 58036
rect 20024 57990 20624 58002
rect 3392 57324 3992 57336
rect 3392 57290 3606 57324
rect 3778 57290 3992 57324
rect 3392 57278 3992 57290
rect 4086 57324 4686 57336
rect 4086 57290 4300 57324
rect 4472 57290 4686 57324
rect 4086 57278 4686 57290
rect 4780 57324 5380 57336
rect 4780 57290 4994 57324
rect 5166 57290 5380 57324
rect 4780 57278 5380 57290
rect 6066 57330 6666 57342
rect 6066 57296 6280 57330
rect 6452 57296 6666 57330
rect 6066 57284 6666 57296
rect 6760 57330 7360 57342
rect 6760 57296 6974 57330
rect 7146 57296 7360 57330
rect 6760 57284 7360 57296
rect 7454 57330 8054 57342
rect 7454 57296 7668 57330
rect 7840 57296 8054 57330
rect 7454 57284 8054 57296
rect 8712 57330 9312 57342
rect 8712 57296 8926 57330
rect 9098 57296 9312 57330
rect 8712 57284 9312 57296
rect 9406 57330 10006 57342
rect 9406 57296 9620 57330
rect 9792 57296 10006 57330
rect 9406 57284 10006 57296
rect 10100 57330 10700 57342
rect 10100 57296 10314 57330
rect 10486 57296 10700 57330
rect 10100 57284 10700 57296
rect 724 56670 1324 56682
rect 724 56636 938 56670
rect 1110 56636 1324 56670
rect 724 56624 1324 56636
rect 1418 56670 2018 56682
rect 1418 56636 1632 56670
rect 1804 56636 2018 56670
rect 1418 56624 2018 56636
rect 2112 56670 2712 56682
rect 2112 56636 2326 56670
rect 2498 56636 2712 56670
rect 2112 56624 2712 56636
rect 11366 57324 11966 57336
rect 11366 57290 11580 57324
rect 11752 57290 11966 57324
rect 11366 57278 11966 57290
rect 12060 57324 12660 57336
rect 12060 57290 12274 57324
rect 12446 57290 12660 57324
rect 12060 57278 12660 57290
rect 12754 57324 13354 57336
rect 12754 57290 12968 57324
rect 13140 57290 13354 57324
rect 12754 57278 13354 57290
rect 14020 57330 14620 57342
rect 14020 57296 14234 57330
rect 14406 57296 14620 57330
rect 14020 57284 14620 57296
rect 14714 57330 15314 57342
rect 14714 57296 14928 57330
rect 15100 57296 15314 57330
rect 14714 57284 15314 57296
rect 15408 57330 16008 57342
rect 15408 57296 15622 57330
rect 15794 57296 16008 57330
rect 15408 57284 16008 57296
rect 16646 57334 17246 57346
rect 16646 57300 16860 57334
rect 17032 57300 17246 57334
rect 16646 57288 17246 57300
rect 17340 57334 17940 57346
rect 17340 57300 17554 57334
rect 17726 57300 17940 57334
rect 17340 57288 17940 57300
rect 18034 57334 18634 57346
rect 18034 57300 18248 57334
rect 18420 57300 18634 57334
rect 18034 57288 18634 57300
rect 19330 57378 19930 57390
rect 19330 57344 19544 57378
rect 19716 57344 19930 57378
rect 19330 57332 19930 57344
rect 20024 57378 20624 57390
rect 20024 57344 20238 57378
rect 20410 57344 20624 57378
rect 20024 57332 20624 57344
rect 3392 56666 3992 56678
rect 3392 56632 3606 56666
rect 3778 56632 3992 56666
rect 3392 56620 3992 56632
rect 4086 56666 4686 56678
rect 4086 56632 4300 56666
rect 4472 56632 4686 56666
rect 4086 56620 4686 56632
rect 4780 56666 5380 56678
rect 4780 56632 4994 56666
rect 5166 56632 5380 56666
rect 4780 56620 5380 56632
rect 6066 56672 6666 56684
rect 6066 56638 6280 56672
rect 6452 56638 6666 56672
rect 6066 56626 6666 56638
rect 6760 56672 7360 56684
rect 6760 56638 6974 56672
rect 7146 56638 7360 56672
rect 6760 56626 7360 56638
rect 7454 56672 8054 56684
rect 7454 56638 7668 56672
rect 7840 56638 8054 56672
rect 7454 56626 8054 56638
rect 8712 56672 9312 56684
rect 8712 56638 8926 56672
rect 9098 56638 9312 56672
rect 8712 56626 9312 56638
rect 9406 56672 10006 56684
rect 9406 56638 9620 56672
rect 9792 56638 10006 56672
rect 9406 56626 10006 56638
rect 10100 56672 10700 56684
rect 10100 56638 10314 56672
rect 10486 56638 10700 56672
rect 10100 56626 10700 56638
rect 724 56012 1324 56024
rect 724 55978 938 56012
rect 1110 55978 1324 56012
rect 724 55966 1324 55978
rect 1418 56012 2018 56024
rect 1418 55978 1632 56012
rect 1804 55978 2018 56012
rect 1418 55966 2018 55978
rect 2112 56012 2712 56024
rect 2112 55978 2326 56012
rect 2498 55978 2712 56012
rect 2112 55966 2712 55978
rect 11366 56666 11966 56678
rect 11366 56632 11580 56666
rect 11752 56632 11966 56666
rect 11366 56620 11966 56632
rect 12060 56666 12660 56678
rect 12060 56632 12274 56666
rect 12446 56632 12660 56666
rect 12060 56620 12660 56632
rect 12754 56666 13354 56678
rect 12754 56632 12968 56666
rect 13140 56632 13354 56666
rect 12754 56620 13354 56632
rect 14020 56672 14620 56684
rect 14020 56638 14234 56672
rect 14406 56638 14620 56672
rect 14020 56626 14620 56638
rect 14714 56672 15314 56684
rect 14714 56638 14928 56672
rect 15100 56638 15314 56672
rect 14714 56626 15314 56638
rect 15408 56672 16008 56684
rect 15408 56638 15622 56672
rect 15794 56638 16008 56672
rect 15408 56626 16008 56638
rect 16646 56676 17246 56688
rect 16646 56642 16860 56676
rect 17032 56642 17246 56676
rect 16646 56630 17246 56642
rect 17340 56676 17940 56688
rect 17340 56642 17554 56676
rect 17726 56642 17940 56676
rect 17340 56630 17940 56642
rect 18034 56676 18634 56688
rect 18034 56642 18248 56676
rect 18420 56642 18634 56676
rect 18034 56630 18634 56642
rect 19330 56720 19930 56732
rect 19330 56686 19544 56720
rect 19716 56686 19930 56720
rect 19330 56674 19930 56686
rect 20024 56720 20624 56732
rect 20024 56686 20238 56720
rect 20410 56686 20624 56720
rect 20024 56674 20624 56686
rect 3392 56008 3992 56020
rect 3392 55974 3606 56008
rect 3778 55974 3992 56008
rect 3392 55962 3992 55974
rect 4086 56008 4686 56020
rect 4086 55974 4300 56008
rect 4472 55974 4686 56008
rect 4086 55962 4686 55974
rect 4780 56008 5380 56020
rect 4780 55974 4994 56008
rect 5166 55974 5380 56008
rect 4780 55962 5380 55974
rect 6066 56014 6666 56026
rect 6066 55980 6280 56014
rect 6452 55980 6666 56014
rect 6066 55968 6666 55980
rect 6760 56014 7360 56026
rect 6760 55980 6974 56014
rect 7146 55980 7360 56014
rect 6760 55968 7360 55980
rect 7454 56014 8054 56026
rect 7454 55980 7668 56014
rect 7840 55980 8054 56014
rect 7454 55968 8054 55980
rect 8712 56014 9312 56026
rect 8712 55980 8926 56014
rect 9098 55980 9312 56014
rect 8712 55968 9312 55980
rect 9406 56014 10006 56026
rect 9406 55980 9620 56014
rect 9792 55980 10006 56014
rect 9406 55968 10006 55980
rect 10100 56014 10700 56026
rect 10100 55980 10314 56014
rect 10486 55980 10700 56014
rect 10100 55968 10700 55980
rect 724 55354 1324 55366
rect 724 55320 938 55354
rect 1110 55320 1324 55354
rect 724 55308 1324 55320
rect 1418 55354 2018 55366
rect 1418 55320 1632 55354
rect 1804 55320 2018 55354
rect 1418 55308 2018 55320
rect 2112 55354 2712 55366
rect 2112 55320 2326 55354
rect 2498 55320 2712 55354
rect 2112 55308 2712 55320
rect 11366 56008 11966 56020
rect 11366 55974 11580 56008
rect 11752 55974 11966 56008
rect 11366 55962 11966 55974
rect 12060 56008 12660 56020
rect 12060 55974 12274 56008
rect 12446 55974 12660 56008
rect 12060 55962 12660 55974
rect 12754 56008 13354 56020
rect 12754 55974 12968 56008
rect 13140 55974 13354 56008
rect 12754 55962 13354 55974
rect 14020 56014 14620 56026
rect 14020 55980 14234 56014
rect 14406 55980 14620 56014
rect 14020 55968 14620 55980
rect 14714 56014 15314 56026
rect 14714 55980 14928 56014
rect 15100 55980 15314 56014
rect 14714 55968 15314 55980
rect 15408 56014 16008 56026
rect 15408 55980 15622 56014
rect 15794 55980 16008 56014
rect 15408 55968 16008 55980
rect 16646 56018 17246 56030
rect 16646 55984 16860 56018
rect 17032 55984 17246 56018
rect 16646 55972 17246 55984
rect 17340 56018 17940 56030
rect 17340 55984 17554 56018
rect 17726 55984 17940 56018
rect 17340 55972 17940 55984
rect 18034 56018 18634 56030
rect 18034 55984 18248 56018
rect 18420 55984 18634 56018
rect 18034 55972 18634 55984
rect 19330 56062 19930 56074
rect 19330 56028 19544 56062
rect 19716 56028 19930 56062
rect 19330 56016 19930 56028
rect 20024 56062 20624 56074
rect 20024 56028 20238 56062
rect 20410 56028 20624 56062
rect 20024 56016 20624 56028
rect 3392 55350 3992 55362
rect 3392 55316 3606 55350
rect 3778 55316 3992 55350
rect 3392 55304 3992 55316
rect 4086 55350 4686 55362
rect 4086 55316 4300 55350
rect 4472 55316 4686 55350
rect 4086 55304 4686 55316
rect 4780 55350 5380 55362
rect 4780 55316 4994 55350
rect 5166 55316 5380 55350
rect 4780 55304 5380 55316
rect 6066 55356 6666 55368
rect 6066 55322 6280 55356
rect 6452 55322 6666 55356
rect 6066 55310 6666 55322
rect 6760 55356 7360 55368
rect 6760 55322 6974 55356
rect 7146 55322 7360 55356
rect 6760 55310 7360 55322
rect 7454 55356 8054 55368
rect 7454 55322 7668 55356
rect 7840 55322 8054 55356
rect 7454 55310 8054 55322
rect 8712 55356 9312 55368
rect 8712 55322 8926 55356
rect 9098 55322 9312 55356
rect 8712 55310 9312 55322
rect 9406 55356 10006 55368
rect 9406 55322 9620 55356
rect 9792 55322 10006 55356
rect 9406 55310 10006 55322
rect 10100 55356 10700 55368
rect 10100 55322 10314 55356
rect 10486 55322 10700 55356
rect 10100 55310 10700 55322
rect 724 54696 1324 54708
rect 724 54662 938 54696
rect 1110 54662 1324 54696
rect 724 54650 1324 54662
rect 1418 54696 2018 54708
rect 1418 54662 1632 54696
rect 1804 54662 2018 54696
rect 1418 54650 2018 54662
rect 2112 54696 2712 54708
rect 2112 54662 2326 54696
rect 2498 54662 2712 54696
rect 2112 54650 2712 54662
rect 11366 55350 11966 55362
rect 11366 55316 11580 55350
rect 11752 55316 11966 55350
rect 11366 55304 11966 55316
rect 12060 55350 12660 55362
rect 12060 55316 12274 55350
rect 12446 55316 12660 55350
rect 12060 55304 12660 55316
rect 12754 55350 13354 55362
rect 12754 55316 12968 55350
rect 13140 55316 13354 55350
rect 12754 55304 13354 55316
rect 14020 55356 14620 55368
rect 14020 55322 14234 55356
rect 14406 55322 14620 55356
rect 14020 55310 14620 55322
rect 14714 55356 15314 55368
rect 14714 55322 14928 55356
rect 15100 55322 15314 55356
rect 14714 55310 15314 55322
rect 15408 55356 16008 55368
rect 15408 55322 15622 55356
rect 15794 55322 16008 55356
rect 15408 55310 16008 55322
rect 16646 55360 17246 55372
rect 16646 55326 16860 55360
rect 17032 55326 17246 55360
rect 16646 55314 17246 55326
rect 17340 55360 17940 55372
rect 17340 55326 17554 55360
rect 17726 55326 17940 55360
rect 17340 55314 17940 55326
rect 18034 55360 18634 55372
rect 18034 55326 18248 55360
rect 18420 55326 18634 55360
rect 18034 55314 18634 55326
rect 19330 55404 19930 55416
rect 19330 55370 19544 55404
rect 19716 55370 19930 55404
rect 19330 55358 19930 55370
rect 20024 55404 20624 55416
rect 20024 55370 20238 55404
rect 20410 55370 20624 55404
rect 20024 55358 20624 55370
rect 3392 54692 3992 54704
rect 3392 54658 3606 54692
rect 3778 54658 3992 54692
rect 3392 54646 3992 54658
rect 4086 54692 4686 54704
rect 4086 54658 4300 54692
rect 4472 54658 4686 54692
rect 4086 54646 4686 54658
rect 4780 54692 5380 54704
rect 4780 54658 4994 54692
rect 5166 54658 5380 54692
rect 4780 54646 5380 54658
rect 6066 54698 6666 54710
rect 6066 54664 6280 54698
rect 6452 54664 6666 54698
rect 6066 54652 6666 54664
rect 6760 54698 7360 54710
rect 6760 54664 6974 54698
rect 7146 54664 7360 54698
rect 6760 54652 7360 54664
rect 7454 54698 8054 54710
rect 7454 54664 7668 54698
rect 7840 54664 8054 54698
rect 7454 54652 8054 54664
rect 8712 54698 9312 54710
rect 8712 54664 8926 54698
rect 9098 54664 9312 54698
rect 8712 54652 9312 54664
rect 9406 54698 10006 54710
rect 9406 54664 9620 54698
rect 9792 54664 10006 54698
rect 9406 54652 10006 54664
rect 10100 54698 10700 54710
rect 10100 54664 10314 54698
rect 10486 54664 10700 54698
rect 10100 54652 10700 54664
rect 724 54038 1324 54050
rect 724 54004 938 54038
rect 1110 54004 1324 54038
rect 724 53992 1324 54004
rect 1418 54038 2018 54050
rect 1418 54004 1632 54038
rect 1804 54004 2018 54038
rect 1418 53992 2018 54004
rect 2112 54038 2712 54050
rect 11366 54692 11966 54704
rect 11366 54658 11580 54692
rect 11752 54658 11966 54692
rect 11366 54646 11966 54658
rect 12060 54692 12660 54704
rect 12060 54658 12274 54692
rect 12446 54658 12660 54692
rect 12060 54646 12660 54658
rect 12754 54692 13354 54704
rect 12754 54658 12968 54692
rect 13140 54658 13354 54692
rect 12754 54646 13354 54658
rect 14020 54698 14620 54710
rect 14020 54664 14234 54698
rect 14406 54664 14620 54698
rect 14020 54652 14620 54664
rect 14714 54698 15314 54710
rect 14714 54664 14928 54698
rect 15100 54664 15314 54698
rect 14714 54652 15314 54664
rect 15408 54698 16008 54710
rect 15408 54664 15622 54698
rect 15794 54664 16008 54698
rect 15408 54652 16008 54664
rect 16646 54702 17246 54714
rect 16646 54668 16860 54702
rect 17032 54668 17246 54702
rect 16646 54656 17246 54668
rect 17340 54702 17940 54714
rect 17340 54668 17554 54702
rect 17726 54668 17940 54702
rect 17340 54656 17940 54668
rect 18034 54702 18634 54714
rect 18034 54668 18248 54702
rect 18420 54668 18634 54702
rect 18034 54656 18634 54668
rect 19330 54746 19930 54758
rect 19330 54712 19544 54746
rect 19716 54712 19930 54746
rect 19330 54700 19930 54712
rect 20024 54746 20624 54758
rect 20024 54712 20238 54746
rect 20410 54712 20624 54746
rect 20024 54700 20624 54712
rect 2112 54004 2326 54038
rect 2498 54004 2712 54038
rect 2112 53992 2712 54004
rect 3392 54034 3992 54046
rect 3392 54000 3606 54034
rect 3778 54000 3992 54034
rect 3392 53988 3992 54000
rect 4086 54034 4686 54046
rect 4086 54000 4300 54034
rect 4472 54000 4686 54034
rect 4086 53988 4686 54000
rect 4780 54034 5380 54046
rect 4780 54000 4994 54034
rect 5166 54000 5380 54034
rect 4780 53988 5380 54000
rect 6066 54040 6666 54052
rect 6066 54006 6280 54040
rect 6452 54006 6666 54040
rect 6066 53994 6666 54006
rect 6760 54040 7360 54052
rect 6760 54006 6974 54040
rect 7146 54006 7360 54040
rect 6760 53994 7360 54006
rect 7454 54040 8054 54052
rect 7454 54006 7668 54040
rect 7840 54006 8054 54040
rect 7454 53994 8054 54006
rect 8712 54040 9312 54052
rect 8712 54006 8926 54040
rect 9098 54006 9312 54040
rect 8712 53994 9312 54006
rect 9406 54040 10006 54052
rect 9406 54006 9620 54040
rect 9792 54006 10006 54040
rect 9406 53994 10006 54006
rect 10100 54040 10700 54052
rect 19330 54088 19930 54100
rect 10100 54006 10314 54040
rect 10486 54006 10700 54040
rect 10100 53994 10700 54006
rect 11366 54034 11966 54046
rect 11366 54000 11580 54034
rect 11752 54000 11966 54034
rect 11366 53988 11966 54000
rect 12060 54034 12660 54046
rect 12060 54000 12274 54034
rect 12446 54000 12660 54034
rect 12060 53988 12660 54000
rect 12754 54034 13354 54046
rect 12754 54000 12968 54034
rect 13140 54000 13354 54034
rect 12754 53988 13354 54000
rect 14020 54040 14620 54052
rect 14020 54006 14234 54040
rect 14406 54006 14620 54040
rect 14020 53994 14620 54006
rect 14714 54040 15314 54052
rect 14714 54006 14928 54040
rect 15100 54006 15314 54040
rect 14714 53994 15314 54006
rect 15408 54040 16008 54052
rect 15408 54006 15622 54040
rect 15794 54006 16008 54040
rect 15408 53994 16008 54006
rect 16646 54044 17246 54056
rect 16646 54010 16860 54044
rect 17032 54010 17246 54044
rect 16646 53998 17246 54010
rect 17340 54044 17940 54056
rect 17340 54010 17554 54044
rect 17726 54010 17940 54044
rect 17340 53998 17940 54010
rect 18034 54044 18634 54056
rect 18034 54010 18248 54044
rect 18420 54010 18634 54044
rect 19330 54054 19544 54088
rect 19716 54054 19930 54088
rect 19330 54042 19930 54054
rect 20024 54088 20624 54100
rect 20024 54054 20238 54088
rect 20410 54054 20624 54088
rect 20024 54042 20624 54054
rect 18034 53998 18634 54010
rect 19330 52986 19930 52998
rect 724 52936 1324 52948
rect 724 52902 938 52936
rect 1110 52902 1324 52936
rect 724 52890 1324 52902
rect 1418 52936 2018 52948
rect 1418 52902 1632 52936
rect 1804 52902 2018 52936
rect 1418 52890 2018 52902
rect 2112 52936 2712 52948
rect 2112 52902 2326 52936
rect 2498 52902 2712 52936
rect 2112 52890 2712 52902
rect 3392 52932 3992 52944
rect 3392 52898 3606 52932
rect 3778 52898 3992 52932
rect 3392 52886 3992 52898
rect 4086 52932 4686 52944
rect 4086 52898 4300 52932
rect 4472 52898 4686 52932
rect 4086 52886 4686 52898
rect 4780 52932 5380 52944
rect 4780 52898 4994 52932
rect 5166 52898 5380 52932
rect 4780 52886 5380 52898
rect 6066 52938 6666 52950
rect 6066 52904 6280 52938
rect 6452 52904 6666 52938
rect 6066 52892 6666 52904
rect 6760 52938 7360 52950
rect 6760 52904 6974 52938
rect 7146 52904 7360 52938
rect 6760 52892 7360 52904
rect 7454 52938 8054 52950
rect 7454 52904 7668 52938
rect 7840 52904 8054 52938
rect 7454 52892 8054 52904
rect 8712 52938 9312 52950
rect 8712 52904 8926 52938
rect 9098 52904 9312 52938
rect 8712 52892 9312 52904
rect 9406 52938 10006 52950
rect 9406 52904 9620 52938
rect 9792 52904 10006 52938
rect 9406 52892 10006 52904
rect 10100 52938 10700 52950
rect 10100 52904 10314 52938
rect 10486 52904 10700 52938
rect 10100 52892 10700 52904
rect 11366 52932 11966 52944
rect 11366 52898 11580 52932
rect 11752 52898 11966 52932
rect 724 52278 1324 52290
rect 724 52244 938 52278
rect 1110 52244 1324 52278
rect 724 52232 1324 52244
rect 1418 52278 2018 52290
rect 1418 52244 1632 52278
rect 1804 52244 2018 52278
rect 1418 52232 2018 52244
rect 2112 52278 2712 52290
rect 2112 52244 2326 52278
rect 2498 52244 2712 52278
rect 2112 52232 2712 52244
rect 11366 52886 11966 52898
rect 12060 52932 12660 52944
rect 12060 52898 12274 52932
rect 12446 52898 12660 52932
rect 12060 52886 12660 52898
rect 12754 52932 13354 52944
rect 12754 52898 12968 52932
rect 13140 52898 13354 52932
rect 12754 52886 13354 52898
rect 14020 52938 14620 52950
rect 14020 52904 14234 52938
rect 14406 52904 14620 52938
rect 14020 52892 14620 52904
rect 14714 52938 15314 52950
rect 14714 52904 14928 52938
rect 15100 52904 15314 52938
rect 14714 52892 15314 52904
rect 15408 52938 16008 52950
rect 15408 52904 15622 52938
rect 15794 52904 16008 52938
rect 15408 52892 16008 52904
rect 16646 52942 17246 52954
rect 16646 52908 16860 52942
rect 17032 52908 17246 52942
rect 16646 52896 17246 52908
rect 17340 52942 17940 52954
rect 17340 52908 17554 52942
rect 17726 52908 17940 52942
rect 17340 52896 17940 52908
rect 18034 52942 18634 52954
rect 18034 52908 18248 52942
rect 18420 52908 18634 52942
rect 19330 52952 19544 52986
rect 19716 52952 19930 52986
rect 19330 52940 19930 52952
rect 20024 52986 20624 52998
rect 20024 52952 20238 52986
rect 20410 52952 20624 52986
rect 20024 52940 20624 52952
rect 18034 52896 18634 52908
rect 3392 52274 3992 52286
rect 3392 52240 3606 52274
rect 3778 52240 3992 52274
rect 3392 52228 3992 52240
rect 4086 52274 4686 52286
rect 4086 52240 4300 52274
rect 4472 52240 4686 52274
rect 4086 52228 4686 52240
rect 4780 52274 5380 52286
rect 4780 52240 4994 52274
rect 5166 52240 5380 52274
rect 4780 52228 5380 52240
rect 6066 52280 6666 52292
rect 6066 52246 6280 52280
rect 6452 52246 6666 52280
rect 6066 52234 6666 52246
rect 6760 52280 7360 52292
rect 6760 52246 6974 52280
rect 7146 52246 7360 52280
rect 6760 52234 7360 52246
rect 7454 52280 8054 52292
rect 7454 52246 7668 52280
rect 7840 52246 8054 52280
rect 7454 52234 8054 52246
rect 8712 52280 9312 52292
rect 8712 52246 8926 52280
rect 9098 52246 9312 52280
rect 8712 52234 9312 52246
rect 9406 52280 10006 52292
rect 9406 52246 9620 52280
rect 9792 52246 10006 52280
rect 9406 52234 10006 52246
rect 10100 52280 10700 52292
rect 10100 52246 10314 52280
rect 10486 52246 10700 52280
rect 10100 52234 10700 52246
rect 724 51620 1324 51632
rect 724 51586 938 51620
rect 1110 51586 1324 51620
rect 724 51574 1324 51586
rect 1418 51620 2018 51632
rect 1418 51586 1632 51620
rect 1804 51586 2018 51620
rect 1418 51574 2018 51586
rect 2112 51620 2712 51632
rect 2112 51586 2326 51620
rect 2498 51586 2712 51620
rect 2112 51574 2712 51586
rect 11366 52274 11966 52286
rect 11366 52240 11580 52274
rect 11752 52240 11966 52274
rect 11366 52228 11966 52240
rect 12060 52274 12660 52286
rect 12060 52240 12274 52274
rect 12446 52240 12660 52274
rect 12060 52228 12660 52240
rect 12754 52274 13354 52286
rect 12754 52240 12968 52274
rect 13140 52240 13354 52274
rect 12754 52228 13354 52240
rect 14020 52280 14620 52292
rect 14020 52246 14234 52280
rect 14406 52246 14620 52280
rect 14020 52234 14620 52246
rect 14714 52280 15314 52292
rect 14714 52246 14928 52280
rect 15100 52246 15314 52280
rect 14714 52234 15314 52246
rect 15408 52280 16008 52292
rect 15408 52246 15622 52280
rect 15794 52246 16008 52280
rect 15408 52234 16008 52246
rect 16646 52284 17246 52296
rect 16646 52250 16860 52284
rect 17032 52250 17246 52284
rect 16646 52238 17246 52250
rect 17340 52284 17940 52296
rect 17340 52250 17554 52284
rect 17726 52250 17940 52284
rect 17340 52238 17940 52250
rect 18034 52284 18634 52296
rect 18034 52250 18248 52284
rect 18420 52250 18634 52284
rect 18034 52238 18634 52250
rect 19330 52328 19930 52340
rect 19330 52294 19544 52328
rect 19716 52294 19930 52328
rect 19330 52282 19930 52294
rect 20024 52328 20624 52340
rect 20024 52294 20238 52328
rect 20410 52294 20624 52328
rect 20024 52282 20624 52294
rect 3392 51616 3992 51628
rect 3392 51582 3606 51616
rect 3778 51582 3992 51616
rect 3392 51570 3992 51582
rect 4086 51616 4686 51628
rect 4086 51582 4300 51616
rect 4472 51582 4686 51616
rect 4086 51570 4686 51582
rect 4780 51616 5380 51628
rect 4780 51582 4994 51616
rect 5166 51582 5380 51616
rect 4780 51570 5380 51582
rect 6066 51622 6666 51634
rect 6066 51588 6280 51622
rect 6452 51588 6666 51622
rect 6066 51576 6666 51588
rect 6760 51622 7360 51634
rect 6760 51588 6974 51622
rect 7146 51588 7360 51622
rect 6760 51576 7360 51588
rect 7454 51622 8054 51634
rect 7454 51588 7668 51622
rect 7840 51588 8054 51622
rect 7454 51576 8054 51588
rect 8712 51622 9312 51634
rect 8712 51588 8926 51622
rect 9098 51588 9312 51622
rect 8712 51576 9312 51588
rect 9406 51622 10006 51634
rect 9406 51588 9620 51622
rect 9792 51588 10006 51622
rect 9406 51576 10006 51588
rect 10100 51622 10700 51634
rect 10100 51588 10314 51622
rect 10486 51588 10700 51622
rect 10100 51576 10700 51588
rect 724 50962 1324 50974
rect 724 50928 938 50962
rect 1110 50928 1324 50962
rect 724 50916 1324 50928
rect 1418 50962 2018 50974
rect 1418 50928 1632 50962
rect 1804 50928 2018 50962
rect 1418 50916 2018 50928
rect 2112 50962 2712 50974
rect 2112 50928 2326 50962
rect 2498 50928 2712 50962
rect 2112 50916 2712 50928
rect 11366 51616 11966 51628
rect 11366 51582 11580 51616
rect 11752 51582 11966 51616
rect 11366 51570 11966 51582
rect 12060 51616 12660 51628
rect 12060 51582 12274 51616
rect 12446 51582 12660 51616
rect 12060 51570 12660 51582
rect 12754 51616 13354 51628
rect 12754 51582 12968 51616
rect 13140 51582 13354 51616
rect 12754 51570 13354 51582
rect 14020 51622 14620 51634
rect 14020 51588 14234 51622
rect 14406 51588 14620 51622
rect 14020 51576 14620 51588
rect 14714 51622 15314 51634
rect 14714 51588 14928 51622
rect 15100 51588 15314 51622
rect 14714 51576 15314 51588
rect 15408 51622 16008 51634
rect 15408 51588 15622 51622
rect 15794 51588 16008 51622
rect 15408 51576 16008 51588
rect 16646 51626 17246 51638
rect 16646 51592 16860 51626
rect 17032 51592 17246 51626
rect 16646 51580 17246 51592
rect 17340 51626 17940 51638
rect 17340 51592 17554 51626
rect 17726 51592 17940 51626
rect 17340 51580 17940 51592
rect 18034 51626 18634 51638
rect 18034 51592 18248 51626
rect 18420 51592 18634 51626
rect 18034 51580 18634 51592
rect 19330 51670 19930 51682
rect 19330 51636 19544 51670
rect 19716 51636 19930 51670
rect 19330 51624 19930 51636
rect 20024 51670 20624 51682
rect 20024 51636 20238 51670
rect 20410 51636 20624 51670
rect 20024 51624 20624 51636
rect 3392 50958 3992 50970
rect 3392 50924 3606 50958
rect 3778 50924 3992 50958
rect 3392 50912 3992 50924
rect 4086 50958 4686 50970
rect 4086 50924 4300 50958
rect 4472 50924 4686 50958
rect 4086 50912 4686 50924
rect 4780 50958 5380 50970
rect 4780 50924 4994 50958
rect 5166 50924 5380 50958
rect 4780 50912 5380 50924
rect 6066 50964 6666 50976
rect 6066 50930 6280 50964
rect 6452 50930 6666 50964
rect 6066 50918 6666 50930
rect 6760 50964 7360 50976
rect 6760 50930 6974 50964
rect 7146 50930 7360 50964
rect 6760 50918 7360 50930
rect 7454 50964 8054 50976
rect 7454 50930 7668 50964
rect 7840 50930 8054 50964
rect 7454 50918 8054 50930
rect 8712 50964 9312 50976
rect 8712 50930 8926 50964
rect 9098 50930 9312 50964
rect 8712 50918 9312 50930
rect 9406 50964 10006 50976
rect 9406 50930 9620 50964
rect 9792 50930 10006 50964
rect 9406 50918 10006 50930
rect 10100 50964 10700 50976
rect 10100 50930 10314 50964
rect 10486 50930 10700 50964
rect 10100 50918 10700 50930
rect 724 50304 1324 50316
rect 724 50270 938 50304
rect 1110 50270 1324 50304
rect 724 50258 1324 50270
rect 1418 50304 2018 50316
rect 1418 50270 1632 50304
rect 1804 50270 2018 50304
rect 1418 50258 2018 50270
rect 2112 50304 2712 50316
rect 2112 50270 2326 50304
rect 2498 50270 2712 50304
rect 2112 50258 2712 50270
rect 11366 50958 11966 50970
rect 11366 50924 11580 50958
rect 11752 50924 11966 50958
rect 11366 50912 11966 50924
rect 12060 50958 12660 50970
rect 12060 50924 12274 50958
rect 12446 50924 12660 50958
rect 12060 50912 12660 50924
rect 12754 50958 13354 50970
rect 12754 50924 12968 50958
rect 13140 50924 13354 50958
rect 12754 50912 13354 50924
rect 14020 50964 14620 50976
rect 14020 50930 14234 50964
rect 14406 50930 14620 50964
rect 14020 50918 14620 50930
rect 14714 50964 15314 50976
rect 14714 50930 14928 50964
rect 15100 50930 15314 50964
rect 14714 50918 15314 50930
rect 15408 50964 16008 50976
rect 15408 50930 15622 50964
rect 15794 50930 16008 50964
rect 15408 50918 16008 50930
rect 16646 50968 17246 50980
rect 16646 50934 16860 50968
rect 17032 50934 17246 50968
rect 16646 50922 17246 50934
rect 17340 50968 17940 50980
rect 17340 50934 17554 50968
rect 17726 50934 17940 50968
rect 17340 50922 17940 50934
rect 18034 50968 18634 50980
rect 18034 50934 18248 50968
rect 18420 50934 18634 50968
rect 18034 50922 18634 50934
rect 19330 51012 19930 51024
rect 19330 50978 19544 51012
rect 19716 50978 19930 51012
rect 19330 50966 19930 50978
rect 20024 51012 20624 51024
rect 20024 50978 20238 51012
rect 20410 50978 20624 51012
rect 20024 50966 20624 50978
rect 3392 50300 3992 50312
rect 3392 50266 3606 50300
rect 3778 50266 3992 50300
rect 3392 50254 3992 50266
rect 4086 50300 4686 50312
rect 4086 50266 4300 50300
rect 4472 50266 4686 50300
rect 4086 50254 4686 50266
rect 4780 50300 5380 50312
rect 4780 50266 4994 50300
rect 5166 50266 5380 50300
rect 4780 50254 5380 50266
rect 6066 50306 6666 50318
rect 6066 50272 6280 50306
rect 6452 50272 6666 50306
rect 6066 50260 6666 50272
rect 6760 50306 7360 50318
rect 6760 50272 6974 50306
rect 7146 50272 7360 50306
rect 6760 50260 7360 50272
rect 7454 50306 8054 50318
rect 7454 50272 7668 50306
rect 7840 50272 8054 50306
rect 7454 50260 8054 50272
rect 8712 50306 9312 50318
rect 8712 50272 8926 50306
rect 9098 50272 9312 50306
rect 8712 50260 9312 50272
rect 9406 50306 10006 50318
rect 9406 50272 9620 50306
rect 9792 50272 10006 50306
rect 9406 50260 10006 50272
rect 10100 50306 10700 50318
rect 10100 50272 10314 50306
rect 10486 50272 10700 50306
rect 10100 50260 10700 50272
rect 724 49646 1324 49658
rect 724 49612 938 49646
rect 1110 49612 1324 49646
rect 724 49600 1324 49612
rect 1418 49646 2018 49658
rect 1418 49612 1632 49646
rect 1804 49612 2018 49646
rect 1418 49600 2018 49612
rect 2112 49646 2712 49658
rect 2112 49612 2326 49646
rect 2498 49612 2712 49646
rect 2112 49600 2712 49612
rect 11366 50300 11966 50312
rect 11366 50266 11580 50300
rect 11752 50266 11966 50300
rect 11366 50254 11966 50266
rect 12060 50300 12660 50312
rect 12060 50266 12274 50300
rect 12446 50266 12660 50300
rect 12060 50254 12660 50266
rect 12754 50300 13354 50312
rect 12754 50266 12968 50300
rect 13140 50266 13354 50300
rect 12754 50254 13354 50266
rect 14020 50306 14620 50318
rect 14020 50272 14234 50306
rect 14406 50272 14620 50306
rect 14020 50260 14620 50272
rect 14714 50306 15314 50318
rect 14714 50272 14928 50306
rect 15100 50272 15314 50306
rect 14714 50260 15314 50272
rect 15408 50306 16008 50318
rect 15408 50272 15622 50306
rect 15794 50272 16008 50306
rect 15408 50260 16008 50272
rect 16646 50310 17246 50322
rect 16646 50276 16860 50310
rect 17032 50276 17246 50310
rect 16646 50264 17246 50276
rect 17340 50310 17940 50322
rect 17340 50276 17554 50310
rect 17726 50276 17940 50310
rect 17340 50264 17940 50276
rect 18034 50310 18634 50322
rect 18034 50276 18248 50310
rect 18420 50276 18634 50310
rect 18034 50264 18634 50276
rect 19330 50354 19930 50366
rect 19330 50320 19544 50354
rect 19716 50320 19930 50354
rect 19330 50308 19930 50320
rect 20024 50354 20624 50366
rect 20024 50320 20238 50354
rect 20410 50320 20624 50354
rect 20024 50308 20624 50320
rect 3392 49642 3992 49654
rect 3392 49608 3606 49642
rect 3778 49608 3992 49642
rect 3392 49596 3992 49608
rect 4086 49642 4686 49654
rect 4086 49608 4300 49642
rect 4472 49608 4686 49642
rect 4086 49596 4686 49608
rect 4780 49642 5380 49654
rect 4780 49608 4994 49642
rect 5166 49608 5380 49642
rect 4780 49596 5380 49608
rect 6066 49648 6666 49660
rect 6066 49614 6280 49648
rect 6452 49614 6666 49648
rect 6066 49602 6666 49614
rect 6760 49648 7360 49660
rect 6760 49614 6974 49648
rect 7146 49614 7360 49648
rect 6760 49602 7360 49614
rect 7454 49648 8054 49660
rect 7454 49614 7668 49648
rect 7840 49614 8054 49648
rect 7454 49602 8054 49614
rect 8712 49648 9312 49660
rect 8712 49614 8926 49648
rect 9098 49614 9312 49648
rect 8712 49602 9312 49614
rect 9406 49648 10006 49660
rect 9406 49614 9620 49648
rect 9792 49614 10006 49648
rect 9406 49602 10006 49614
rect 10100 49648 10700 49660
rect 10100 49614 10314 49648
rect 10486 49614 10700 49648
rect 10100 49602 10700 49614
rect 724 48988 1324 49000
rect 724 48954 938 48988
rect 1110 48954 1324 48988
rect 724 48942 1324 48954
rect 1418 48988 2018 49000
rect 1418 48954 1632 48988
rect 1804 48954 2018 48988
rect 1418 48942 2018 48954
rect 2112 48988 2712 49000
rect 2112 48954 2326 48988
rect 2498 48954 2712 48988
rect 2112 48942 2712 48954
rect 11366 49642 11966 49654
rect 11366 49608 11580 49642
rect 11752 49608 11966 49642
rect 11366 49596 11966 49608
rect 12060 49642 12660 49654
rect 12060 49608 12274 49642
rect 12446 49608 12660 49642
rect 12060 49596 12660 49608
rect 12754 49642 13354 49654
rect 12754 49608 12968 49642
rect 13140 49608 13354 49642
rect 12754 49596 13354 49608
rect 14020 49648 14620 49660
rect 14020 49614 14234 49648
rect 14406 49614 14620 49648
rect 14020 49602 14620 49614
rect 14714 49648 15314 49660
rect 14714 49614 14928 49648
rect 15100 49614 15314 49648
rect 14714 49602 15314 49614
rect 15408 49648 16008 49660
rect 15408 49614 15622 49648
rect 15794 49614 16008 49648
rect 15408 49602 16008 49614
rect 16646 49652 17246 49664
rect 16646 49618 16860 49652
rect 17032 49618 17246 49652
rect 16646 49606 17246 49618
rect 17340 49652 17940 49664
rect 17340 49618 17554 49652
rect 17726 49618 17940 49652
rect 17340 49606 17940 49618
rect 18034 49652 18634 49664
rect 18034 49618 18248 49652
rect 18420 49618 18634 49652
rect 18034 49606 18634 49618
rect 19330 49696 19930 49708
rect 19330 49662 19544 49696
rect 19716 49662 19930 49696
rect 19330 49650 19930 49662
rect 20024 49696 20624 49708
rect 20024 49662 20238 49696
rect 20410 49662 20624 49696
rect 20024 49650 20624 49662
rect 3392 48984 3992 48996
rect 3392 48950 3606 48984
rect 3778 48950 3992 48984
rect 3392 48938 3992 48950
rect 4086 48984 4686 48996
rect 4086 48950 4300 48984
rect 4472 48950 4686 48984
rect 4086 48938 4686 48950
rect 4780 48984 5380 48996
rect 4780 48950 4994 48984
rect 5166 48950 5380 48984
rect 4780 48938 5380 48950
rect 6066 48990 6666 49002
rect 6066 48956 6280 48990
rect 6452 48956 6666 48990
rect 6066 48944 6666 48956
rect 6760 48990 7360 49002
rect 6760 48956 6974 48990
rect 7146 48956 7360 48990
rect 6760 48944 7360 48956
rect 7454 48990 8054 49002
rect 7454 48956 7668 48990
rect 7840 48956 8054 48990
rect 7454 48944 8054 48956
rect 8712 48990 9312 49002
rect 8712 48956 8926 48990
rect 9098 48956 9312 48990
rect 8712 48944 9312 48956
rect 9406 48990 10006 49002
rect 9406 48956 9620 48990
rect 9792 48956 10006 48990
rect 9406 48944 10006 48956
rect 10100 48990 10700 49002
rect 10100 48956 10314 48990
rect 10486 48956 10700 48990
rect 10100 48944 10700 48956
rect 724 48330 1324 48342
rect 724 48296 938 48330
rect 1110 48296 1324 48330
rect 724 48284 1324 48296
rect 1418 48330 2018 48342
rect 1418 48296 1632 48330
rect 1804 48296 2018 48330
rect 1418 48284 2018 48296
rect 2112 48330 2712 48342
rect 2112 48296 2326 48330
rect 2498 48296 2712 48330
rect 2112 48284 2712 48296
rect 11366 48984 11966 48996
rect 11366 48950 11580 48984
rect 11752 48950 11966 48984
rect 11366 48938 11966 48950
rect 12060 48984 12660 48996
rect 12060 48950 12274 48984
rect 12446 48950 12660 48984
rect 12060 48938 12660 48950
rect 12754 48984 13354 48996
rect 12754 48950 12968 48984
rect 13140 48950 13354 48984
rect 12754 48938 13354 48950
rect 14020 48990 14620 49002
rect 14020 48956 14234 48990
rect 14406 48956 14620 48990
rect 14020 48944 14620 48956
rect 14714 48990 15314 49002
rect 14714 48956 14928 48990
rect 15100 48956 15314 48990
rect 14714 48944 15314 48956
rect 15408 48990 16008 49002
rect 15408 48956 15622 48990
rect 15794 48956 16008 48990
rect 15408 48944 16008 48956
rect 16646 48994 17246 49006
rect 16646 48960 16860 48994
rect 17032 48960 17246 48994
rect 16646 48948 17246 48960
rect 17340 48994 17940 49006
rect 17340 48960 17554 48994
rect 17726 48960 17940 48994
rect 17340 48948 17940 48960
rect 18034 48994 18634 49006
rect 18034 48960 18248 48994
rect 18420 48960 18634 48994
rect 18034 48948 18634 48960
rect 19330 49038 19930 49050
rect 19330 49004 19544 49038
rect 19716 49004 19930 49038
rect 19330 48992 19930 49004
rect 20024 49038 20624 49050
rect 20024 49004 20238 49038
rect 20410 49004 20624 49038
rect 20024 48992 20624 49004
rect 3392 48326 3992 48338
rect 3392 48292 3606 48326
rect 3778 48292 3992 48326
rect 3392 48280 3992 48292
rect 4086 48326 4686 48338
rect 4086 48292 4300 48326
rect 4472 48292 4686 48326
rect 4086 48280 4686 48292
rect 4780 48326 5380 48338
rect 4780 48292 4994 48326
rect 5166 48292 5380 48326
rect 4780 48280 5380 48292
rect 6066 48332 6666 48344
rect 6066 48298 6280 48332
rect 6452 48298 6666 48332
rect 6066 48286 6666 48298
rect 6760 48332 7360 48344
rect 6760 48298 6974 48332
rect 7146 48298 7360 48332
rect 6760 48286 7360 48298
rect 7454 48332 8054 48344
rect 7454 48298 7668 48332
rect 7840 48298 8054 48332
rect 7454 48286 8054 48298
rect 8712 48332 9312 48344
rect 8712 48298 8926 48332
rect 9098 48298 9312 48332
rect 8712 48286 9312 48298
rect 9406 48332 10006 48344
rect 9406 48298 9620 48332
rect 9792 48298 10006 48332
rect 9406 48286 10006 48298
rect 10100 48332 10700 48344
rect 10100 48298 10314 48332
rect 10486 48298 10700 48332
rect 10100 48286 10700 48298
rect 724 47672 1324 47684
rect 724 47638 938 47672
rect 1110 47638 1324 47672
rect 724 47626 1324 47638
rect 1418 47672 2018 47684
rect 1418 47638 1632 47672
rect 1804 47638 2018 47672
rect 1418 47626 2018 47638
rect 2112 47672 2712 47684
rect 11366 48326 11966 48338
rect 11366 48292 11580 48326
rect 11752 48292 11966 48326
rect 11366 48280 11966 48292
rect 12060 48326 12660 48338
rect 12060 48292 12274 48326
rect 12446 48292 12660 48326
rect 12060 48280 12660 48292
rect 12754 48326 13354 48338
rect 12754 48292 12968 48326
rect 13140 48292 13354 48326
rect 12754 48280 13354 48292
rect 14020 48332 14620 48344
rect 14020 48298 14234 48332
rect 14406 48298 14620 48332
rect 14020 48286 14620 48298
rect 14714 48332 15314 48344
rect 14714 48298 14928 48332
rect 15100 48298 15314 48332
rect 14714 48286 15314 48298
rect 15408 48332 16008 48344
rect 15408 48298 15622 48332
rect 15794 48298 16008 48332
rect 15408 48286 16008 48298
rect 16646 48336 17246 48348
rect 16646 48302 16860 48336
rect 17032 48302 17246 48336
rect 16646 48290 17246 48302
rect 17340 48336 17940 48348
rect 17340 48302 17554 48336
rect 17726 48302 17940 48336
rect 17340 48290 17940 48302
rect 18034 48336 18634 48348
rect 18034 48302 18248 48336
rect 18420 48302 18634 48336
rect 18034 48290 18634 48302
rect 19330 48380 19930 48392
rect 19330 48346 19544 48380
rect 19716 48346 19930 48380
rect 19330 48334 19930 48346
rect 20024 48380 20624 48392
rect 20024 48346 20238 48380
rect 20410 48346 20624 48380
rect 20024 48334 20624 48346
rect 2112 47638 2326 47672
rect 2498 47638 2712 47672
rect 2112 47626 2712 47638
rect 3392 47668 3992 47680
rect 3392 47634 3606 47668
rect 3778 47634 3992 47668
rect 3392 47622 3992 47634
rect 4086 47668 4686 47680
rect 4086 47634 4300 47668
rect 4472 47634 4686 47668
rect 4086 47622 4686 47634
rect 4780 47668 5380 47680
rect 4780 47634 4994 47668
rect 5166 47634 5380 47668
rect 4780 47622 5380 47634
rect 6066 47674 6666 47686
rect 6066 47640 6280 47674
rect 6452 47640 6666 47674
rect 6066 47628 6666 47640
rect 6760 47674 7360 47686
rect 6760 47640 6974 47674
rect 7146 47640 7360 47674
rect 6760 47628 7360 47640
rect 7454 47674 8054 47686
rect 7454 47640 7668 47674
rect 7840 47640 8054 47674
rect 7454 47628 8054 47640
rect 8712 47674 9312 47686
rect 8712 47640 8926 47674
rect 9098 47640 9312 47674
rect 8712 47628 9312 47640
rect 9406 47674 10006 47686
rect 9406 47640 9620 47674
rect 9792 47640 10006 47674
rect 9406 47628 10006 47640
rect 10100 47674 10700 47686
rect 19330 47722 19930 47734
rect 10100 47640 10314 47674
rect 10486 47640 10700 47674
rect 10100 47628 10700 47640
rect 11366 47668 11966 47680
rect 11366 47634 11580 47668
rect 11752 47634 11966 47668
rect 11366 47622 11966 47634
rect 12060 47668 12660 47680
rect 12060 47634 12274 47668
rect 12446 47634 12660 47668
rect 12060 47622 12660 47634
rect 12754 47668 13354 47680
rect 12754 47634 12968 47668
rect 13140 47634 13354 47668
rect 12754 47622 13354 47634
rect 14020 47674 14620 47686
rect 14020 47640 14234 47674
rect 14406 47640 14620 47674
rect 14020 47628 14620 47640
rect 14714 47674 15314 47686
rect 14714 47640 14928 47674
rect 15100 47640 15314 47674
rect 14714 47628 15314 47640
rect 15408 47674 16008 47686
rect 15408 47640 15622 47674
rect 15794 47640 16008 47674
rect 15408 47628 16008 47640
rect 16646 47678 17246 47690
rect 16646 47644 16860 47678
rect 17032 47644 17246 47678
rect 16646 47632 17246 47644
rect 17340 47678 17940 47690
rect 17340 47644 17554 47678
rect 17726 47644 17940 47678
rect 17340 47632 17940 47644
rect 18034 47678 18634 47690
rect 18034 47644 18248 47678
rect 18420 47644 18634 47678
rect 19330 47688 19544 47722
rect 19716 47688 19930 47722
rect 19330 47676 19930 47688
rect 20024 47722 20624 47734
rect 20024 47688 20238 47722
rect 20410 47688 20624 47722
rect 20024 47676 20624 47688
rect 18034 47632 18634 47644
rect 42188 65740 42788 65752
rect 42188 65706 42402 65740
rect 42574 65706 42788 65740
rect 42188 65694 42788 65706
rect 42882 65740 43482 65752
rect 42882 65706 43096 65740
rect 43268 65706 43482 65740
rect 42882 65694 43482 65706
rect 43576 65740 44176 65752
rect 43576 65706 43790 65740
rect 43962 65706 44176 65740
rect 43576 65694 44176 65706
rect 44270 65740 44870 65752
rect 44270 65706 44484 65740
rect 44656 65706 44870 65740
rect 44270 65694 44870 65706
rect 44964 65740 45564 65752
rect 44964 65706 45178 65740
rect 45350 65706 45564 65740
rect 44964 65694 45564 65706
rect 46182 65740 46782 65752
rect 46182 65706 46396 65740
rect 46568 65706 46782 65740
rect 46182 65694 46782 65706
rect 46876 65740 47476 65752
rect 46876 65706 47090 65740
rect 47262 65706 47476 65740
rect 46876 65694 47476 65706
rect 47570 65740 48170 65752
rect 47570 65706 47784 65740
rect 47956 65706 48170 65740
rect 47570 65694 48170 65706
rect 48264 65740 48864 65752
rect 48264 65706 48478 65740
rect 48650 65706 48864 65740
rect 48264 65694 48864 65706
rect 48958 65740 49558 65752
rect 48958 65706 49172 65740
rect 49344 65706 49558 65740
rect 48958 65694 49558 65706
rect 50204 65740 50804 65752
rect 50204 65706 50418 65740
rect 50590 65706 50804 65740
rect 50204 65694 50804 65706
rect 50898 65740 51498 65752
rect 50898 65706 51112 65740
rect 51284 65706 51498 65740
rect 50898 65694 51498 65706
rect 51592 65740 52192 65752
rect 51592 65706 51806 65740
rect 51978 65706 52192 65740
rect 51592 65694 52192 65706
rect 52286 65740 52886 65752
rect 52286 65706 52500 65740
rect 52672 65706 52886 65740
rect 52286 65694 52886 65706
rect 52980 65740 53580 65752
rect 52980 65706 53194 65740
rect 53366 65706 53580 65740
rect 52980 65694 53580 65706
rect 54226 65740 54826 65752
rect 54226 65706 54440 65740
rect 54612 65706 54826 65740
rect 54226 65694 54826 65706
rect 54920 65740 55520 65752
rect 54920 65706 55134 65740
rect 55306 65706 55520 65740
rect 54920 65694 55520 65706
rect 55614 65740 56214 65752
rect 55614 65706 55828 65740
rect 56000 65706 56214 65740
rect 55614 65694 56214 65706
rect 56308 65740 56908 65752
rect 56308 65706 56522 65740
rect 56694 65706 56908 65740
rect 56308 65694 56908 65706
rect 57002 65740 57602 65752
rect 57002 65706 57216 65740
rect 57388 65706 57602 65740
rect 57002 65694 57602 65706
rect 71294 66402 71306 66574
rect 71340 66402 71352 66574
rect 71294 66188 71352 66402
rect 71952 66574 72010 66788
rect 71952 66402 71964 66574
rect 71998 66402 72010 66574
rect 71952 66188 72010 66402
rect 72610 66574 72668 66788
rect 72610 66402 72622 66574
rect 72656 66402 72668 66574
rect 72610 66188 72668 66402
rect 73268 66574 73326 66788
rect 73268 66402 73280 66574
rect 73314 66402 73326 66574
rect 73268 66188 73326 66402
rect 73926 66574 73984 66788
rect 73926 66402 73938 66574
rect 73972 66402 73984 66574
rect 75158 69158 75170 69330
rect 75204 69158 75216 69330
rect 75158 68944 75216 69158
rect 75816 69330 75874 69544
rect 75816 69158 75828 69330
rect 75862 69158 75874 69330
rect 75816 68944 75874 69158
rect 76474 69330 76532 69544
rect 76474 69158 76486 69330
rect 76520 69158 76532 69330
rect 76474 68944 76532 69158
rect 77132 69330 77190 69544
rect 77132 69158 77144 69330
rect 77178 69158 77190 69330
rect 77132 68944 77190 69158
rect 77790 69330 77848 69544
rect 79008 69344 79066 69558
rect 77790 69158 77802 69330
rect 77836 69158 77848 69330
rect 77790 68944 77848 69158
rect 75158 68636 75216 68850
rect 75158 68464 75170 68636
rect 75204 68464 75216 68636
rect 75158 68250 75216 68464
rect 75816 68636 75874 68850
rect 75816 68464 75828 68636
rect 75862 68464 75874 68636
rect 75816 68250 75874 68464
rect 76474 68636 76532 68850
rect 76474 68464 76486 68636
rect 76520 68464 76532 68636
rect 76474 68250 76532 68464
rect 77132 68636 77190 68850
rect 77132 68464 77144 68636
rect 77178 68464 77190 68636
rect 77132 68250 77190 68464
rect 77790 68636 77848 68850
rect 77790 68464 77802 68636
rect 77836 68464 77848 68636
rect 77790 68250 77848 68464
rect 75158 67942 75216 68156
rect 75158 67770 75170 67942
rect 75204 67770 75216 67942
rect 75158 67556 75216 67770
rect 75816 67942 75874 68156
rect 75816 67770 75828 67942
rect 75862 67770 75874 67942
rect 75816 67556 75874 67770
rect 76474 67942 76532 68156
rect 76474 67770 76486 67942
rect 76520 67770 76532 67942
rect 76474 67556 76532 67770
rect 77132 67942 77190 68156
rect 77132 67770 77144 67942
rect 77178 67770 77190 67942
rect 77132 67556 77190 67770
rect 77790 67942 77848 68156
rect 77790 67770 77802 67942
rect 77836 67770 77848 67942
rect 77790 67556 77848 67770
rect 75158 67248 75216 67462
rect 75158 67076 75170 67248
rect 75204 67076 75216 67248
rect 75158 66862 75216 67076
rect 75816 67248 75874 67462
rect 75816 67076 75828 67248
rect 75862 67076 75874 67248
rect 75816 66862 75874 67076
rect 76474 67248 76532 67462
rect 76474 67076 76486 67248
rect 76520 67076 76532 67248
rect 76474 66862 76532 67076
rect 77132 67248 77190 67462
rect 77132 67076 77144 67248
rect 77178 67076 77190 67248
rect 77132 66862 77190 67076
rect 77790 67248 77848 67462
rect 77790 67076 77802 67248
rect 77836 67076 77848 67248
rect 77790 66862 77848 67076
rect 75158 66554 75216 66768
rect 73926 66188 73984 66402
rect 75158 66382 75170 66554
rect 75204 66382 75216 66554
rect 75158 66168 75216 66382
rect 75816 66554 75874 66768
rect 75816 66382 75828 66554
rect 75862 66382 75874 66554
rect 75816 66168 75874 66382
rect 76474 66554 76532 66768
rect 76474 66382 76486 66554
rect 76520 66382 76532 66554
rect 76474 66168 76532 66382
rect 77132 66554 77190 66768
rect 77132 66382 77144 66554
rect 77178 66382 77190 66554
rect 77132 66168 77190 66382
rect 77790 66554 77848 66768
rect 77790 66382 77802 66554
rect 77836 66382 77848 66554
rect 79008 69172 79020 69344
rect 79054 69172 79066 69344
rect 79008 68958 79066 69172
rect 79666 69344 79724 69558
rect 79666 69172 79678 69344
rect 79712 69172 79724 69344
rect 79666 68958 79724 69172
rect 80324 69344 80382 69558
rect 80324 69172 80336 69344
rect 80370 69172 80382 69344
rect 80324 68958 80382 69172
rect 80982 69344 81040 69558
rect 80982 69172 80994 69344
rect 81028 69172 81040 69344
rect 80982 68958 81040 69172
rect 81640 69344 81698 69558
rect 81640 69172 81652 69344
rect 81686 69172 81698 69344
rect 81640 68958 81698 69172
rect 79008 68650 79066 68864
rect 79008 68478 79020 68650
rect 79054 68478 79066 68650
rect 79008 68264 79066 68478
rect 79666 68650 79724 68864
rect 79666 68478 79678 68650
rect 79712 68478 79724 68650
rect 79666 68264 79724 68478
rect 80324 68650 80382 68864
rect 80324 68478 80336 68650
rect 80370 68478 80382 68650
rect 80324 68264 80382 68478
rect 80982 68650 81040 68864
rect 80982 68478 80994 68650
rect 81028 68478 81040 68650
rect 80982 68264 81040 68478
rect 81640 68650 81698 68864
rect 81640 68478 81652 68650
rect 81686 68478 81698 68650
rect 81640 68264 81698 68478
rect 79008 67956 79066 68170
rect 79008 67784 79020 67956
rect 79054 67784 79066 67956
rect 79008 67570 79066 67784
rect 79666 67956 79724 68170
rect 79666 67784 79678 67956
rect 79712 67784 79724 67956
rect 79666 67570 79724 67784
rect 80324 67956 80382 68170
rect 80324 67784 80336 67956
rect 80370 67784 80382 67956
rect 80324 67570 80382 67784
rect 80982 67956 81040 68170
rect 80982 67784 80994 67956
rect 81028 67784 81040 67956
rect 80982 67570 81040 67784
rect 81640 67956 81698 68170
rect 81640 67784 81652 67956
rect 81686 67784 81698 67956
rect 81640 67570 81698 67784
rect 79008 67262 79066 67476
rect 79008 67090 79020 67262
rect 79054 67090 79066 67262
rect 79008 66876 79066 67090
rect 79666 67262 79724 67476
rect 79666 67090 79678 67262
rect 79712 67090 79724 67262
rect 79666 66876 79724 67090
rect 80324 67262 80382 67476
rect 80324 67090 80336 67262
rect 80370 67090 80382 67262
rect 80324 66876 80382 67090
rect 80982 67262 81040 67476
rect 80982 67090 80994 67262
rect 81028 67090 81040 67262
rect 80982 66876 81040 67090
rect 81640 67262 81698 67476
rect 81640 67090 81652 67262
rect 81686 67090 81698 67262
rect 81640 66876 81698 67090
rect 79008 66568 79066 66782
rect 77790 66168 77848 66382
rect 79008 66396 79020 66568
rect 79054 66396 79066 66568
rect 79008 66182 79066 66396
rect 79666 66568 79724 66782
rect 79666 66396 79678 66568
rect 79712 66396 79724 66568
rect 79666 66182 79724 66396
rect 80324 66568 80382 66782
rect 80324 66396 80336 66568
rect 80370 66396 80382 66568
rect 80324 66182 80382 66396
rect 80982 66568 81040 66782
rect 80982 66396 80994 66568
rect 81028 66396 81040 66568
rect 80982 66182 81040 66396
rect 81640 66568 81698 66782
rect 81640 66396 81652 66568
rect 81686 66396 81698 66568
rect 81640 66182 81698 66396
rect 71294 65580 71352 65794
rect 42176 64556 42776 64568
rect 42176 64522 42390 64556
rect 42562 64522 42776 64556
rect 42176 64510 42776 64522
rect 42870 64556 43470 64568
rect 42870 64522 43084 64556
rect 43256 64522 43470 64556
rect 42870 64510 43470 64522
rect 43564 64556 44164 64568
rect 43564 64522 43778 64556
rect 43950 64522 44164 64556
rect 43564 64510 44164 64522
rect 44258 64556 44858 64568
rect 44258 64522 44472 64556
rect 44644 64522 44858 64556
rect 44258 64510 44858 64522
rect 44952 64556 45552 64568
rect 44952 64522 45166 64556
rect 45338 64522 45552 64556
rect 44952 64510 45552 64522
rect 46184 64554 46784 64566
rect 46184 64520 46398 64554
rect 46570 64520 46784 64554
rect 46184 64508 46784 64520
rect 46878 64554 47478 64566
rect 46878 64520 47092 64554
rect 47264 64520 47478 64554
rect 46878 64508 47478 64520
rect 47572 64554 48172 64566
rect 47572 64520 47786 64554
rect 47958 64520 48172 64554
rect 47572 64508 48172 64520
rect 48266 64554 48866 64566
rect 48266 64520 48480 64554
rect 48652 64520 48866 64554
rect 48266 64508 48866 64520
rect 48960 64554 49560 64566
rect 48960 64520 49174 64554
rect 49346 64520 49560 64554
rect 48960 64508 49560 64520
rect 50196 64554 50796 64566
rect 50196 64520 50410 64554
rect 50582 64520 50796 64554
rect 50196 64508 50796 64520
rect 50890 64554 51490 64566
rect 50890 64520 51104 64554
rect 51276 64520 51490 64554
rect 50890 64508 51490 64520
rect 51584 64554 52184 64566
rect 51584 64520 51798 64554
rect 51970 64520 52184 64554
rect 51584 64508 52184 64520
rect 52278 64554 52878 64566
rect 52278 64520 52492 64554
rect 52664 64520 52878 64554
rect 52278 64508 52878 64520
rect 52972 64554 53572 64566
rect 52972 64520 53186 64554
rect 53358 64520 53572 64554
rect 52972 64508 53572 64520
rect 54206 64554 54806 64566
rect 54206 64520 54420 64554
rect 54592 64520 54806 64554
rect 54206 64508 54806 64520
rect 54900 64554 55500 64566
rect 54900 64520 55114 64554
rect 55286 64520 55500 64554
rect 54900 64508 55500 64520
rect 55594 64554 56194 64566
rect 55594 64520 55808 64554
rect 55980 64520 56194 64554
rect 55594 64508 56194 64520
rect 56288 64554 56888 64566
rect 56288 64520 56502 64554
rect 56674 64520 56888 64554
rect 56288 64508 56888 64520
rect 56982 64554 57582 64566
rect 56982 64520 57196 64554
rect 57368 64520 57582 64554
rect 56982 64508 57582 64520
rect 42176 63898 42776 63910
rect 42176 63864 42390 63898
rect 42562 63864 42776 63898
rect 42176 63852 42776 63864
rect 42870 63898 43470 63910
rect 42870 63864 43084 63898
rect 43256 63864 43470 63898
rect 42870 63852 43470 63864
rect 43564 63898 44164 63910
rect 43564 63864 43778 63898
rect 43950 63864 44164 63898
rect 43564 63852 44164 63864
rect 44258 63898 44858 63910
rect 44258 63864 44472 63898
rect 44644 63864 44858 63898
rect 44258 63852 44858 63864
rect 44952 63898 45552 63910
rect 44952 63864 45166 63898
rect 45338 63864 45552 63898
rect 44952 63852 45552 63864
rect 46184 63896 46784 63908
rect 46184 63862 46398 63896
rect 46570 63862 46784 63896
rect 46184 63850 46784 63862
rect 46878 63896 47478 63908
rect 46878 63862 47092 63896
rect 47264 63862 47478 63896
rect 46878 63850 47478 63862
rect 47572 63896 48172 63908
rect 47572 63862 47786 63896
rect 47958 63862 48172 63896
rect 47572 63850 48172 63862
rect 48266 63896 48866 63908
rect 48266 63862 48480 63896
rect 48652 63862 48866 63896
rect 48266 63850 48866 63862
rect 48960 63896 49560 63908
rect 48960 63862 49174 63896
rect 49346 63862 49560 63896
rect 48960 63850 49560 63862
rect 50196 63896 50796 63908
rect 50196 63862 50410 63896
rect 50582 63862 50796 63896
rect 50196 63850 50796 63862
rect 50890 63896 51490 63908
rect 50890 63862 51104 63896
rect 51276 63862 51490 63896
rect 50890 63850 51490 63862
rect 51584 63896 52184 63908
rect 51584 63862 51798 63896
rect 51970 63862 52184 63896
rect 51584 63850 52184 63862
rect 52278 63896 52878 63908
rect 52278 63862 52492 63896
rect 52664 63862 52878 63896
rect 52278 63850 52878 63862
rect 52972 63896 53572 63908
rect 52972 63862 53186 63896
rect 53358 63862 53572 63896
rect 52972 63850 53572 63862
rect 54206 63896 54806 63908
rect 54206 63862 54420 63896
rect 54592 63862 54806 63896
rect 54206 63850 54806 63862
rect 54900 63896 55500 63908
rect 54900 63862 55114 63896
rect 55286 63862 55500 63896
rect 54900 63850 55500 63862
rect 55594 63896 56194 63908
rect 55594 63862 55808 63896
rect 55980 63862 56194 63896
rect 55594 63850 56194 63862
rect 56288 63896 56888 63908
rect 56288 63862 56502 63896
rect 56674 63862 56888 63896
rect 56288 63850 56888 63862
rect 56982 63896 57582 63908
rect 56982 63862 57196 63896
rect 57368 63862 57582 63896
rect 56982 63850 57582 63862
rect 42176 63240 42776 63252
rect 42176 63206 42390 63240
rect 42562 63206 42776 63240
rect 42176 63194 42776 63206
rect 42870 63240 43470 63252
rect 42870 63206 43084 63240
rect 43256 63206 43470 63240
rect 42870 63194 43470 63206
rect 43564 63240 44164 63252
rect 43564 63206 43778 63240
rect 43950 63206 44164 63240
rect 43564 63194 44164 63206
rect 44258 63240 44858 63252
rect 44258 63206 44472 63240
rect 44644 63206 44858 63240
rect 44258 63194 44858 63206
rect 44952 63240 45552 63252
rect 44952 63206 45166 63240
rect 45338 63206 45552 63240
rect 44952 63194 45552 63206
rect 46184 63238 46784 63250
rect 46184 63204 46398 63238
rect 46570 63204 46784 63238
rect 46184 63192 46784 63204
rect 46878 63238 47478 63250
rect 46878 63204 47092 63238
rect 47264 63204 47478 63238
rect 46878 63192 47478 63204
rect 47572 63238 48172 63250
rect 47572 63204 47786 63238
rect 47958 63204 48172 63238
rect 47572 63192 48172 63204
rect 48266 63238 48866 63250
rect 48266 63204 48480 63238
rect 48652 63204 48866 63238
rect 48266 63192 48866 63204
rect 48960 63238 49560 63250
rect 48960 63204 49174 63238
rect 49346 63204 49560 63238
rect 48960 63192 49560 63204
rect 50196 63238 50796 63250
rect 50196 63204 50410 63238
rect 50582 63204 50796 63238
rect 50196 63192 50796 63204
rect 50890 63238 51490 63250
rect 50890 63204 51104 63238
rect 51276 63204 51490 63238
rect 50890 63192 51490 63204
rect 51584 63238 52184 63250
rect 51584 63204 51798 63238
rect 51970 63204 52184 63238
rect 51584 63192 52184 63204
rect 52278 63238 52878 63250
rect 52278 63204 52492 63238
rect 52664 63204 52878 63238
rect 52278 63192 52878 63204
rect 52972 63238 53572 63250
rect 52972 63204 53186 63238
rect 53358 63204 53572 63238
rect 52972 63192 53572 63204
rect 54206 63238 54806 63250
rect 54206 63204 54420 63238
rect 54592 63204 54806 63238
rect 54206 63192 54806 63204
rect 54900 63238 55500 63250
rect 54900 63204 55114 63238
rect 55286 63204 55500 63238
rect 54900 63192 55500 63204
rect 55594 63238 56194 63250
rect 55594 63204 55808 63238
rect 55980 63204 56194 63238
rect 55594 63192 56194 63204
rect 56288 63238 56888 63250
rect 56288 63204 56502 63238
rect 56674 63204 56888 63238
rect 56288 63192 56888 63204
rect 56982 63238 57582 63250
rect 56982 63204 57196 63238
rect 57368 63204 57582 63238
rect 56982 63192 57582 63204
rect 42176 62582 42776 62594
rect 42176 62548 42390 62582
rect 42562 62548 42776 62582
rect 42176 62536 42776 62548
rect 42870 62582 43470 62594
rect 42870 62548 43084 62582
rect 43256 62548 43470 62582
rect 42870 62536 43470 62548
rect 43564 62582 44164 62594
rect 43564 62548 43778 62582
rect 43950 62548 44164 62582
rect 43564 62536 44164 62548
rect 44258 62582 44858 62594
rect 44258 62548 44472 62582
rect 44644 62548 44858 62582
rect 44258 62536 44858 62548
rect 44952 62582 45552 62594
rect 44952 62548 45166 62582
rect 45338 62548 45552 62582
rect 44952 62536 45552 62548
rect 46184 62580 46784 62592
rect 46184 62546 46398 62580
rect 46570 62546 46784 62580
rect 46184 62534 46784 62546
rect 46878 62580 47478 62592
rect 46878 62546 47092 62580
rect 47264 62546 47478 62580
rect 46878 62534 47478 62546
rect 47572 62580 48172 62592
rect 47572 62546 47786 62580
rect 47958 62546 48172 62580
rect 47572 62534 48172 62546
rect 48266 62580 48866 62592
rect 48266 62546 48480 62580
rect 48652 62546 48866 62580
rect 48266 62534 48866 62546
rect 48960 62580 49560 62592
rect 48960 62546 49174 62580
rect 49346 62546 49560 62580
rect 48960 62534 49560 62546
rect 50196 62580 50796 62592
rect 50196 62546 50410 62580
rect 50582 62546 50796 62580
rect 50196 62534 50796 62546
rect 50890 62580 51490 62592
rect 50890 62546 51104 62580
rect 51276 62546 51490 62580
rect 50890 62534 51490 62546
rect 51584 62580 52184 62592
rect 51584 62546 51798 62580
rect 51970 62546 52184 62580
rect 51584 62534 52184 62546
rect 52278 62580 52878 62592
rect 52278 62546 52492 62580
rect 52664 62546 52878 62580
rect 52278 62534 52878 62546
rect 52972 62580 53572 62592
rect 52972 62546 53186 62580
rect 53358 62546 53572 62580
rect 52972 62534 53572 62546
rect 54206 62580 54806 62592
rect 54206 62546 54420 62580
rect 54592 62546 54806 62580
rect 54206 62534 54806 62546
rect 54900 62580 55500 62592
rect 54900 62546 55114 62580
rect 55286 62546 55500 62580
rect 54900 62534 55500 62546
rect 55594 62580 56194 62592
rect 55594 62546 55808 62580
rect 55980 62546 56194 62580
rect 55594 62534 56194 62546
rect 56288 62580 56888 62592
rect 56288 62546 56502 62580
rect 56674 62546 56888 62580
rect 56288 62534 56888 62546
rect 56982 62580 57582 62592
rect 56982 62546 57196 62580
rect 57368 62546 57582 62580
rect 56982 62534 57582 62546
rect 42176 61924 42776 61936
rect 42176 61890 42390 61924
rect 42562 61890 42776 61924
rect 42176 61878 42776 61890
rect 42870 61924 43470 61936
rect 42870 61890 43084 61924
rect 43256 61890 43470 61924
rect 42870 61878 43470 61890
rect 43564 61924 44164 61936
rect 43564 61890 43778 61924
rect 43950 61890 44164 61924
rect 43564 61878 44164 61890
rect 44258 61924 44858 61936
rect 44258 61890 44472 61924
rect 44644 61890 44858 61924
rect 44258 61878 44858 61890
rect 44952 61924 45552 61936
rect 44952 61890 45166 61924
rect 45338 61890 45552 61924
rect 44952 61878 45552 61890
rect 71294 65408 71306 65580
rect 71340 65408 71352 65580
rect 71294 65194 71352 65408
rect 71952 65580 72010 65794
rect 71952 65408 71964 65580
rect 71998 65408 72010 65580
rect 71952 65194 72010 65408
rect 72610 65580 72668 65794
rect 72610 65408 72622 65580
rect 72656 65408 72668 65580
rect 72610 65194 72668 65408
rect 73268 65580 73326 65794
rect 73268 65408 73280 65580
rect 73314 65408 73326 65580
rect 73268 65194 73326 65408
rect 73926 65580 73984 65794
rect 73926 65408 73938 65580
rect 73972 65408 73984 65580
rect 75158 65560 75216 65774
rect 73926 65194 73984 65408
rect 71294 64886 71352 65100
rect 71294 64714 71306 64886
rect 71340 64714 71352 64886
rect 71294 64500 71352 64714
rect 71952 64886 72010 65100
rect 71952 64714 71964 64886
rect 71998 64714 72010 64886
rect 71952 64500 72010 64714
rect 72610 64886 72668 65100
rect 72610 64714 72622 64886
rect 72656 64714 72668 64886
rect 72610 64500 72668 64714
rect 73268 64886 73326 65100
rect 73268 64714 73280 64886
rect 73314 64714 73326 64886
rect 73268 64500 73326 64714
rect 73926 64886 73984 65100
rect 73926 64714 73938 64886
rect 73972 64714 73984 64886
rect 73926 64500 73984 64714
rect 71294 64192 71352 64406
rect 71294 64020 71306 64192
rect 71340 64020 71352 64192
rect 71294 63806 71352 64020
rect 71952 64192 72010 64406
rect 71952 64020 71964 64192
rect 71998 64020 72010 64192
rect 71952 63806 72010 64020
rect 72610 64192 72668 64406
rect 72610 64020 72622 64192
rect 72656 64020 72668 64192
rect 72610 63806 72668 64020
rect 73268 64192 73326 64406
rect 73268 64020 73280 64192
rect 73314 64020 73326 64192
rect 73268 63806 73326 64020
rect 73926 64192 73984 64406
rect 73926 64020 73938 64192
rect 73972 64020 73984 64192
rect 73926 63806 73984 64020
rect 71294 63498 71352 63712
rect 71294 63326 71306 63498
rect 71340 63326 71352 63498
rect 71294 63112 71352 63326
rect 71952 63498 72010 63712
rect 71952 63326 71964 63498
rect 71998 63326 72010 63498
rect 71952 63112 72010 63326
rect 72610 63498 72668 63712
rect 72610 63326 72622 63498
rect 72656 63326 72668 63498
rect 72610 63112 72668 63326
rect 73268 63498 73326 63712
rect 73268 63326 73280 63498
rect 73314 63326 73326 63498
rect 73268 63112 73326 63326
rect 73926 63498 73984 63712
rect 73926 63326 73938 63498
rect 73972 63326 73984 63498
rect 73926 63112 73984 63326
rect 46184 61922 46784 61934
rect 46184 61888 46398 61922
rect 46570 61888 46784 61922
rect 46184 61876 46784 61888
rect 46878 61922 47478 61934
rect 46878 61888 47092 61922
rect 47264 61888 47478 61922
rect 46878 61876 47478 61888
rect 47572 61922 48172 61934
rect 47572 61888 47786 61922
rect 47958 61888 48172 61922
rect 47572 61876 48172 61888
rect 48266 61922 48866 61934
rect 48266 61888 48480 61922
rect 48652 61888 48866 61922
rect 48266 61876 48866 61888
rect 48960 61922 49560 61934
rect 48960 61888 49174 61922
rect 49346 61888 49560 61922
rect 48960 61876 49560 61888
rect 50196 61922 50796 61934
rect 50196 61888 50410 61922
rect 50582 61888 50796 61922
rect 50196 61876 50796 61888
rect 50890 61922 51490 61934
rect 50890 61888 51104 61922
rect 51276 61888 51490 61922
rect 50890 61876 51490 61888
rect 51584 61922 52184 61934
rect 51584 61888 51798 61922
rect 51970 61888 52184 61922
rect 51584 61876 52184 61888
rect 52278 61922 52878 61934
rect 52278 61888 52492 61922
rect 52664 61888 52878 61922
rect 52278 61876 52878 61888
rect 52972 61922 53572 61934
rect 52972 61888 53186 61922
rect 53358 61888 53572 61922
rect 52972 61876 53572 61888
rect 54206 61922 54806 61934
rect 54206 61888 54420 61922
rect 54592 61888 54806 61922
rect 54206 61876 54806 61888
rect 54900 61922 55500 61934
rect 54900 61888 55114 61922
rect 55286 61888 55500 61922
rect 54900 61876 55500 61888
rect 55594 61922 56194 61934
rect 55594 61888 55808 61922
rect 55980 61888 56194 61922
rect 55594 61876 56194 61888
rect 56288 61922 56888 61934
rect 56288 61888 56502 61922
rect 56674 61888 56888 61922
rect 56288 61876 56888 61888
rect 56982 61922 57582 61934
rect 56982 61888 57196 61922
rect 57368 61888 57582 61922
rect 56982 61876 57582 61888
rect 42176 61266 42776 61278
rect 42176 61232 42390 61266
rect 42562 61232 42776 61266
rect 42176 61220 42776 61232
rect 42870 61266 43470 61278
rect 42870 61232 43084 61266
rect 43256 61232 43470 61266
rect 42870 61220 43470 61232
rect 43564 61266 44164 61278
rect 43564 61232 43778 61266
rect 43950 61232 44164 61266
rect 43564 61220 44164 61232
rect 44258 61266 44858 61278
rect 44258 61232 44472 61266
rect 44644 61232 44858 61266
rect 44258 61220 44858 61232
rect 44952 61266 45552 61278
rect 71294 62804 71352 63018
rect 71294 62632 71306 62804
rect 71340 62632 71352 62804
rect 71294 62418 71352 62632
rect 71952 62804 72010 63018
rect 71952 62632 71964 62804
rect 71998 62632 72010 62804
rect 71952 62418 72010 62632
rect 72610 62804 72668 63018
rect 72610 62632 72622 62804
rect 72656 62632 72668 62804
rect 72610 62418 72668 62632
rect 73268 62804 73326 63018
rect 73268 62632 73280 62804
rect 73314 62632 73326 62804
rect 73268 62418 73326 62632
rect 73926 62804 73984 63018
rect 73926 62632 73938 62804
rect 73972 62632 73984 62804
rect 75158 65388 75170 65560
rect 75204 65388 75216 65560
rect 75158 65174 75216 65388
rect 75816 65560 75874 65774
rect 75816 65388 75828 65560
rect 75862 65388 75874 65560
rect 75816 65174 75874 65388
rect 76474 65560 76532 65774
rect 76474 65388 76486 65560
rect 76520 65388 76532 65560
rect 76474 65174 76532 65388
rect 77132 65560 77190 65774
rect 77132 65388 77144 65560
rect 77178 65388 77190 65560
rect 77132 65174 77190 65388
rect 77790 65560 77848 65774
rect 79008 65574 79066 65788
rect 77790 65388 77802 65560
rect 77836 65388 77848 65560
rect 77790 65174 77848 65388
rect 75158 64866 75216 65080
rect 75158 64694 75170 64866
rect 75204 64694 75216 64866
rect 75158 64480 75216 64694
rect 75816 64866 75874 65080
rect 75816 64694 75828 64866
rect 75862 64694 75874 64866
rect 75816 64480 75874 64694
rect 76474 64866 76532 65080
rect 76474 64694 76486 64866
rect 76520 64694 76532 64866
rect 76474 64480 76532 64694
rect 77132 64866 77190 65080
rect 77132 64694 77144 64866
rect 77178 64694 77190 64866
rect 77132 64480 77190 64694
rect 77790 64866 77848 65080
rect 77790 64694 77802 64866
rect 77836 64694 77848 64866
rect 77790 64480 77848 64694
rect 75158 64172 75216 64386
rect 75158 64000 75170 64172
rect 75204 64000 75216 64172
rect 75158 63786 75216 64000
rect 75816 64172 75874 64386
rect 75816 64000 75828 64172
rect 75862 64000 75874 64172
rect 75816 63786 75874 64000
rect 76474 64172 76532 64386
rect 76474 64000 76486 64172
rect 76520 64000 76532 64172
rect 76474 63786 76532 64000
rect 77132 64172 77190 64386
rect 77132 64000 77144 64172
rect 77178 64000 77190 64172
rect 77132 63786 77190 64000
rect 77790 64172 77848 64386
rect 77790 64000 77802 64172
rect 77836 64000 77848 64172
rect 77790 63786 77848 64000
rect 75158 63478 75216 63692
rect 75158 63306 75170 63478
rect 75204 63306 75216 63478
rect 75158 63092 75216 63306
rect 75816 63478 75874 63692
rect 75816 63306 75828 63478
rect 75862 63306 75874 63478
rect 75816 63092 75874 63306
rect 76474 63478 76532 63692
rect 76474 63306 76486 63478
rect 76520 63306 76532 63478
rect 76474 63092 76532 63306
rect 77132 63478 77190 63692
rect 77132 63306 77144 63478
rect 77178 63306 77190 63478
rect 77132 63092 77190 63306
rect 77790 63478 77848 63692
rect 77790 63306 77802 63478
rect 77836 63306 77848 63478
rect 77790 63092 77848 63306
rect 75158 62784 75216 62998
rect 73926 62418 73984 62632
rect 75158 62612 75170 62784
rect 75204 62612 75216 62784
rect 75158 62398 75216 62612
rect 75816 62784 75874 62998
rect 75816 62612 75828 62784
rect 75862 62612 75874 62784
rect 75816 62398 75874 62612
rect 76474 62784 76532 62998
rect 76474 62612 76486 62784
rect 76520 62612 76532 62784
rect 76474 62398 76532 62612
rect 77132 62784 77190 62998
rect 77132 62612 77144 62784
rect 77178 62612 77190 62784
rect 77132 62398 77190 62612
rect 77790 62784 77848 62998
rect 77790 62612 77802 62784
rect 77836 62612 77848 62784
rect 79008 65402 79020 65574
rect 79054 65402 79066 65574
rect 79008 65188 79066 65402
rect 79666 65574 79724 65788
rect 79666 65402 79678 65574
rect 79712 65402 79724 65574
rect 79666 65188 79724 65402
rect 80324 65574 80382 65788
rect 80324 65402 80336 65574
rect 80370 65402 80382 65574
rect 80324 65188 80382 65402
rect 80982 65574 81040 65788
rect 80982 65402 80994 65574
rect 81028 65402 81040 65574
rect 80982 65188 81040 65402
rect 81640 65574 81698 65788
rect 81640 65402 81652 65574
rect 81686 65402 81698 65574
rect 81640 65188 81698 65402
rect 79008 64880 79066 65094
rect 79008 64708 79020 64880
rect 79054 64708 79066 64880
rect 79008 64494 79066 64708
rect 79666 64880 79724 65094
rect 79666 64708 79678 64880
rect 79712 64708 79724 64880
rect 79666 64494 79724 64708
rect 80324 64880 80382 65094
rect 80324 64708 80336 64880
rect 80370 64708 80382 64880
rect 80324 64494 80382 64708
rect 80982 64880 81040 65094
rect 80982 64708 80994 64880
rect 81028 64708 81040 64880
rect 80982 64494 81040 64708
rect 81640 64880 81698 65094
rect 81640 64708 81652 64880
rect 81686 64708 81698 64880
rect 81640 64494 81698 64708
rect 79008 64186 79066 64400
rect 79008 64014 79020 64186
rect 79054 64014 79066 64186
rect 79008 63800 79066 64014
rect 79666 64186 79724 64400
rect 79666 64014 79678 64186
rect 79712 64014 79724 64186
rect 79666 63800 79724 64014
rect 80324 64186 80382 64400
rect 80324 64014 80336 64186
rect 80370 64014 80382 64186
rect 80324 63800 80382 64014
rect 80982 64186 81040 64400
rect 80982 64014 80994 64186
rect 81028 64014 81040 64186
rect 80982 63800 81040 64014
rect 81640 64186 81698 64400
rect 81640 64014 81652 64186
rect 81686 64014 81698 64186
rect 81640 63800 81698 64014
rect 79008 63492 79066 63706
rect 79008 63320 79020 63492
rect 79054 63320 79066 63492
rect 79008 63106 79066 63320
rect 79666 63492 79724 63706
rect 79666 63320 79678 63492
rect 79712 63320 79724 63492
rect 79666 63106 79724 63320
rect 80324 63492 80382 63706
rect 80324 63320 80336 63492
rect 80370 63320 80382 63492
rect 80324 63106 80382 63320
rect 80982 63492 81040 63706
rect 80982 63320 80994 63492
rect 81028 63320 81040 63492
rect 80982 63106 81040 63320
rect 81640 63492 81698 63706
rect 81640 63320 81652 63492
rect 81686 63320 81698 63492
rect 81640 63106 81698 63320
rect 79008 62798 79066 63012
rect 77790 62398 77848 62612
rect 79008 62626 79020 62798
rect 79054 62626 79066 62798
rect 79008 62412 79066 62626
rect 79666 62798 79724 63012
rect 79666 62626 79678 62798
rect 79712 62626 79724 62798
rect 79666 62412 79724 62626
rect 80324 62798 80382 63012
rect 80324 62626 80336 62798
rect 80370 62626 80382 62798
rect 80324 62412 80382 62626
rect 80982 62798 81040 63012
rect 80982 62626 80994 62798
rect 81028 62626 81040 62798
rect 80982 62412 81040 62626
rect 81640 62798 81698 63012
rect 81640 62626 81652 62798
rect 81686 62626 81698 62798
rect 81640 62412 81698 62626
rect 44952 61232 45166 61266
rect 45338 61232 45552 61266
rect 44952 61220 45552 61232
rect 46184 61264 46784 61276
rect 46184 61230 46398 61264
rect 46570 61230 46784 61264
rect 46184 61218 46784 61230
rect 46878 61264 47478 61276
rect 46878 61230 47092 61264
rect 47264 61230 47478 61264
rect 46878 61218 47478 61230
rect 47572 61264 48172 61276
rect 47572 61230 47786 61264
rect 47958 61230 48172 61264
rect 47572 61218 48172 61230
rect 48266 61264 48866 61276
rect 48266 61230 48480 61264
rect 48652 61230 48866 61264
rect 48266 61218 48866 61230
rect 48960 61264 49560 61276
rect 48960 61230 49174 61264
rect 49346 61230 49560 61264
rect 48960 61218 49560 61230
rect 50196 61264 50796 61276
rect 50196 61230 50410 61264
rect 50582 61230 50796 61264
rect 50196 61218 50796 61230
rect 50890 61264 51490 61276
rect 50890 61230 51104 61264
rect 51276 61230 51490 61264
rect 50890 61218 51490 61230
rect 51584 61264 52184 61276
rect 51584 61230 51798 61264
rect 51970 61230 52184 61264
rect 51584 61218 52184 61230
rect 52278 61264 52878 61276
rect 52278 61230 52492 61264
rect 52664 61230 52878 61264
rect 52278 61218 52878 61230
rect 52972 61264 53572 61276
rect 52972 61230 53186 61264
rect 53358 61230 53572 61264
rect 52972 61218 53572 61230
rect 54206 61264 54806 61276
rect 54206 61230 54420 61264
rect 54592 61230 54806 61264
rect 54206 61218 54806 61230
rect 54900 61264 55500 61276
rect 54900 61230 55114 61264
rect 55286 61230 55500 61264
rect 54900 61218 55500 61230
rect 55594 61264 56194 61276
rect 55594 61230 55808 61264
rect 55980 61230 56194 61264
rect 55594 61218 56194 61230
rect 56288 61264 56888 61276
rect 56288 61230 56502 61264
rect 56674 61230 56888 61264
rect 56288 61218 56888 61230
rect 56982 61264 57582 61276
rect 56982 61230 57196 61264
rect 57368 61230 57582 61264
rect 56982 61218 57582 61230
rect 42168 60358 42768 60370
rect 42168 60324 42382 60358
rect 42554 60324 42768 60358
rect 42168 60312 42768 60324
rect 42862 60358 43462 60370
rect 42862 60324 43076 60358
rect 43248 60324 43462 60358
rect 42862 60312 43462 60324
rect 43556 60358 44156 60370
rect 43556 60324 43770 60358
rect 43942 60324 44156 60358
rect 43556 60312 44156 60324
rect 44250 60358 44850 60370
rect 44250 60324 44464 60358
rect 44636 60324 44850 60358
rect 44250 60312 44850 60324
rect 44944 60358 45544 60370
rect 44944 60324 45158 60358
rect 45330 60324 45544 60358
rect 44944 60312 45544 60324
rect 46162 60358 46762 60370
rect 46162 60324 46376 60358
rect 46548 60324 46762 60358
rect 46162 60312 46762 60324
rect 46856 60358 47456 60370
rect 46856 60324 47070 60358
rect 47242 60324 47456 60358
rect 46856 60312 47456 60324
rect 47550 60358 48150 60370
rect 47550 60324 47764 60358
rect 47936 60324 48150 60358
rect 47550 60312 48150 60324
rect 48244 60358 48844 60370
rect 48244 60324 48458 60358
rect 48630 60324 48844 60358
rect 48244 60312 48844 60324
rect 48938 60358 49538 60370
rect 48938 60324 49152 60358
rect 49324 60324 49538 60358
rect 48938 60312 49538 60324
rect 50184 60358 50784 60370
rect 50184 60324 50398 60358
rect 50570 60324 50784 60358
rect 50184 60312 50784 60324
rect 50878 60358 51478 60370
rect 50878 60324 51092 60358
rect 51264 60324 51478 60358
rect 50878 60312 51478 60324
rect 51572 60358 52172 60370
rect 51572 60324 51786 60358
rect 51958 60324 52172 60358
rect 51572 60312 52172 60324
rect 52266 60358 52866 60370
rect 52266 60324 52480 60358
rect 52652 60324 52866 60358
rect 52266 60312 52866 60324
rect 52960 60358 53560 60370
rect 52960 60324 53174 60358
rect 53346 60324 53560 60358
rect 52960 60312 53560 60324
rect 54206 60358 54806 60370
rect 54206 60324 54420 60358
rect 54592 60324 54806 60358
rect 54206 60312 54806 60324
rect 54900 60358 55500 60370
rect 54900 60324 55114 60358
rect 55286 60324 55500 60358
rect 54900 60312 55500 60324
rect 55594 60358 56194 60370
rect 55594 60324 55808 60358
rect 55980 60324 56194 60358
rect 55594 60312 56194 60324
rect 56288 60358 56888 60370
rect 56288 60324 56502 60358
rect 56674 60324 56888 60358
rect 56288 60312 56888 60324
rect 56982 60358 57582 60370
rect 56982 60324 57196 60358
rect 57368 60324 57582 60358
rect 56982 60312 57582 60324
rect 42168 59700 42768 59712
rect 42168 59666 42382 59700
rect 42554 59666 42768 59700
rect 42168 59654 42768 59666
rect 42862 59700 43462 59712
rect 42862 59666 43076 59700
rect 43248 59666 43462 59700
rect 42862 59654 43462 59666
rect 43556 59700 44156 59712
rect 43556 59666 43770 59700
rect 43942 59666 44156 59700
rect 43556 59654 44156 59666
rect 44250 59700 44850 59712
rect 44250 59666 44464 59700
rect 44636 59666 44850 59700
rect 44250 59654 44850 59666
rect 44944 59700 45544 59712
rect 44944 59666 45158 59700
rect 45330 59666 45544 59700
rect 44944 59654 45544 59666
rect 46162 59700 46762 59712
rect 46162 59666 46376 59700
rect 46548 59666 46762 59700
rect 46162 59654 46762 59666
rect 46856 59700 47456 59712
rect 46856 59666 47070 59700
rect 47242 59666 47456 59700
rect 46856 59654 47456 59666
rect 47550 59700 48150 59712
rect 47550 59666 47764 59700
rect 47936 59666 48150 59700
rect 47550 59654 48150 59666
rect 48244 59700 48844 59712
rect 48244 59666 48458 59700
rect 48630 59666 48844 59700
rect 48244 59654 48844 59666
rect 48938 59700 49538 59712
rect 48938 59666 49152 59700
rect 49324 59666 49538 59700
rect 48938 59654 49538 59666
rect 50184 59700 50784 59712
rect 50184 59666 50398 59700
rect 50570 59666 50784 59700
rect 50184 59654 50784 59666
rect 50878 59700 51478 59712
rect 50878 59666 51092 59700
rect 51264 59666 51478 59700
rect 50878 59654 51478 59666
rect 51572 59700 52172 59712
rect 51572 59666 51786 59700
rect 51958 59666 52172 59700
rect 51572 59654 52172 59666
rect 52266 59700 52866 59712
rect 52266 59666 52480 59700
rect 52652 59666 52866 59700
rect 52266 59654 52866 59666
rect 52960 59700 53560 59712
rect 52960 59666 53174 59700
rect 53346 59666 53560 59700
rect 52960 59654 53560 59666
rect 54206 59700 54806 59712
rect 54206 59666 54420 59700
rect 54592 59666 54806 59700
rect 54206 59654 54806 59666
rect 54900 59700 55500 59712
rect 54900 59666 55114 59700
rect 55286 59666 55500 59700
rect 54900 59654 55500 59666
rect 55594 59700 56194 59712
rect 55594 59666 55808 59700
rect 55980 59666 56194 59700
rect 55594 59654 56194 59666
rect 56288 59700 56888 59712
rect 56288 59666 56502 59700
rect 56674 59666 56888 59700
rect 56288 59654 56888 59666
rect 56982 59700 57582 59712
rect 56982 59666 57196 59700
rect 57368 59666 57582 59700
rect 56982 59654 57582 59666
rect 42168 59042 42768 59054
rect 42168 59008 42382 59042
rect 42554 59008 42768 59042
rect 42168 58996 42768 59008
rect 42862 59042 43462 59054
rect 42862 59008 43076 59042
rect 43248 59008 43462 59042
rect 42862 58996 43462 59008
rect 43556 59042 44156 59054
rect 43556 59008 43770 59042
rect 43942 59008 44156 59042
rect 43556 58996 44156 59008
rect 44250 59042 44850 59054
rect 44250 59008 44464 59042
rect 44636 59008 44850 59042
rect 44250 58996 44850 59008
rect 44944 59042 45544 59054
rect 44944 59008 45158 59042
rect 45330 59008 45544 59042
rect 44944 58996 45544 59008
rect 46162 59042 46762 59054
rect 46162 59008 46376 59042
rect 46548 59008 46762 59042
rect 46162 58996 46762 59008
rect 46856 59042 47456 59054
rect 46856 59008 47070 59042
rect 47242 59008 47456 59042
rect 46856 58996 47456 59008
rect 47550 59042 48150 59054
rect 47550 59008 47764 59042
rect 47936 59008 48150 59042
rect 47550 58996 48150 59008
rect 48244 59042 48844 59054
rect 48244 59008 48458 59042
rect 48630 59008 48844 59042
rect 48244 58996 48844 59008
rect 48938 59042 49538 59054
rect 48938 59008 49152 59042
rect 49324 59008 49538 59042
rect 48938 58996 49538 59008
rect 50184 59042 50784 59054
rect 50184 59008 50398 59042
rect 50570 59008 50784 59042
rect 50184 58996 50784 59008
rect 50878 59042 51478 59054
rect 50878 59008 51092 59042
rect 51264 59008 51478 59042
rect 50878 58996 51478 59008
rect 51572 59042 52172 59054
rect 51572 59008 51786 59042
rect 51958 59008 52172 59042
rect 51572 58996 52172 59008
rect 52266 59042 52866 59054
rect 52266 59008 52480 59042
rect 52652 59008 52866 59042
rect 52266 58996 52866 59008
rect 52960 59042 53560 59054
rect 52960 59008 53174 59042
rect 53346 59008 53560 59042
rect 52960 58996 53560 59008
rect 54206 59042 54806 59054
rect 54206 59008 54420 59042
rect 54592 59008 54806 59042
rect 54206 58996 54806 59008
rect 54900 59042 55500 59054
rect 54900 59008 55114 59042
rect 55286 59008 55500 59042
rect 54900 58996 55500 59008
rect 55594 59042 56194 59054
rect 55594 59008 55808 59042
rect 55980 59008 56194 59042
rect 55594 58996 56194 59008
rect 56288 59042 56888 59054
rect 56288 59008 56502 59042
rect 56674 59008 56888 59042
rect 56288 58996 56888 59008
rect 56982 59042 57582 59054
rect 56982 59008 57196 59042
rect 57368 59008 57582 59042
rect 56982 58996 57582 59008
rect 42168 58384 42768 58396
rect 42168 58350 42382 58384
rect 42554 58350 42768 58384
rect 42168 58338 42768 58350
rect 42862 58384 43462 58396
rect 42862 58350 43076 58384
rect 43248 58350 43462 58384
rect 42862 58338 43462 58350
rect 43556 58384 44156 58396
rect 43556 58350 43770 58384
rect 43942 58350 44156 58384
rect 43556 58338 44156 58350
rect 44250 58384 44850 58396
rect 44250 58350 44464 58384
rect 44636 58350 44850 58384
rect 44250 58338 44850 58350
rect 44944 58384 45544 58396
rect 44944 58350 45158 58384
rect 45330 58350 45544 58384
rect 44944 58338 45544 58350
rect 46162 58384 46762 58396
rect 46162 58350 46376 58384
rect 46548 58350 46762 58384
rect 46162 58338 46762 58350
rect 46856 58384 47456 58396
rect 46856 58350 47070 58384
rect 47242 58350 47456 58384
rect 46856 58338 47456 58350
rect 47550 58384 48150 58396
rect 47550 58350 47764 58384
rect 47936 58350 48150 58384
rect 47550 58338 48150 58350
rect 48244 58384 48844 58396
rect 48244 58350 48458 58384
rect 48630 58350 48844 58384
rect 48244 58338 48844 58350
rect 48938 58384 49538 58396
rect 48938 58350 49152 58384
rect 49324 58350 49538 58384
rect 48938 58338 49538 58350
rect 50184 58384 50784 58396
rect 50184 58350 50398 58384
rect 50570 58350 50784 58384
rect 50184 58338 50784 58350
rect 50878 58384 51478 58396
rect 50878 58350 51092 58384
rect 51264 58350 51478 58384
rect 50878 58338 51478 58350
rect 51572 58384 52172 58396
rect 51572 58350 51786 58384
rect 51958 58350 52172 58384
rect 51572 58338 52172 58350
rect 52266 58384 52866 58396
rect 52266 58350 52480 58384
rect 52652 58350 52866 58384
rect 52266 58338 52866 58350
rect 52960 58384 53560 58396
rect 52960 58350 53174 58384
rect 53346 58350 53560 58384
rect 52960 58338 53560 58350
rect 54206 58384 54806 58396
rect 54206 58350 54420 58384
rect 54592 58350 54806 58384
rect 54206 58338 54806 58350
rect 54900 58384 55500 58396
rect 54900 58350 55114 58384
rect 55286 58350 55500 58384
rect 54900 58338 55500 58350
rect 55594 58384 56194 58396
rect 55594 58350 55808 58384
rect 55980 58350 56194 58384
rect 55594 58338 56194 58350
rect 56288 58384 56888 58396
rect 56288 58350 56502 58384
rect 56674 58350 56888 58384
rect 56288 58338 56888 58350
rect 56982 58384 57582 58396
rect 56982 58350 57196 58384
rect 57368 58350 57582 58384
rect 56982 58338 57582 58350
rect 42168 57726 42768 57738
rect 42168 57692 42382 57726
rect 42554 57692 42768 57726
rect 42168 57680 42768 57692
rect 42862 57726 43462 57738
rect 42862 57692 43076 57726
rect 43248 57692 43462 57726
rect 42862 57680 43462 57692
rect 43556 57726 44156 57738
rect 43556 57692 43770 57726
rect 43942 57692 44156 57726
rect 43556 57680 44156 57692
rect 44250 57726 44850 57738
rect 44250 57692 44464 57726
rect 44636 57692 44850 57726
rect 44250 57680 44850 57692
rect 44944 57726 45544 57738
rect 44944 57692 45158 57726
rect 45330 57692 45544 57726
rect 44944 57680 45544 57692
rect 46162 57726 46762 57738
rect 46162 57692 46376 57726
rect 46548 57692 46762 57726
rect 46162 57680 46762 57692
rect 46856 57726 47456 57738
rect 46856 57692 47070 57726
rect 47242 57692 47456 57726
rect 46856 57680 47456 57692
rect 47550 57726 48150 57738
rect 47550 57692 47764 57726
rect 47936 57692 48150 57726
rect 47550 57680 48150 57692
rect 48244 57726 48844 57738
rect 48244 57692 48458 57726
rect 48630 57692 48844 57726
rect 48244 57680 48844 57692
rect 48938 57726 49538 57738
rect 48938 57692 49152 57726
rect 49324 57692 49538 57726
rect 48938 57680 49538 57692
rect 50184 57726 50784 57738
rect 50184 57692 50398 57726
rect 50570 57692 50784 57726
rect 50184 57680 50784 57692
rect 50878 57726 51478 57738
rect 50878 57692 51092 57726
rect 51264 57692 51478 57726
rect 50878 57680 51478 57692
rect 51572 57726 52172 57738
rect 51572 57692 51786 57726
rect 51958 57692 52172 57726
rect 51572 57680 52172 57692
rect 52266 57726 52866 57738
rect 52266 57692 52480 57726
rect 52652 57692 52866 57726
rect 52266 57680 52866 57692
rect 52960 57726 53560 57738
rect 52960 57692 53174 57726
rect 53346 57692 53560 57726
rect 52960 57680 53560 57692
rect 54206 57726 54806 57738
rect 54206 57692 54420 57726
rect 54592 57692 54806 57726
rect 54206 57680 54806 57692
rect 54900 57726 55500 57738
rect 54900 57692 55114 57726
rect 55286 57692 55500 57726
rect 54900 57680 55500 57692
rect 55594 57726 56194 57738
rect 55594 57692 55808 57726
rect 55980 57692 56194 57726
rect 55594 57680 56194 57692
rect 56288 57726 56888 57738
rect 56288 57692 56502 57726
rect 56674 57692 56888 57726
rect 56288 57680 56888 57692
rect 56982 57726 57582 57738
rect 56982 57692 57196 57726
rect 57368 57692 57582 57726
rect 56982 57680 57582 57692
rect 71294 61816 71352 62030
rect 71294 61644 71306 61816
rect 71340 61644 71352 61816
rect 71294 61430 71352 61644
rect 71952 61816 72010 62030
rect 71952 61644 71964 61816
rect 71998 61644 72010 61816
rect 71952 61430 72010 61644
rect 72610 61816 72668 62030
rect 72610 61644 72622 61816
rect 72656 61644 72668 61816
rect 72610 61430 72668 61644
rect 73268 61816 73326 62030
rect 73268 61644 73280 61816
rect 73314 61644 73326 61816
rect 73268 61430 73326 61644
rect 73926 61816 73984 62030
rect 73926 61644 73938 61816
rect 73972 61644 73984 61816
rect 75158 61796 75216 62010
rect 73926 61430 73984 61644
rect 71294 61122 71352 61336
rect 71294 60950 71306 61122
rect 71340 60950 71352 61122
rect 71294 60736 71352 60950
rect 71952 61122 72010 61336
rect 71952 60950 71964 61122
rect 71998 60950 72010 61122
rect 71952 60736 72010 60950
rect 72610 61122 72668 61336
rect 72610 60950 72622 61122
rect 72656 60950 72668 61122
rect 72610 60736 72668 60950
rect 73268 61122 73326 61336
rect 73268 60950 73280 61122
rect 73314 60950 73326 61122
rect 73268 60736 73326 60950
rect 73926 61122 73984 61336
rect 73926 60950 73938 61122
rect 73972 60950 73984 61122
rect 73926 60736 73984 60950
rect 71294 60428 71352 60642
rect 71294 60256 71306 60428
rect 71340 60256 71352 60428
rect 71294 60042 71352 60256
rect 71952 60428 72010 60642
rect 71952 60256 71964 60428
rect 71998 60256 72010 60428
rect 71952 60042 72010 60256
rect 72610 60428 72668 60642
rect 72610 60256 72622 60428
rect 72656 60256 72668 60428
rect 72610 60042 72668 60256
rect 73268 60428 73326 60642
rect 73268 60256 73280 60428
rect 73314 60256 73326 60428
rect 73268 60042 73326 60256
rect 73926 60428 73984 60642
rect 73926 60256 73938 60428
rect 73972 60256 73984 60428
rect 73926 60042 73984 60256
rect 71294 59734 71352 59948
rect 71294 59562 71306 59734
rect 71340 59562 71352 59734
rect 71294 59348 71352 59562
rect 71952 59734 72010 59948
rect 71952 59562 71964 59734
rect 71998 59562 72010 59734
rect 71952 59348 72010 59562
rect 72610 59734 72668 59948
rect 72610 59562 72622 59734
rect 72656 59562 72668 59734
rect 72610 59348 72668 59562
rect 73268 59734 73326 59948
rect 73268 59562 73280 59734
rect 73314 59562 73326 59734
rect 73268 59348 73326 59562
rect 73926 59734 73984 59948
rect 73926 59562 73938 59734
rect 73972 59562 73984 59734
rect 73926 59348 73984 59562
rect 71294 59040 71352 59254
rect 71294 58868 71306 59040
rect 71340 58868 71352 59040
rect 71294 58654 71352 58868
rect 71952 59040 72010 59254
rect 71952 58868 71964 59040
rect 71998 58868 72010 59040
rect 71952 58654 72010 58868
rect 72610 59040 72668 59254
rect 72610 58868 72622 59040
rect 72656 58868 72668 59040
rect 72610 58654 72668 58868
rect 73268 59040 73326 59254
rect 73268 58868 73280 59040
rect 73314 58868 73326 59040
rect 73268 58654 73326 58868
rect 73926 59040 73984 59254
rect 73926 58868 73938 59040
rect 73972 58868 73984 59040
rect 75158 61624 75170 61796
rect 75204 61624 75216 61796
rect 75158 61410 75216 61624
rect 75816 61796 75874 62010
rect 75816 61624 75828 61796
rect 75862 61624 75874 61796
rect 75816 61410 75874 61624
rect 76474 61796 76532 62010
rect 76474 61624 76486 61796
rect 76520 61624 76532 61796
rect 76474 61410 76532 61624
rect 77132 61796 77190 62010
rect 77132 61624 77144 61796
rect 77178 61624 77190 61796
rect 77132 61410 77190 61624
rect 77790 61796 77848 62010
rect 79008 61810 79066 62024
rect 77790 61624 77802 61796
rect 77836 61624 77848 61796
rect 77790 61410 77848 61624
rect 75158 61102 75216 61316
rect 75158 60930 75170 61102
rect 75204 60930 75216 61102
rect 75158 60716 75216 60930
rect 75816 61102 75874 61316
rect 75816 60930 75828 61102
rect 75862 60930 75874 61102
rect 75816 60716 75874 60930
rect 76474 61102 76532 61316
rect 76474 60930 76486 61102
rect 76520 60930 76532 61102
rect 76474 60716 76532 60930
rect 77132 61102 77190 61316
rect 77132 60930 77144 61102
rect 77178 60930 77190 61102
rect 77132 60716 77190 60930
rect 77790 61102 77848 61316
rect 77790 60930 77802 61102
rect 77836 60930 77848 61102
rect 77790 60716 77848 60930
rect 75158 60408 75216 60622
rect 75158 60236 75170 60408
rect 75204 60236 75216 60408
rect 75158 60022 75216 60236
rect 75816 60408 75874 60622
rect 75816 60236 75828 60408
rect 75862 60236 75874 60408
rect 75816 60022 75874 60236
rect 76474 60408 76532 60622
rect 76474 60236 76486 60408
rect 76520 60236 76532 60408
rect 76474 60022 76532 60236
rect 77132 60408 77190 60622
rect 77132 60236 77144 60408
rect 77178 60236 77190 60408
rect 77132 60022 77190 60236
rect 77790 60408 77848 60622
rect 77790 60236 77802 60408
rect 77836 60236 77848 60408
rect 77790 60022 77848 60236
rect 75158 59714 75216 59928
rect 75158 59542 75170 59714
rect 75204 59542 75216 59714
rect 75158 59328 75216 59542
rect 75816 59714 75874 59928
rect 75816 59542 75828 59714
rect 75862 59542 75874 59714
rect 75816 59328 75874 59542
rect 76474 59714 76532 59928
rect 76474 59542 76486 59714
rect 76520 59542 76532 59714
rect 76474 59328 76532 59542
rect 77132 59714 77190 59928
rect 77132 59542 77144 59714
rect 77178 59542 77190 59714
rect 77132 59328 77190 59542
rect 77790 59714 77848 59928
rect 77790 59542 77802 59714
rect 77836 59542 77848 59714
rect 77790 59328 77848 59542
rect 75158 59020 75216 59234
rect 73926 58654 73984 58868
rect 75158 58848 75170 59020
rect 75204 58848 75216 59020
rect 75158 58634 75216 58848
rect 75816 59020 75874 59234
rect 75816 58848 75828 59020
rect 75862 58848 75874 59020
rect 75816 58634 75874 58848
rect 76474 59020 76532 59234
rect 76474 58848 76486 59020
rect 76520 58848 76532 59020
rect 76474 58634 76532 58848
rect 77132 59020 77190 59234
rect 77132 58848 77144 59020
rect 77178 58848 77190 59020
rect 77132 58634 77190 58848
rect 77790 59020 77848 59234
rect 77790 58848 77802 59020
rect 77836 58848 77848 59020
rect 79008 61638 79020 61810
rect 79054 61638 79066 61810
rect 79008 61424 79066 61638
rect 79666 61810 79724 62024
rect 79666 61638 79678 61810
rect 79712 61638 79724 61810
rect 79666 61424 79724 61638
rect 80324 61810 80382 62024
rect 80324 61638 80336 61810
rect 80370 61638 80382 61810
rect 80324 61424 80382 61638
rect 80982 61810 81040 62024
rect 80982 61638 80994 61810
rect 81028 61638 81040 61810
rect 80982 61424 81040 61638
rect 81640 61810 81698 62024
rect 81640 61638 81652 61810
rect 81686 61638 81698 61810
rect 81640 61424 81698 61638
rect 79008 61116 79066 61330
rect 79008 60944 79020 61116
rect 79054 60944 79066 61116
rect 79008 60730 79066 60944
rect 79666 61116 79724 61330
rect 79666 60944 79678 61116
rect 79712 60944 79724 61116
rect 79666 60730 79724 60944
rect 80324 61116 80382 61330
rect 80324 60944 80336 61116
rect 80370 60944 80382 61116
rect 80324 60730 80382 60944
rect 80982 61116 81040 61330
rect 80982 60944 80994 61116
rect 81028 60944 81040 61116
rect 80982 60730 81040 60944
rect 81640 61116 81698 61330
rect 81640 60944 81652 61116
rect 81686 60944 81698 61116
rect 81640 60730 81698 60944
rect 79008 60422 79066 60636
rect 79008 60250 79020 60422
rect 79054 60250 79066 60422
rect 79008 60036 79066 60250
rect 79666 60422 79724 60636
rect 79666 60250 79678 60422
rect 79712 60250 79724 60422
rect 79666 60036 79724 60250
rect 80324 60422 80382 60636
rect 80324 60250 80336 60422
rect 80370 60250 80382 60422
rect 80324 60036 80382 60250
rect 80982 60422 81040 60636
rect 80982 60250 80994 60422
rect 81028 60250 81040 60422
rect 80982 60036 81040 60250
rect 81640 60422 81698 60636
rect 81640 60250 81652 60422
rect 81686 60250 81698 60422
rect 81640 60036 81698 60250
rect 79008 59728 79066 59942
rect 79008 59556 79020 59728
rect 79054 59556 79066 59728
rect 79008 59342 79066 59556
rect 79666 59728 79724 59942
rect 79666 59556 79678 59728
rect 79712 59556 79724 59728
rect 79666 59342 79724 59556
rect 80324 59728 80382 59942
rect 80324 59556 80336 59728
rect 80370 59556 80382 59728
rect 80324 59342 80382 59556
rect 80982 59728 81040 59942
rect 80982 59556 80994 59728
rect 81028 59556 81040 59728
rect 80982 59342 81040 59556
rect 81640 59728 81698 59942
rect 81640 59556 81652 59728
rect 81686 59556 81698 59728
rect 81640 59342 81698 59556
rect 79008 59034 79066 59248
rect 77790 58634 77848 58848
rect 79008 58862 79020 59034
rect 79054 58862 79066 59034
rect 79008 58648 79066 58862
rect 79666 59034 79724 59248
rect 79666 58862 79678 59034
rect 79712 58862 79724 59034
rect 79666 58648 79724 58862
rect 80324 59034 80382 59248
rect 80324 58862 80336 59034
rect 80370 58862 80382 59034
rect 80324 58648 80382 58862
rect 80982 59034 81040 59248
rect 80982 58862 80994 59034
rect 81028 58862 81040 59034
rect 80982 58648 81040 58862
rect 81640 59034 81698 59248
rect 81640 58862 81652 59034
rect 81686 58862 81698 59034
rect 81640 58648 81698 58862
rect 42168 57068 42768 57080
rect 42168 57034 42382 57068
rect 42554 57034 42768 57068
rect 42168 57022 42768 57034
rect 42862 57068 43462 57080
rect 42862 57034 43076 57068
rect 43248 57034 43462 57068
rect 42862 57022 43462 57034
rect 43556 57068 44156 57080
rect 43556 57034 43770 57068
rect 43942 57034 44156 57068
rect 43556 57022 44156 57034
rect 44250 57068 44850 57080
rect 44250 57034 44464 57068
rect 44636 57034 44850 57068
rect 44250 57022 44850 57034
rect 44944 57068 45544 57080
rect 44944 57034 45158 57068
rect 45330 57034 45544 57068
rect 44944 57022 45544 57034
rect 46162 57068 46762 57080
rect 46162 57034 46376 57068
rect 46548 57034 46762 57068
rect 46162 57022 46762 57034
rect 46856 57068 47456 57080
rect 46856 57034 47070 57068
rect 47242 57034 47456 57068
rect 46856 57022 47456 57034
rect 47550 57068 48150 57080
rect 47550 57034 47764 57068
rect 47936 57034 48150 57068
rect 47550 57022 48150 57034
rect 48244 57068 48844 57080
rect 48244 57034 48458 57068
rect 48630 57034 48844 57068
rect 48244 57022 48844 57034
rect 48938 57068 49538 57080
rect 48938 57034 49152 57068
rect 49324 57034 49538 57068
rect 48938 57022 49538 57034
rect 50184 57068 50784 57080
rect 50184 57034 50398 57068
rect 50570 57034 50784 57068
rect 50184 57022 50784 57034
rect 50878 57068 51478 57080
rect 50878 57034 51092 57068
rect 51264 57034 51478 57068
rect 50878 57022 51478 57034
rect 51572 57068 52172 57080
rect 51572 57034 51786 57068
rect 51958 57034 52172 57068
rect 51572 57022 52172 57034
rect 52266 57068 52866 57080
rect 52266 57034 52480 57068
rect 52652 57034 52866 57068
rect 52266 57022 52866 57034
rect 52960 57068 53560 57080
rect 52960 57034 53174 57068
rect 53346 57034 53560 57068
rect 52960 57022 53560 57034
rect 54206 57068 54806 57080
rect 54206 57034 54420 57068
rect 54592 57034 54806 57068
rect 54206 57022 54806 57034
rect 54900 57068 55500 57080
rect 54900 57034 55114 57068
rect 55286 57034 55500 57068
rect 54900 57022 55500 57034
rect 55594 57068 56194 57080
rect 55594 57034 55808 57068
rect 55980 57034 56194 57068
rect 55594 57022 56194 57034
rect 56288 57068 56888 57080
rect 56288 57034 56502 57068
rect 56674 57034 56888 57068
rect 56288 57022 56888 57034
rect 56982 57068 57582 57080
rect 56982 57034 57196 57068
rect 57368 57034 57582 57068
rect 56982 57022 57582 57034
rect 42120 55968 42720 55980
rect 42120 55934 42334 55968
rect 42506 55934 42720 55968
rect 42120 55922 42720 55934
rect 42814 55968 43414 55980
rect 42814 55934 43028 55968
rect 43200 55934 43414 55968
rect 42814 55922 43414 55934
rect 43508 55968 44108 55980
rect 43508 55934 43722 55968
rect 43894 55934 44108 55968
rect 43508 55922 44108 55934
rect 44202 55968 44802 55980
rect 44202 55934 44416 55968
rect 44588 55934 44802 55968
rect 44202 55922 44802 55934
rect 44896 55968 45496 55980
rect 44896 55934 45110 55968
rect 45282 55934 45496 55968
rect 44896 55922 45496 55934
rect 46128 55966 46728 55978
rect 46128 55932 46342 55966
rect 46514 55932 46728 55966
rect 46128 55920 46728 55932
rect 46822 55966 47422 55978
rect 46822 55932 47036 55966
rect 47208 55932 47422 55966
rect 46822 55920 47422 55932
rect 47516 55966 48116 55978
rect 47516 55932 47730 55966
rect 47902 55932 48116 55966
rect 47516 55920 48116 55932
rect 48210 55966 48810 55978
rect 48210 55932 48424 55966
rect 48596 55932 48810 55966
rect 48210 55920 48810 55932
rect 48904 55966 49504 55978
rect 48904 55932 49118 55966
rect 49290 55932 49504 55966
rect 48904 55920 49504 55932
rect 50140 55966 50740 55978
rect 50140 55932 50354 55966
rect 50526 55932 50740 55966
rect 50140 55920 50740 55932
rect 50834 55966 51434 55978
rect 50834 55932 51048 55966
rect 51220 55932 51434 55966
rect 50834 55920 51434 55932
rect 51528 55966 52128 55978
rect 51528 55932 51742 55966
rect 51914 55932 52128 55966
rect 51528 55920 52128 55932
rect 52222 55966 52822 55978
rect 52222 55932 52436 55966
rect 52608 55932 52822 55966
rect 52222 55920 52822 55932
rect 52916 55966 53516 55978
rect 52916 55932 53130 55966
rect 53302 55932 53516 55966
rect 52916 55920 53516 55932
rect 54150 55966 54750 55978
rect 54150 55932 54364 55966
rect 54536 55932 54750 55966
rect 54150 55920 54750 55932
rect 54844 55966 55444 55978
rect 54844 55932 55058 55966
rect 55230 55932 55444 55966
rect 54844 55920 55444 55932
rect 55538 55966 56138 55978
rect 55538 55932 55752 55966
rect 55924 55932 56138 55966
rect 55538 55920 56138 55932
rect 56232 55966 56832 55978
rect 56232 55932 56446 55966
rect 56618 55932 56832 55966
rect 56232 55920 56832 55932
rect 56926 55966 57526 55978
rect 56926 55932 57140 55966
rect 57312 55932 57526 55966
rect 56926 55920 57526 55932
rect 42120 55310 42720 55322
rect 42120 55276 42334 55310
rect 42506 55276 42720 55310
rect 42120 55264 42720 55276
rect 42814 55310 43414 55322
rect 42814 55276 43028 55310
rect 43200 55276 43414 55310
rect 42814 55264 43414 55276
rect 43508 55310 44108 55322
rect 43508 55276 43722 55310
rect 43894 55276 44108 55310
rect 43508 55264 44108 55276
rect 44202 55310 44802 55322
rect 44202 55276 44416 55310
rect 44588 55276 44802 55310
rect 44202 55264 44802 55276
rect 44896 55310 45496 55322
rect 44896 55276 45110 55310
rect 45282 55276 45496 55310
rect 44896 55264 45496 55276
rect 46128 55308 46728 55320
rect 46128 55274 46342 55308
rect 46514 55274 46728 55308
rect 46128 55262 46728 55274
rect 46822 55308 47422 55320
rect 46822 55274 47036 55308
rect 47208 55274 47422 55308
rect 46822 55262 47422 55274
rect 47516 55308 48116 55320
rect 47516 55274 47730 55308
rect 47902 55274 48116 55308
rect 47516 55262 48116 55274
rect 48210 55308 48810 55320
rect 48210 55274 48424 55308
rect 48596 55274 48810 55308
rect 48210 55262 48810 55274
rect 48904 55308 49504 55320
rect 48904 55274 49118 55308
rect 49290 55274 49504 55308
rect 48904 55262 49504 55274
rect 50140 55308 50740 55320
rect 50140 55274 50354 55308
rect 50526 55274 50740 55308
rect 50140 55262 50740 55274
rect 50834 55308 51434 55320
rect 50834 55274 51048 55308
rect 51220 55274 51434 55308
rect 50834 55262 51434 55274
rect 51528 55308 52128 55320
rect 51528 55274 51742 55308
rect 51914 55274 52128 55308
rect 51528 55262 52128 55274
rect 52222 55308 52822 55320
rect 52222 55274 52436 55308
rect 52608 55274 52822 55308
rect 52222 55262 52822 55274
rect 52916 55308 53516 55320
rect 52916 55274 53130 55308
rect 53302 55274 53516 55308
rect 52916 55262 53516 55274
rect 54150 55308 54750 55320
rect 54150 55274 54364 55308
rect 54536 55274 54750 55308
rect 54150 55262 54750 55274
rect 54844 55308 55444 55320
rect 54844 55274 55058 55308
rect 55230 55274 55444 55308
rect 54844 55262 55444 55274
rect 55538 55308 56138 55320
rect 55538 55274 55752 55308
rect 55924 55274 56138 55308
rect 55538 55262 56138 55274
rect 56232 55308 56832 55320
rect 56232 55274 56446 55308
rect 56618 55274 56832 55308
rect 56232 55262 56832 55274
rect 56926 55308 57526 55320
rect 56926 55274 57140 55308
rect 57312 55274 57526 55308
rect 56926 55262 57526 55274
rect 42120 54652 42720 54664
rect 42120 54618 42334 54652
rect 42506 54618 42720 54652
rect 42120 54606 42720 54618
rect 42814 54652 43414 54664
rect 42814 54618 43028 54652
rect 43200 54618 43414 54652
rect 42814 54606 43414 54618
rect 43508 54652 44108 54664
rect 43508 54618 43722 54652
rect 43894 54618 44108 54652
rect 43508 54606 44108 54618
rect 44202 54652 44802 54664
rect 44202 54618 44416 54652
rect 44588 54618 44802 54652
rect 44202 54606 44802 54618
rect 44896 54652 45496 54664
rect 44896 54618 45110 54652
rect 45282 54618 45496 54652
rect 44896 54606 45496 54618
rect 46128 54650 46728 54662
rect 46128 54616 46342 54650
rect 46514 54616 46728 54650
rect 46128 54604 46728 54616
rect 46822 54650 47422 54662
rect 46822 54616 47036 54650
rect 47208 54616 47422 54650
rect 46822 54604 47422 54616
rect 47516 54650 48116 54662
rect 47516 54616 47730 54650
rect 47902 54616 48116 54650
rect 47516 54604 48116 54616
rect 48210 54650 48810 54662
rect 48210 54616 48424 54650
rect 48596 54616 48810 54650
rect 48210 54604 48810 54616
rect 48904 54650 49504 54662
rect 48904 54616 49118 54650
rect 49290 54616 49504 54650
rect 48904 54604 49504 54616
rect 50140 54650 50740 54662
rect 50140 54616 50354 54650
rect 50526 54616 50740 54650
rect 50140 54604 50740 54616
rect 50834 54650 51434 54662
rect 50834 54616 51048 54650
rect 51220 54616 51434 54650
rect 50834 54604 51434 54616
rect 51528 54650 52128 54662
rect 51528 54616 51742 54650
rect 51914 54616 52128 54650
rect 51528 54604 52128 54616
rect 52222 54650 52822 54662
rect 52222 54616 52436 54650
rect 52608 54616 52822 54650
rect 52222 54604 52822 54616
rect 52916 54650 53516 54662
rect 52916 54616 53130 54650
rect 53302 54616 53516 54650
rect 52916 54604 53516 54616
rect 54150 54650 54750 54662
rect 54150 54616 54364 54650
rect 54536 54616 54750 54650
rect 54150 54604 54750 54616
rect 54844 54650 55444 54662
rect 54844 54616 55058 54650
rect 55230 54616 55444 54650
rect 54844 54604 55444 54616
rect 55538 54650 56138 54662
rect 55538 54616 55752 54650
rect 55924 54616 56138 54650
rect 55538 54604 56138 54616
rect 56232 54650 56832 54662
rect 56232 54616 56446 54650
rect 56618 54616 56832 54650
rect 56232 54604 56832 54616
rect 56926 54650 57526 54662
rect 56926 54616 57140 54650
rect 57312 54616 57526 54650
rect 56926 54604 57526 54616
rect 42120 53994 42720 54006
rect 42120 53960 42334 53994
rect 42506 53960 42720 53994
rect 42120 53948 42720 53960
rect 42814 53994 43414 54006
rect 42814 53960 43028 53994
rect 43200 53960 43414 53994
rect 42814 53948 43414 53960
rect 43508 53994 44108 54006
rect 43508 53960 43722 53994
rect 43894 53960 44108 53994
rect 43508 53948 44108 53960
rect 44202 53994 44802 54006
rect 44202 53960 44416 53994
rect 44588 53960 44802 53994
rect 44202 53948 44802 53960
rect 44896 53994 45496 54006
rect 44896 53960 45110 53994
rect 45282 53960 45496 53994
rect 44896 53948 45496 53960
rect 46128 53992 46728 54004
rect 46128 53958 46342 53992
rect 46514 53958 46728 53992
rect 46128 53946 46728 53958
rect 46822 53992 47422 54004
rect 46822 53958 47036 53992
rect 47208 53958 47422 53992
rect 46822 53946 47422 53958
rect 47516 53992 48116 54004
rect 47516 53958 47730 53992
rect 47902 53958 48116 53992
rect 47516 53946 48116 53958
rect 48210 53992 48810 54004
rect 48210 53958 48424 53992
rect 48596 53958 48810 53992
rect 48210 53946 48810 53958
rect 48904 53992 49504 54004
rect 48904 53958 49118 53992
rect 49290 53958 49504 53992
rect 48904 53946 49504 53958
rect 50140 53992 50740 54004
rect 50140 53958 50354 53992
rect 50526 53958 50740 53992
rect 50140 53946 50740 53958
rect 50834 53992 51434 54004
rect 50834 53958 51048 53992
rect 51220 53958 51434 53992
rect 50834 53946 51434 53958
rect 51528 53992 52128 54004
rect 51528 53958 51742 53992
rect 51914 53958 52128 53992
rect 51528 53946 52128 53958
rect 52222 53992 52822 54004
rect 52222 53958 52436 53992
rect 52608 53958 52822 53992
rect 52222 53946 52822 53958
rect 52916 53992 53516 54004
rect 52916 53958 53130 53992
rect 53302 53958 53516 53992
rect 52916 53946 53516 53958
rect 54150 53992 54750 54004
rect 54150 53958 54364 53992
rect 54536 53958 54750 53992
rect 54150 53946 54750 53958
rect 54844 53992 55444 54004
rect 54844 53958 55058 53992
rect 55230 53958 55444 53992
rect 54844 53946 55444 53958
rect 55538 53992 56138 54004
rect 55538 53958 55752 53992
rect 55924 53958 56138 53992
rect 55538 53946 56138 53958
rect 56232 53992 56832 54004
rect 56232 53958 56446 53992
rect 56618 53958 56832 53992
rect 56232 53946 56832 53958
rect 56926 53992 57526 54004
rect 56926 53958 57140 53992
rect 57312 53958 57526 53992
rect 56926 53946 57526 53958
rect 42120 53336 42720 53348
rect 42120 53302 42334 53336
rect 42506 53302 42720 53336
rect 42120 53290 42720 53302
rect 42814 53336 43414 53348
rect 42814 53302 43028 53336
rect 43200 53302 43414 53336
rect 42814 53290 43414 53302
rect 43508 53336 44108 53348
rect 43508 53302 43722 53336
rect 43894 53302 44108 53336
rect 43508 53290 44108 53302
rect 44202 53336 44802 53348
rect 44202 53302 44416 53336
rect 44588 53302 44802 53336
rect 44202 53290 44802 53302
rect 44896 53336 45496 53348
rect 44896 53302 45110 53336
rect 45282 53302 45496 53336
rect 44896 53290 45496 53302
rect 71294 58040 71352 58254
rect 71294 57868 71306 58040
rect 71340 57868 71352 58040
rect 71294 57654 71352 57868
rect 71952 58040 72010 58254
rect 71952 57868 71964 58040
rect 71998 57868 72010 58040
rect 71952 57654 72010 57868
rect 72610 58040 72668 58254
rect 72610 57868 72622 58040
rect 72656 57868 72668 58040
rect 72610 57654 72668 57868
rect 73268 58040 73326 58254
rect 73268 57868 73280 58040
rect 73314 57868 73326 58040
rect 73268 57654 73326 57868
rect 73926 58040 73984 58254
rect 73926 57868 73938 58040
rect 73972 57868 73984 58040
rect 75158 58020 75216 58234
rect 73926 57654 73984 57868
rect 71294 57346 71352 57560
rect 71294 57174 71306 57346
rect 71340 57174 71352 57346
rect 71294 56960 71352 57174
rect 71952 57346 72010 57560
rect 71952 57174 71964 57346
rect 71998 57174 72010 57346
rect 71952 56960 72010 57174
rect 72610 57346 72668 57560
rect 72610 57174 72622 57346
rect 72656 57174 72668 57346
rect 72610 56960 72668 57174
rect 73268 57346 73326 57560
rect 73268 57174 73280 57346
rect 73314 57174 73326 57346
rect 73268 56960 73326 57174
rect 73926 57346 73984 57560
rect 73926 57174 73938 57346
rect 73972 57174 73984 57346
rect 73926 56960 73984 57174
rect 71294 56652 71352 56866
rect 71294 56480 71306 56652
rect 71340 56480 71352 56652
rect 71294 56266 71352 56480
rect 71952 56652 72010 56866
rect 71952 56480 71964 56652
rect 71998 56480 72010 56652
rect 71952 56266 72010 56480
rect 72610 56652 72668 56866
rect 72610 56480 72622 56652
rect 72656 56480 72668 56652
rect 72610 56266 72668 56480
rect 73268 56652 73326 56866
rect 73268 56480 73280 56652
rect 73314 56480 73326 56652
rect 73268 56266 73326 56480
rect 73926 56652 73984 56866
rect 73926 56480 73938 56652
rect 73972 56480 73984 56652
rect 73926 56266 73984 56480
rect 71294 55958 71352 56172
rect 71294 55786 71306 55958
rect 71340 55786 71352 55958
rect 71294 55572 71352 55786
rect 71952 55958 72010 56172
rect 71952 55786 71964 55958
rect 71998 55786 72010 55958
rect 71952 55572 72010 55786
rect 72610 55958 72668 56172
rect 72610 55786 72622 55958
rect 72656 55786 72668 55958
rect 72610 55572 72668 55786
rect 73268 55958 73326 56172
rect 73268 55786 73280 55958
rect 73314 55786 73326 55958
rect 73268 55572 73326 55786
rect 73926 55958 73984 56172
rect 73926 55786 73938 55958
rect 73972 55786 73984 55958
rect 73926 55572 73984 55786
rect 71294 55264 71352 55478
rect 71294 55092 71306 55264
rect 71340 55092 71352 55264
rect 71294 54878 71352 55092
rect 71952 55264 72010 55478
rect 71952 55092 71964 55264
rect 71998 55092 72010 55264
rect 71952 54878 72010 55092
rect 72610 55264 72668 55478
rect 72610 55092 72622 55264
rect 72656 55092 72668 55264
rect 72610 54878 72668 55092
rect 73268 55264 73326 55478
rect 73268 55092 73280 55264
rect 73314 55092 73326 55264
rect 73268 54878 73326 55092
rect 73926 55264 73984 55478
rect 73926 55092 73938 55264
rect 73972 55092 73984 55264
rect 75158 57848 75170 58020
rect 75204 57848 75216 58020
rect 75158 57634 75216 57848
rect 75816 58020 75874 58234
rect 75816 57848 75828 58020
rect 75862 57848 75874 58020
rect 75816 57634 75874 57848
rect 76474 58020 76532 58234
rect 76474 57848 76486 58020
rect 76520 57848 76532 58020
rect 76474 57634 76532 57848
rect 77132 58020 77190 58234
rect 77132 57848 77144 58020
rect 77178 57848 77190 58020
rect 77132 57634 77190 57848
rect 77790 58020 77848 58234
rect 79008 58034 79066 58248
rect 77790 57848 77802 58020
rect 77836 57848 77848 58020
rect 77790 57634 77848 57848
rect 75158 57326 75216 57540
rect 75158 57154 75170 57326
rect 75204 57154 75216 57326
rect 75158 56940 75216 57154
rect 75816 57326 75874 57540
rect 75816 57154 75828 57326
rect 75862 57154 75874 57326
rect 75816 56940 75874 57154
rect 76474 57326 76532 57540
rect 76474 57154 76486 57326
rect 76520 57154 76532 57326
rect 76474 56940 76532 57154
rect 77132 57326 77190 57540
rect 77132 57154 77144 57326
rect 77178 57154 77190 57326
rect 77132 56940 77190 57154
rect 77790 57326 77848 57540
rect 77790 57154 77802 57326
rect 77836 57154 77848 57326
rect 77790 56940 77848 57154
rect 75158 56632 75216 56846
rect 75158 56460 75170 56632
rect 75204 56460 75216 56632
rect 75158 56246 75216 56460
rect 75816 56632 75874 56846
rect 75816 56460 75828 56632
rect 75862 56460 75874 56632
rect 75816 56246 75874 56460
rect 76474 56632 76532 56846
rect 76474 56460 76486 56632
rect 76520 56460 76532 56632
rect 76474 56246 76532 56460
rect 77132 56632 77190 56846
rect 77132 56460 77144 56632
rect 77178 56460 77190 56632
rect 77132 56246 77190 56460
rect 77790 56632 77848 56846
rect 77790 56460 77802 56632
rect 77836 56460 77848 56632
rect 77790 56246 77848 56460
rect 75158 55938 75216 56152
rect 75158 55766 75170 55938
rect 75204 55766 75216 55938
rect 75158 55552 75216 55766
rect 75816 55938 75874 56152
rect 75816 55766 75828 55938
rect 75862 55766 75874 55938
rect 75816 55552 75874 55766
rect 76474 55938 76532 56152
rect 76474 55766 76486 55938
rect 76520 55766 76532 55938
rect 76474 55552 76532 55766
rect 77132 55938 77190 56152
rect 77132 55766 77144 55938
rect 77178 55766 77190 55938
rect 77132 55552 77190 55766
rect 77790 55938 77848 56152
rect 77790 55766 77802 55938
rect 77836 55766 77848 55938
rect 77790 55552 77848 55766
rect 75158 55244 75216 55458
rect 73926 54878 73984 55092
rect 75158 55072 75170 55244
rect 75204 55072 75216 55244
rect 75158 54858 75216 55072
rect 75816 55244 75874 55458
rect 75816 55072 75828 55244
rect 75862 55072 75874 55244
rect 75816 54858 75874 55072
rect 76474 55244 76532 55458
rect 76474 55072 76486 55244
rect 76520 55072 76532 55244
rect 76474 54858 76532 55072
rect 77132 55244 77190 55458
rect 77132 55072 77144 55244
rect 77178 55072 77190 55244
rect 77132 54858 77190 55072
rect 77790 55244 77848 55458
rect 77790 55072 77802 55244
rect 77836 55072 77848 55244
rect 79008 57862 79020 58034
rect 79054 57862 79066 58034
rect 79008 57648 79066 57862
rect 79666 58034 79724 58248
rect 79666 57862 79678 58034
rect 79712 57862 79724 58034
rect 79666 57648 79724 57862
rect 80324 58034 80382 58248
rect 80324 57862 80336 58034
rect 80370 57862 80382 58034
rect 80324 57648 80382 57862
rect 80982 58034 81040 58248
rect 80982 57862 80994 58034
rect 81028 57862 81040 58034
rect 80982 57648 81040 57862
rect 81640 58034 81698 58248
rect 81640 57862 81652 58034
rect 81686 57862 81698 58034
rect 81640 57648 81698 57862
rect 79008 57340 79066 57554
rect 79008 57168 79020 57340
rect 79054 57168 79066 57340
rect 79008 56954 79066 57168
rect 79666 57340 79724 57554
rect 79666 57168 79678 57340
rect 79712 57168 79724 57340
rect 79666 56954 79724 57168
rect 80324 57340 80382 57554
rect 80324 57168 80336 57340
rect 80370 57168 80382 57340
rect 80324 56954 80382 57168
rect 80982 57340 81040 57554
rect 80982 57168 80994 57340
rect 81028 57168 81040 57340
rect 80982 56954 81040 57168
rect 81640 57340 81698 57554
rect 81640 57168 81652 57340
rect 81686 57168 81698 57340
rect 81640 56954 81698 57168
rect 79008 56646 79066 56860
rect 79008 56474 79020 56646
rect 79054 56474 79066 56646
rect 79008 56260 79066 56474
rect 79666 56646 79724 56860
rect 79666 56474 79678 56646
rect 79712 56474 79724 56646
rect 79666 56260 79724 56474
rect 80324 56646 80382 56860
rect 80324 56474 80336 56646
rect 80370 56474 80382 56646
rect 80324 56260 80382 56474
rect 80982 56646 81040 56860
rect 80982 56474 80994 56646
rect 81028 56474 81040 56646
rect 80982 56260 81040 56474
rect 81640 56646 81698 56860
rect 81640 56474 81652 56646
rect 81686 56474 81698 56646
rect 81640 56260 81698 56474
rect 79008 55952 79066 56166
rect 79008 55780 79020 55952
rect 79054 55780 79066 55952
rect 79008 55566 79066 55780
rect 79666 55952 79724 56166
rect 79666 55780 79678 55952
rect 79712 55780 79724 55952
rect 79666 55566 79724 55780
rect 80324 55952 80382 56166
rect 80324 55780 80336 55952
rect 80370 55780 80382 55952
rect 80324 55566 80382 55780
rect 80982 55952 81040 56166
rect 80982 55780 80994 55952
rect 81028 55780 81040 55952
rect 80982 55566 81040 55780
rect 81640 55952 81698 56166
rect 81640 55780 81652 55952
rect 81686 55780 81698 55952
rect 81640 55566 81698 55780
rect 79008 55258 79066 55472
rect 77790 54858 77848 55072
rect 79008 55086 79020 55258
rect 79054 55086 79066 55258
rect 79008 54872 79066 55086
rect 79666 55258 79724 55472
rect 79666 55086 79678 55258
rect 79712 55086 79724 55258
rect 79666 54872 79724 55086
rect 80324 55258 80382 55472
rect 80324 55086 80336 55258
rect 80370 55086 80382 55258
rect 80324 54872 80382 55086
rect 80982 55258 81040 55472
rect 80982 55086 80994 55258
rect 81028 55086 81040 55258
rect 80982 54872 81040 55086
rect 81640 55258 81698 55472
rect 81640 55086 81652 55258
rect 81686 55086 81698 55258
rect 81640 54872 81698 55086
rect 46128 53334 46728 53346
rect 46128 53300 46342 53334
rect 46514 53300 46728 53334
rect 46128 53288 46728 53300
rect 46822 53334 47422 53346
rect 46822 53300 47036 53334
rect 47208 53300 47422 53334
rect 46822 53288 47422 53300
rect 47516 53334 48116 53346
rect 47516 53300 47730 53334
rect 47902 53300 48116 53334
rect 47516 53288 48116 53300
rect 48210 53334 48810 53346
rect 48210 53300 48424 53334
rect 48596 53300 48810 53334
rect 48210 53288 48810 53300
rect 48904 53334 49504 53346
rect 48904 53300 49118 53334
rect 49290 53300 49504 53334
rect 48904 53288 49504 53300
rect 50140 53334 50740 53346
rect 50140 53300 50354 53334
rect 50526 53300 50740 53334
rect 50140 53288 50740 53300
rect 50834 53334 51434 53346
rect 50834 53300 51048 53334
rect 51220 53300 51434 53334
rect 50834 53288 51434 53300
rect 51528 53334 52128 53346
rect 51528 53300 51742 53334
rect 51914 53300 52128 53334
rect 51528 53288 52128 53300
rect 52222 53334 52822 53346
rect 52222 53300 52436 53334
rect 52608 53300 52822 53334
rect 52222 53288 52822 53300
rect 52916 53334 53516 53346
rect 52916 53300 53130 53334
rect 53302 53300 53516 53334
rect 52916 53288 53516 53300
rect 54150 53334 54750 53346
rect 54150 53300 54364 53334
rect 54536 53300 54750 53334
rect 54150 53288 54750 53300
rect 54844 53334 55444 53346
rect 54844 53300 55058 53334
rect 55230 53300 55444 53334
rect 54844 53288 55444 53300
rect 55538 53334 56138 53346
rect 55538 53300 55752 53334
rect 55924 53300 56138 53334
rect 55538 53288 56138 53300
rect 56232 53334 56832 53346
rect 56232 53300 56446 53334
rect 56618 53300 56832 53334
rect 56232 53288 56832 53300
rect 56926 53334 57526 53346
rect 56926 53300 57140 53334
rect 57312 53300 57526 53334
rect 56926 53288 57526 53300
rect 42120 52678 42720 52690
rect 42120 52644 42334 52678
rect 42506 52644 42720 52678
rect 42120 52632 42720 52644
rect 42814 52678 43414 52690
rect 42814 52644 43028 52678
rect 43200 52644 43414 52678
rect 42814 52632 43414 52644
rect 43508 52678 44108 52690
rect 43508 52644 43722 52678
rect 43894 52644 44108 52678
rect 43508 52632 44108 52644
rect 44202 52678 44802 52690
rect 44202 52644 44416 52678
rect 44588 52644 44802 52678
rect 44202 52632 44802 52644
rect 44896 52678 45496 52690
rect 44896 52644 45110 52678
rect 45282 52644 45496 52678
rect 44896 52632 45496 52644
rect 46128 52676 46728 52688
rect 46128 52642 46342 52676
rect 46514 52642 46728 52676
rect 46128 52630 46728 52642
rect 46822 52676 47422 52688
rect 46822 52642 47036 52676
rect 47208 52642 47422 52676
rect 46822 52630 47422 52642
rect 47516 52676 48116 52688
rect 47516 52642 47730 52676
rect 47902 52642 48116 52676
rect 47516 52630 48116 52642
rect 48210 52676 48810 52688
rect 48210 52642 48424 52676
rect 48596 52642 48810 52676
rect 48210 52630 48810 52642
rect 48904 52676 49504 52688
rect 48904 52642 49118 52676
rect 49290 52642 49504 52676
rect 48904 52630 49504 52642
rect 50140 52676 50740 52688
rect 50140 52642 50354 52676
rect 50526 52642 50740 52676
rect 50140 52630 50740 52642
rect 50834 52676 51434 52688
rect 50834 52642 51048 52676
rect 51220 52642 51434 52676
rect 50834 52630 51434 52642
rect 51528 52676 52128 52688
rect 51528 52642 51742 52676
rect 51914 52642 52128 52676
rect 51528 52630 52128 52642
rect 52222 52676 52822 52688
rect 52222 52642 52436 52676
rect 52608 52642 52822 52676
rect 52222 52630 52822 52642
rect 52916 52676 53516 52688
rect 52916 52642 53130 52676
rect 53302 52642 53516 52676
rect 52916 52630 53516 52642
rect 54150 52676 54750 52688
rect 54150 52642 54364 52676
rect 54536 52642 54750 52676
rect 54150 52630 54750 52642
rect 54844 52676 55444 52688
rect 54844 52642 55058 52676
rect 55230 52642 55444 52676
rect 54844 52630 55444 52642
rect 55538 52676 56138 52688
rect 55538 52642 55752 52676
rect 55924 52642 56138 52676
rect 55538 52630 56138 52642
rect 56232 52676 56832 52688
rect 56232 52642 56446 52676
rect 56618 52642 56832 52676
rect 56232 52630 56832 52642
rect 56926 52676 57526 52688
rect 56926 52642 57140 52676
rect 57312 52642 57526 52676
rect 56926 52630 57526 52642
rect 42112 51770 42712 51782
rect 42112 51736 42326 51770
rect 42498 51736 42712 51770
rect 42112 51724 42712 51736
rect 42806 51770 43406 51782
rect 42806 51736 43020 51770
rect 43192 51736 43406 51770
rect 42806 51724 43406 51736
rect 43500 51770 44100 51782
rect 43500 51736 43714 51770
rect 43886 51736 44100 51770
rect 43500 51724 44100 51736
rect 44194 51770 44794 51782
rect 44194 51736 44408 51770
rect 44580 51736 44794 51770
rect 44194 51724 44794 51736
rect 44888 51770 45488 51782
rect 44888 51736 45102 51770
rect 45274 51736 45488 51770
rect 44888 51724 45488 51736
rect 46106 51770 46706 51782
rect 46106 51736 46320 51770
rect 46492 51736 46706 51770
rect 46106 51724 46706 51736
rect 46800 51770 47400 51782
rect 46800 51736 47014 51770
rect 47186 51736 47400 51770
rect 46800 51724 47400 51736
rect 47494 51770 48094 51782
rect 47494 51736 47708 51770
rect 47880 51736 48094 51770
rect 47494 51724 48094 51736
rect 48188 51770 48788 51782
rect 48188 51736 48402 51770
rect 48574 51736 48788 51770
rect 48188 51724 48788 51736
rect 48882 51770 49482 51782
rect 48882 51736 49096 51770
rect 49268 51736 49482 51770
rect 48882 51724 49482 51736
rect 50128 51770 50728 51782
rect 50128 51736 50342 51770
rect 50514 51736 50728 51770
rect 50128 51724 50728 51736
rect 50822 51770 51422 51782
rect 50822 51736 51036 51770
rect 51208 51736 51422 51770
rect 50822 51724 51422 51736
rect 51516 51770 52116 51782
rect 51516 51736 51730 51770
rect 51902 51736 52116 51770
rect 51516 51724 52116 51736
rect 52210 51770 52810 51782
rect 52210 51736 52424 51770
rect 52596 51736 52810 51770
rect 52210 51724 52810 51736
rect 52904 51770 53504 51782
rect 52904 51736 53118 51770
rect 53290 51736 53504 51770
rect 52904 51724 53504 51736
rect 54150 51770 54750 51782
rect 54150 51736 54364 51770
rect 54536 51736 54750 51770
rect 54150 51724 54750 51736
rect 54844 51770 55444 51782
rect 54844 51736 55058 51770
rect 55230 51736 55444 51770
rect 54844 51724 55444 51736
rect 55538 51770 56138 51782
rect 55538 51736 55752 51770
rect 55924 51736 56138 51770
rect 55538 51724 56138 51736
rect 56232 51770 56832 51782
rect 56232 51736 56446 51770
rect 56618 51736 56832 51770
rect 56232 51724 56832 51736
rect 56926 51770 57526 51782
rect 56926 51736 57140 51770
rect 57312 51736 57526 51770
rect 56926 51724 57526 51736
rect 71298 54268 71356 54482
rect 71298 54096 71310 54268
rect 71344 54096 71356 54268
rect 71298 53882 71356 54096
rect 71956 54268 72014 54482
rect 71956 54096 71968 54268
rect 72002 54096 72014 54268
rect 71956 53882 72014 54096
rect 72614 54268 72672 54482
rect 72614 54096 72626 54268
rect 72660 54096 72672 54268
rect 72614 53882 72672 54096
rect 73272 54268 73330 54482
rect 73272 54096 73284 54268
rect 73318 54096 73330 54268
rect 73272 53882 73330 54096
rect 73930 54268 73988 54482
rect 73930 54096 73942 54268
rect 73976 54096 73988 54268
rect 75162 54248 75220 54462
rect 73930 53882 73988 54096
rect 71298 53574 71356 53788
rect 71298 53402 71310 53574
rect 71344 53402 71356 53574
rect 71298 53188 71356 53402
rect 71956 53574 72014 53788
rect 71956 53402 71968 53574
rect 72002 53402 72014 53574
rect 71956 53188 72014 53402
rect 72614 53574 72672 53788
rect 72614 53402 72626 53574
rect 72660 53402 72672 53574
rect 72614 53188 72672 53402
rect 73272 53574 73330 53788
rect 73272 53402 73284 53574
rect 73318 53402 73330 53574
rect 73272 53188 73330 53402
rect 73930 53574 73988 53788
rect 73930 53402 73942 53574
rect 73976 53402 73988 53574
rect 73930 53188 73988 53402
rect 71298 52880 71356 53094
rect 71298 52708 71310 52880
rect 71344 52708 71356 52880
rect 71298 52494 71356 52708
rect 71956 52880 72014 53094
rect 71956 52708 71968 52880
rect 72002 52708 72014 52880
rect 71956 52494 72014 52708
rect 72614 52880 72672 53094
rect 72614 52708 72626 52880
rect 72660 52708 72672 52880
rect 72614 52494 72672 52708
rect 73272 52880 73330 53094
rect 73272 52708 73284 52880
rect 73318 52708 73330 52880
rect 73272 52494 73330 52708
rect 73930 52880 73988 53094
rect 73930 52708 73942 52880
rect 73976 52708 73988 52880
rect 73930 52494 73988 52708
rect 71298 52186 71356 52400
rect 71298 52014 71310 52186
rect 71344 52014 71356 52186
rect 71298 51800 71356 52014
rect 71956 52186 72014 52400
rect 71956 52014 71968 52186
rect 72002 52014 72014 52186
rect 71956 51800 72014 52014
rect 72614 52186 72672 52400
rect 72614 52014 72626 52186
rect 72660 52014 72672 52186
rect 72614 51800 72672 52014
rect 73272 52186 73330 52400
rect 73272 52014 73284 52186
rect 73318 52014 73330 52186
rect 73272 51800 73330 52014
rect 73930 52186 73988 52400
rect 73930 52014 73942 52186
rect 73976 52014 73988 52186
rect 73930 51800 73988 52014
rect 42112 51112 42712 51124
rect 42112 51078 42326 51112
rect 42498 51078 42712 51112
rect 42112 51066 42712 51078
rect 42806 51112 43406 51124
rect 42806 51078 43020 51112
rect 43192 51078 43406 51112
rect 42806 51066 43406 51078
rect 43500 51112 44100 51124
rect 43500 51078 43714 51112
rect 43886 51078 44100 51112
rect 43500 51066 44100 51078
rect 44194 51112 44794 51124
rect 44194 51078 44408 51112
rect 44580 51078 44794 51112
rect 44194 51066 44794 51078
rect 44888 51112 45488 51124
rect 44888 51078 45102 51112
rect 45274 51078 45488 51112
rect 44888 51066 45488 51078
rect 46106 51112 46706 51124
rect 46106 51078 46320 51112
rect 46492 51078 46706 51112
rect 46106 51066 46706 51078
rect 46800 51112 47400 51124
rect 46800 51078 47014 51112
rect 47186 51078 47400 51112
rect 46800 51066 47400 51078
rect 47494 51112 48094 51124
rect 47494 51078 47708 51112
rect 47880 51078 48094 51112
rect 47494 51066 48094 51078
rect 48188 51112 48788 51124
rect 48188 51078 48402 51112
rect 48574 51078 48788 51112
rect 48188 51066 48788 51078
rect 48882 51112 49482 51124
rect 48882 51078 49096 51112
rect 49268 51078 49482 51112
rect 48882 51066 49482 51078
rect 50128 51112 50728 51124
rect 50128 51078 50342 51112
rect 50514 51078 50728 51112
rect 50128 51066 50728 51078
rect 50822 51112 51422 51124
rect 50822 51078 51036 51112
rect 51208 51078 51422 51112
rect 50822 51066 51422 51078
rect 51516 51112 52116 51124
rect 51516 51078 51730 51112
rect 51902 51078 52116 51112
rect 51516 51066 52116 51078
rect 52210 51112 52810 51124
rect 52210 51078 52424 51112
rect 52596 51078 52810 51112
rect 52210 51066 52810 51078
rect 52904 51112 53504 51124
rect 52904 51078 53118 51112
rect 53290 51078 53504 51112
rect 52904 51066 53504 51078
rect 54150 51112 54750 51124
rect 54150 51078 54364 51112
rect 54536 51078 54750 51112
rect 54150 51066 54750 51078
rect 54844 51112 55444 51124
rect 54844 51078 55058 51112
rect 55230 51078 55444 51112
rect 54844 51066 55444 51078
rect 55538 51112 56138 51124
rect 55538 51078 55752 51112
rect 55924 51078 56138 51112
rect 55538 51066 56138 51078
rect 56232 51112 56832 51124
rect 56232 51078 56446 51112
rect 56618 51078 56832 51112
rect 56232 51066 56832 51078
rect 56926 51112 57526 51124
rect 56926 51078 57140 51112
rect 57312 51078 57526 51112
rect 56926 51066 57526 51078
rect 71298 51492 71356 51706
rect 71298 51320 71310 51492
rect 71344 51320 71356 51492
rect 71298 51106 71356 51320
rect 71956 51492 72014 51706
rect 71956 51320 71968 51492
rect 72002 51320 72014 51492
rect 71956 51106 72014 51320
rect 72614 51492 72672 51706
rect 72614 51320 72626 51492
rect 72660 51320 72672 51492
rect 72614 51106 72672 51320
rect 73272 51492 73330 51706
rect 73272 51320 73284 51492
rect 73318 51320 73330 51492
rect 73272 51106 73330 51320
rect 73930 51492 73988 51706
rect 73930 51320 73942 51492
rect 73976 51320 73988 51492
rect 75162 54076 75174 54248
rect 75208 54076 75220 54248
rect 75162 53862 75220 54076
rect 75820 54248 75878 54462
rect 75820 54076 75832 54248
rect 75866 54076 75878 54248
rect 75820 53862 75878 54076
rect 76478 54248 76536 54462
rect 76478 54076 76490 54248
rect 76524 54076 76536 54248
rect 76478 53862 76536 54076
rect 77136 54248 77194 54462
rect 77136 54076 77148 54248
rect 77182 54076 77194 54248
rect 77136 53862 77194 54076
rect 77794 54248 77852 54462
rect 79012 54262 79070 54476
rect 77794 54076 77806 54248
rect 77840 54076 77852 54248
rect 77794 53862 77852 54076
rect 75162 53554 75220 53768
rect 75162 53382 75174 53554
rect 75208 53382 75220 53554
rect 75162 53168 75220 53382
rect 75820 53554 75878 53768
rect 75820 53382 75832 53554
rect 75866 53382 75878 53554
rect 75820 53168 75878 53382
rect 76478 53554 76536 53768
rect 76478 53382 76490 53554
rect 76524 53382 76536 53554
rect 76478 53168 76536 53382
rect 77136 53554 77194 53768
rect 77136 53382 77148 53554
rect 77182 53382 77194 53554
rect 77136 53168 77194 53382
rect 77794 53554 77852 53768
rect 77794 53382 77806 53554
rect 77840 53382 77852 53554
rect 77794 53168 77852 53382
rect 75162 52860 75220 53074
rect 75162 52688 75174 52860
rect 75208 52688 75220 52860
rect 75162 52474 75220 52688
rect 75820 52860 75878 53074
rect 75820 52688 75832 52860
rect 75866 52688 75878 52860
rect 75820 52474 75878 52688
rect 76478 52860 76536 53074
rect 76478 52688 76490 52860
rect 76524 52688 76536 52860
rect 76478 52474 76536 52688
rect 77136 52860 77194 53074
rect 77136 52688 77148 52860
rect 77182 52688 77194 52860
rect 77136 52474 77194 52688
rect 77794 52860 77852 53074
rect 77794 52688 77806 52860
rect 77840 52688 77852 52860
rect 77794 52474 77852 52688
rect 75162 52166 75220 52380
rect 75162 51994 75174 52166
rect 75208 51994 75220 52166
rect 75162 51780 75220 51994
rect 75820 52166 75878 52380
rect 75820 51994 75832 52166
rect 75866 51994 75878 52166
rect 75820 51780 75878 51994
rect 76478 52166 76536 52380
rect 76478 51994 76490 52166
rect 76524 51994 76536 52166
rect 76478 51780 76536 51994
rect 77136 52166 77194 52380
rect 77136 51994 77148 52166
rect 77182 51994 77194 52166
rect 77136 51780 77194 51994
rect 77794 52166 77852 52380
rect 77794 51994 77806 52166
rect 77840 51994 77852 52166
rect 77794 51780 77852 51994
rect 75162 51472 75220 51686
rect 73930 51106 73988 51320
rect 75162 51300 75174 51472
rect 75208 51300 75220 51472
rect 75162 51086 75220 51300
rect 75820 51472 75878 51686
rect 75820 51300 75832 51472
rect 75866 51300 75878 51472
rect 75820 51086 75878 51300
rect 76478 51472 76536 51686
rect 76478 51300 76490 51472
rect 76524 51300 76536 51472
rect 76478 51086 76536 51300
rect 77136 51472 77194 51686
rect 77136 51300 77148 51472
rect 77182 51300 77194 51472
rect 77136 51086 77194 51300
rect 77794 51472 77852 51686
rect 77794 51300 77806 51472
rect 77840 51300 77852 51472
rect 79012 54090 79024 54262
rect 79058 54090 79070 54262
rect 79012 53876 79070 54090
rect 79670 54262 79728 54476
rect 79670 54090 79682 54262
rect 79716 54090 79728 54262
rect 79670 53876 79728 54090
rect 80328 54262 80386 54476
rect 80328 54090 80340 54262
rect 80374 54090 80386 54262
rect 80328 53876 80386 54090
rect 80986 54262 81044 54476
rect 80986 54090 80998 54262
rect 81032 54090 81044 54262
rect 80986 53876 81044 54090
rect 81644 54262 81702 54476
rect 81644 54090 81656 54262
rect 81690 54090 81702 54262
rect 81644 53876 81702 54090
rect 79012 53568 79070 53782
rect 79012 53396 79024 53568
rect 79058 53396 79070 53568
rect 79012 53182 79070 53396
rect 79670 53568 79728 53782
rect 79670 53396 79682 53568
rect 79716 53396 79728 53568
rect 79670 53182 79728 53396
rect 80328 53568 80386 53782
rect 80328 53396 80340 53568
rect 80374 53396 80386 53568
rect 80328 53182 80386 53396
rect 80986 53568 81044 53782
rect 80986 53396 80998 53568
rect 81032 53396 81044 53568
rect 80986 53182 81044 53396
rect 81644 53568 81702 53782
rect 81644 53396 81656 53568
rect 81690 53396 81702 53568
rect 81644 53182 81702 53396
rect 79012 52874 79070 53088
rect 79012 52702 79024 52874
rect 79058 52702 79070 52874
rect 79012 52488 79070 52702
rect 79670 52874 79728 53088
rect 79670 52702 79682 52874
rect 79716 52702 79728 52874
rect 79670 52488 79728 52702
rect 80328 52874 80386 53088
rect 80328 52702 80340 52874
rect 80374 52702 80386 52874
rect 80328 52488 80386 52702
rect 80986 52874 81044 53088
rect 80986 52702 80998 52874
rect 81032 52702 81044 52874
rect 80986 52488 81044 52702
rect 81644 52874 81702 53088
rect 81644 52702 81656 52874
rect 81690 52702 81702 52874
rect 81644 52488 81702 52702
rect 79012 52180 79070 52394
rect 79012 52008 79024 52180
rect 79058 52008 79070 52180
rect 79012 51794 79070 52008
rect 79670 52180 79728 52394
rect 79670 52008 79682 52180
rect 79716 52008 79728 52180
rect 79670 51794 79728 52008
rect 80328 52180 80386 52394
rect 80328 52008 80340 52180
rect 80374 52008 80386 52180
rect 80328 51794 80386 52008
rect 80986 52180 81044 52394
rect 80986 52008 80998 52180
rect 81032 52008 81044 52180
rect 80986 51794 81044 52008
rect 81644 52180 81702 52394
rect 81644 52008 81656 52180
rect 81690 52008 81702 52180
rect 81644 51794 81702 52008
rect 79012 51486 79070 51700
rect 77794 51086 77852 51300
rect 79012 51314 79024 51486
rect 79058 51314 79070 51486
rect 79012 51100 79070 51314
rect 79670 51486 79728 51700
rect 79670 51314 79682 51486
rect 79716 51314 79728 51486
rect 79670 51100 79728 51314
rect 80328 51486 80386 51700
rect 80328 51314 80340 51486
rect 80374 51314 80386 51486
rect 80328 51100 80386 51314
rect 80986 51486 81044 51700
rect 80986 51314 80998 51486
rect 81032 51314 81044 51486
rect 80986 51100 81044 51314
rect 81644 51486 81702 51700
rect 81644 51314 81656 51486
rect 81690 51314 81702 51486
rect 81644 51100 81702 51314
rect 84834 53998 84891 54011
rect 83302 53943 83355 53955
rect 83302 53909 83310 53943
rect 83344 53909 83355 53943
rect 83302 53851 83355 53909
rect 83302 53817 83310 53851
rect 83344 53817 83355 53851
rect 83302 53805 83355 53817
rect 83455 53947 83511 53955
rect 83455 53913 83466 53947
rect 83500 53913 83511 53947
rect 83455 53847 83511 53913
rect 83455 53813 83466 53847
rect 83500 53813 83511 53847
rect 83455 53805 83511 53813
rect 83611 53943 83664 53955
rect 83611 53909 83622 53943
rect 83656 53909 83664 53943
rect 83611 53851 83664 53909
rect 83724 53942 83781 53984
rect 83724 53908 83736 53942
rect 83770 53908 83781 53942
rect 83724 53900 83781 53908
rect 83881 53976 83937 53984
rect 83881 53942 83892 53976
rect 83926 53942 83937 53976
rect 83881 53900 83937 53942
rect 84037 53942 84093 53984
rect 84037 53908 84048 53942
rect 84082 53908 84093 53942
rect 84037 53900 84093 53908
rect 84193 53950 84249 53984
rect 84193 53916 84204 53950
rect 84238 53916 84249 53950
rect 84193 53900 84249 53916
rect 84349 53900 84391 53984
rect 84491 53961 84563 53984
rect 84491 53927 84502 53961
rect 84536 53927 84563 53961
rect 84491 53900 84563 53927
rect 84663 53950 84720 53984
rect 84663 53916 84674 53950
rect 84708 53916 84720 53950
rect 84663 53900 84720 53916
rect 84834 53964 84846 53998
rect 84880 53964 84891 53998
rect 83611 53817 83622 53851
rect 83656 53817 83664 53851
rect 83611 53805 83664 53817
rect 84834 53811 84891 53964
rect 84991 53853 85047 54011
rect 84991 53819 85002 53853
rect 85036 53819 85047 53853
rect 84991 53811 85047 53819
rect 85147 54003 85204 54011
rect 85147 53969 85158 54003
rect 85192 53969 85204 54003
rect 85147 53928 85204 53969
rect 85147 53894 85158 53928
rect 85192 53895 85204 53928
rect 86108 53999 86161 54011
rect 86108 53965 86116 53999
rect 86150 53965 86161 53999
rect 86108 53919 86161 53965
rect 85192 53894 85226 53895
rect 85147 53853 85226 53894
rect 85147 53819 85158 53853
rect 85192 53819 85226 53853
rect 85147 53811 85226 53819
rect 85326 53811 85368 53895
rect 85468 53870 85545 53895
rect 85468 53836 85479 53870
rect 85513 53836 85545 53870
rect 85468 53811 85545 53836
rect 85645 53870 85701 53895
rect 85645 53836 85656 53870
rect 85690 53836 85701 53870
rect 85645 53811 85701 53836
rect 85801 53883 85858 53895
rect 85801 53849 85812 53883
rect 85846 53849 85858 53883
rect 86108 53885 86116 53919
rect 86150 53885 86161 53919
rect 86108 53861 86161 53885
rect 85801 53811 85858 53849
rect 85929 53853 85986 53861
rect 85929 53819 85941 53853
rect 85975 53819 85986 53853
rect 85929 53753 85986 53819
rect 85929 53719 85941 53753
rect 85975 53719 85986 53753
rect 85929 53711 85986 53719
rect 86086 53837 86161 53861
rect 86086 53803 86116 53837
rect 86150 53803 86161 53837
rect 86086 53757 86161 53803
rect 86086 53723 86116 53757
rect 86150 53723 86161 53757
rect 86086 53711 86161 53723
rect 86261 53999 86314 54011
rect 86261 53965 86272 53999
rect 86306 53965 86314 53999
rect 86261 53919 86314 53965
rect 86261 53885 86272 53919
rect 86306 53885 86314 53919
rect 86261 53837 86314 53885
rect 86261 53803 86272 53837
rect 86306 53803 86314 53837
rect 86261 53757 86314 53803
rect 86261 53723 86272 53757
rect 86306 53723 86314 53757
rect 86261 53711 86314 53723
rect 42112 50454 42712 50466
rect 42112 50420 42326 50454
rect 42498 50420 42712 50454
rect 42112 50408 42712 50420
rect 42806 50454 43406 50466
rect 42806 50420 43020 50454
rect 43192 50420 43406 50454
rect 42806 50408 43406 50420
rect 43500 50454 44100 50466
rect 43500 50420 43714 50454
rect 43886 50420 44100 50454
rect 43500 50408 44100 50420
rect 44194 50454 44794 50466
rect 44194 50420 44408 50454
rect 44580 50420 44794 50454
rect 44194 50408 44794 50420
rect 44888 50454 45488 50466
rect 44888 50420 45102 50454
rect 45274 50420 45488 50454
rect 44888 50408 45488 50420
rect 46106 50454 46706 50466
rect 46106 50420 46320 50454
rect 46492 50420 46706 50454
rect 46106 50408 46706 50420
rect 46800 50454 47400 50466
rect 46800 50420 47014 50454
rect 47186 50420 47400 50454
rect 46800 50408 47400 50420
rect 47494 50454 48094 50466
rect 47494 50420 47708 50454
rect 47880 50420 48094 50454
rect 47494 50408 48094 50420
rect 48188 50454 48788 50466
rect 48188 50420 48402 50454
rect 48574 50420 48788 50454
rect 48188 50408 48788 50420
rect 48882 50454 49482 50466
rect 48882 50420 49096 50454
rect 49268 50420 49482 50454
rect 48882 50408 49482 50420
rect 50128 50454 50728 50466
rect 50128 50420 50342 50454
rect 50514 50420 50728 50454
rect 50128 50408 50728 50420
rect 50822 50454 51422 50466
rect 50822 50420 51036 50454
rect 51208 50420 51422 50454
rect 50822 50408 51422 50420
rect 51516 50454 52116 50466
rect 51516 50420 51730 50454
rect 51902 50420 52116 50454
rect 51516 50408 52116 50420
rect 52210 50454 52810 50466
rect 52210 50420 52424 50454
rect 52596 50420 52810 50454
rect 52210 50408 52810 50420
rect 52904 50454 53504 50466
rect 52904 50420 53118 50454
rect 53290 50420 53504 50454
rect 52904 50408 53504 50420
rect 54150 50454 54750 50466
rect 54150 50420 54364 50454
rect 54536 50420 54750 50454
rect 54150 50408 54750 50420
rect 54844 50454 55444 50466
rect 54844 50420 55058 50454
rect 55230 50420 55444 50454
rect 54844 50408 55444 50420
rect 55538 50454 56138 50466
rect 55538 50420 55752 50454
rect 55924 50420 56138 50454
rect 55538 50408 56138 50420
rect 56232 50454 56832 50466
rect 56232 50420 56446 50454
rect 56618 50420 56832 50454
rect 56232 50408 56832 50420
rect 56926 50454 57526 50466
rect 56926 50420 57140 50454
rect 57312 50420 57526 50454
rect 56926 50408 57526 50420
rect 42112 49796 42712 49808
rect 42112 49762 42326 49796
rect 42498 49762 42712 49796
rect 42112 49750 42712 49762
rect 42806 49796 43406 49808
rect 42806 49762 43020 49796
rect 43192 49762 43406 49796
rect 42806 49750 43406 49762
rect 43500 49796 44100 49808
rect 43500 49762 43714 49796
rect 43886 49762 44100 49796
rect 43500 49750 44100 49762
rect 44194 49796 44794 49808
rect 44194 49762 44408 49796
rect 44580 49762 44794 49796
rect 44194 49750 44794 49762
rect 44888 49796 45488 49808
rect 44888 49762 45102 49796
rect 45274 49762 45488 49796
rect 44888 49750 45488 49762
rect 46106 49796 46706 49808
rect 46106 49762 46320 49796
rect 46492 49762 46706 49796
rect 46106 49750 46706 49762
rect 46800 49796 47400 49808
rect 46800 49762 47014 49796
rect 47186 49762 47400 49796
rect 46800 49750 47400 49762
rect 47494 49796 48094 49808
rect 47494 49762 47708 49796
rect 47880 49762 48094 49796
rect 47494 49750 48094 49762
rect 48188 49796 48788 49808
rect 48188 49762 48402 49796
rect 48574 49762 48788 49796
rect 48188 49750 48788 49762
rect 48882 49796 49482 49808
rect 48882 49762 49096 49796
rect 49268 49762 49482 49796
rect 48882 49750 49482 49762
rect 50128 49796 50728 49808
rect 50128 49762 50342 49796
rect 50514 49762 50728 49796
rect 50128 49750 50728 49762
rect 50822 49796 51422 49808
rect 50822 49762 51036 49796
rect 51208 49762 51422 49796
rect 50822 49750 51422 49762
rect 51516 49796 52116 49808
rect 51516 49762 51730 49796
rect 51902 49762 52116 49796
rect 51516 49750 52116 49762
rect 52210 49796 52810 49808
rect 52210 49762 52424 49796
rect 52596 49762 52810 49796
rect 52210 49750 52810 49762
rect 52904 49796 53504 49808
rect 52904 49762 53118 49796
rect 53290 49762 53504 49796
rect 52904 49750 53504 49762
rect 54150 49796 54750 49808
rect 54150 49762 54364 49796
rect 54536 49762 54750 49796
rect 54150 49750 54750 49762
rect 54844 49796 55444 49808
rect 54844 49762 55058 49796
rect 55230 49762 55444 49796
rect 54844 49750 55444 49762
rect 55538 49796 56138 49808
rect 55538 49762 55752 49796
rect 55924 49762 56138 49796
rect 55538 49750 56138 49762
rect 56232 49796 56832 49808
rect 56232 49762 56446 49796
rect 56618 49762 56832 49796
rect 56232 49750 56832 49762
rect 56926 49796 57526 49808
rect 56926 49762 57140 49796
rect 57312 49762 57526 49796
rect 56926 49750 57526 49762
rect 42112 49138 42712 49150
rect 42112 49104 42326 49138
rect 42498 49104 42712 49138
rect 42112 49092 42712 49104
rect 42806 49138 43406 49150
rect 42806 49104 43020 49138
rect 43192 49104 43406 49138
rect 42806 49092 43406 49104
rect 43500 49138 44100 49150
rect 43500 49104 43714 49138
rect 43886 49104 44100 49138
rect 43500 49092 44100 49104
rect 44194 49138 44794 49150
rect 44194 49104 44408 49138
rect 44580 49104 44794 49138
rect 44194 49092 44794 49104
rect 44888 49138 45488 49150
rect 44888 49104 45102 49138
rect 45274 49104 45488 49138
rect 44888 49092 45488 49104
rect 46106 49138 46706 49150
rect 46106 49104 46320 49138
rect 46492 49104 46706 49138
rect 46106 49092 46706 49104
rect 46800 49138 47400 49150
rect 46800 49104 47014 49138
rect 47186 49104 47400 49138
rect 46800 49092 47400 49104
rect 47494 49138 48094 49150
rect 47494 49104 47708 49138
rect 47880 49104 48094 49138
rect 47494 49092 48094 49104
rect 48188 49138 48788 49150
rect 48188 49104 48402 49138
rect 48574 49104 48788 49138
rect 48188 49092 48788 49104
rect 48882 49138 49482 49150
rect 48882 49104 49096 49138
rect 49268 49104 49482 49138
rect 48882 49092 49482 49104
rect 50128 49138 50728 49150
rect 50128 49104 50342 49138
rect 50514 49104 50728 49138
rect 50128 49092 50728 49104
rect 50822 49138 51422 49150
rect 50822 49104 51036 49138
rect 51208 49104 51422 49138
rect 50822 49092 51422 49104
rect 51516 49138 52116 49150
rect 51516 49104 51730 49138
rect 51902 49104 52116 49138
rect 51516 49092 52116 49104
rect 52210 49138 52810 49150
rect 52210 49104 52424 49138
rect 52596 49104 52810 49138
rect 52210 49092 52810 49104
rect 52904 49138 53504 49150
rect 52904 49104 53118 49138
rect 53290 49104 53504 49138
rect 52904 49092 53504 49104
rect 54150 49138 54750 49150
rect 54150 49104 54364 49138
rect 54536 49104 54750 49138
rect 54150 49092 54750 49104
rect 54844 49138 55444 49150
rect 54844 49104 55058 49138
rect 55230 49104 55444 49138
rect 54844 49092 55444 49104
rect 55538 49138 56138 49150
rect 55538 49104 55752 49138
rect 55924 49104 56138 49138
rect 55538 49092 56138 49104
rect 56232 49138 56832 49150
rect 56232 49104 56446 49138
rect 56618 49104 56832 49138
rect 56232 49092 56832 49104
rect 56926 49138 57526 49150
rect 56926 49104 57140 49138
rect 57312 49104 57526 49138
rect 56926 49092 57526 49104
rect 42112 48480 42712 48492
rect 42112 48446 42326 48480
rect 42498 48446 42712 48480
rect 42112 48434 42712 48446
rect 42806 48480 43406 48492
rect 42806 48446 43020 48480
rect 43192 48446 43406 48480
rect 42806 48434 43406 48446
rect 43500 48480 44100 48492
rect 43500 48446 43714 48480
rect 43886 48446 44100 48480
rect 43500 48434 44100 48446
rect 44194 48480 44794 48492
rect 44194 48446 44408 48480
rect 44580 48446 44794 48480
rect 44194 48434 44794 48446
rect 44888 48480 45488 48492
rect 44888 48446 45102 48480
rect 45274 48446 45488 48480
rect 44888 48434 45488 48446
rect 46106 48480 46706 48492
rect 46106 48446 46320 48480
rect 46492 48446 46706 48480
rect 46106 48434 46706 48446
rect 46800 48480 47400 48492
rect 46800 48446 47014 48480
rect 47186 48446 47400 48480
rect 46800 48434 47400 48446
rect 47494 48480 48094 48492
rect 47494 48446 47708 48480
rect 47880 48446 48094 48480
rect 47494 48434 48094 48446
rect 48188 48480 48788 48492
rect 48188 48446 48402 48480
rect 48574 48446 48788 48480
rect 48188 48434 48788 48446
rect 48882 48480 49482 48492
rect 48882 48446 49096 48480
rect 49268 48446 49482 48480
rect 48882 48434 49482 48446
rect 50128 48480 50728 48492
rect 50128 48446 50342 48480
rect 50514 48446 50728 48480
rect 50128 48434 50728 48446
rect 50822 48480 51422 48492
rect 50822 48446 51036 48480
rect 51208 48446 51422 48480
rect 50822 48434 51422 48446
rect 51516 48480 52116 48492
rect 51516 48446 51730 48480
rect 51902 48446 52116 48480
rect 51516 48434 52116 48446
rect 52210 48480 52810 48492
rect 52210 48446 52424 48480
rect 52596 48446 52810 48480
rect 52210 48434 52810 48446
rect 52904 48480 53504 48492
rect 52904 48446 53118 48480
rect 53290 48446 53504 48480
rect 52904 48434 53504 48446
rect 54150 48480 54750 48492
rect 54150 48446 54364 48480
rect 54536 48446 54750 48480
rect 54150 48434 54750 48446
rect 54844 48480 55444 48492
rect 54844 48446 55058 48480
rect 55230 48446 55444 48480
rect 54844 48434 55444 48446
rect 55538 48480 56138 48492
rect 55538 48446 55752 48480
rect 55924 48446 56138 48480
rect 55538 48434 56138 48446
rect 56232 48480 56832 48492
rect 56232 48446 56446 48480
rect 56618 48446 56832 48480
rect 56232 48434 56832 48446
rect 56926 48480 57526 48492
rect 56926 48446 57140 48480
rect 57312 48446 57526 48480
rect 56926 48434 57526 48446
<< mvndiffc >>
rect 23634 57446 23806 57480
rect 24328 57446 24500 57480
rect 25022 57446 25194 57480
rect 25716 57446 25888 57480
rect 26410 57446 26582 57480
rect 27104 57446 27276 57480
rect 27798 57446 27970 57480
rect 28492 57446 28664 57480
rect 29186 57446 29358 57480
rect 29880 57446 30052 57480
rect 23634 56788 23806 56822
rect 24328 56788 24500 56822
rect 25022 56788 25194 56822
rect 25716 56788 25888 56822
rect 26410 56788 26582 56822
rect 27104 56788 27276 56822
rect 27798 56788 27970 56822
rect 28492 56788 28664 56822
rect 29186 56788 29358 56822
rect 29880 56788 30052 56822
rect 23634 56130 23806 56164
rect 24328 56130 24500 56164
rect 25022 56130 25194 56164
rect 25716 56130 25888 56164
rect 26410 56130 26582 56164
rect 27104 56130 27276 56164
rect 27798 56130 27970 56164
rect 28492 56130 28664 56164
rect 29186 56130 29358 56164
rect 29880 56130 30052 56164
rect 23640 55556 23812 55590
rect 24334 55556 24506 55590
rect 25028 55556 25200 55590
rect 25722 55556 25894 55590
rect 26416 55556 26588 55590
rect 27110 55556 27282 55590
rect 27804 55556 27976 55590
rect 28498 55556 28670 55590
rect 29192 55556 29364 55590
rect 29886 55556 30058 55590
rect 23640 54898 23812 54932
rect 24334 54898 24506 54932
rect 25028 54898 25200 54932
rect 25722 54898 25894 54932
rect 26416 54898 26588 54932
rect 27110 54898 27282 54932
rect 27804 54898 27976 54932
rect 28498 54898 28670 54932
rect 29192 54898 29364 54932
rect 29886 54898 30058 54932
rect 23640 54240 23812 54274
rect 24334 54240 24506 54274
rect 25028 54240 25200 54274
rect 25722 54240 25894 54274
rect 26416 54240 26588 54274
rect 27110 54240 27282 54274
rect 27804 54240 27976 54274
rect 28498 54240 28670 54274
rect 29192 54240 29364 54274
rect 29886 54240 30058 54274
rect 23656 53614 23828 53648
rect 24350 53614 24522 53648
rect 25044 53614 25216 53648
rect 25738 53614 25910 53648
rect 26432 53614 26604 53648
rect 27126 53614 27298 53648
rect 27820 53614 27992 53648
rect 28514 53614 28686 53648
rect 29208 53614 29380 53648
rect 29902 53614 30074 53648
rect 23656 52956 23828 52990
rect 24350 52956 24522 52990
rect 25044 52956 25216 52990
rect 25738 52956 25910 52990
rect 26432 52956 26604 52990
rect 27126 52956 27298 52990
rect 27820 52956 27992 52990
rect 28514 52956 28686 52990
rect 29208 52956 29380 52990
rect 29902 52956 30074 52990
rect 23656 52298 23828 52332
rect 24350 52298 24522 52332
rect 25044 52298 25216 52332
rect 25738 52298 25910 52332
rect 26432 52298 26604 52332
rect 27126 52298 27298 52332
rect 27820 52298 27992 52332
rect 28514 52298 28686 52332
rect 29208 52298 29380 52332
rect 29902 52298 30074 52332
rect 83764 53466 83798 53500
rect 83314 53400 83348 53434
rect 83470 53400 83504 53434
rect 84062 53466 84096 53500
rect 84218 53466 84252 53500
rect 83626 53400 83660 53434
rect 84844 53403 84878 53437
rect 85016 53483 85050 53517
rect 85016 53391 85050 53425
rect 85174 53483 85208 53517
rect 85933 53500 85967 53534
rect 86112 53517 86146 53551
rect 85174 53391 85208 53425
rect 85514 53400 85548 53434
rect 85812 53400 85846 53434
rect 86112 53417 86146 53451
rect 86268 53517 86302 53551
rect 86268 53417 86302 53451
rect 1958 42760 1992 43052
rect 3016 42760 3050 43052
rect 4074 42760 4108 43052
rect 5132 42760 5166 43052
rect 6190 42760 6224 43052
rect 7248 42760 7282 43052
rect 8472 42768 8506 43060
rect 9530 42768 9564 43060
rect 10588 42768 10622 43060
rect 11646 42768 11680 43060
rect 12704 42768 12738 43060
rect 13762 42768 13796 43060
rect 14978 42776 15012 43068
rect 16036 42776 16070 43068
rect 17094 42776 17128 43068
rect 18152 42776 18186 43068
rect 19210 42776 19244 43068
rect 20268 42776 20302 43068
rect 21468 42760 21502 43052
rect 22526 42760 22560 43052
rect 23584 42760 23618 43052
rect 24642 42760 24676 43052
rect 25700 42760 25734 43052
rect 26758 42760 26792 43052
rect 27990 42776 28024 43068
rect 29048 42776 29082 43068
rect 30106 42776 30140 43068
rect 31164 42776 31198 43068
rect 32222 42776 32256 43068
rect 33280 42776 33314 43068
rect 34500 42782 34534 43074
rect 35558 42782 35592 43074
rect 36616 42782 36650 43074
rect 37674 42782 37708 43074
rect 38732 42782 38766 43074
rect 39790 42782 39824 43074
rect 40990 42782 41024 43074
rect 42048 42782 42082 43074
rect 43106 42782 43140 43074
rect 44164 42782 44198 43074
rect 45222 42782 45256 43074
rect 46280 42782 46314 43074
rect 47578 42804 47612 43096
rect 48636 42804 48670 43096
rect 49694 42804 49728 43096
rect 50752 42804 50786 43096
rect 51810 42804 51844 43096
rect 52868 42804 52902 43096
rect 54092 42818 54126 43110
rect 55150 42818 55184 43110
rect 56208 42818 56242 43110
rect 57266 42818 57300 43110
rect 58324 42818 58358 43110
rect 59382 42818 59416 43110
rect 1958 41666 1992 41958
rect 3016 41666 3050 41958
rect 4074 41666 4108 41958
rect 5132 41666 5166 41958
rect 6190 41666 6224 41958
rect 7248 41666 7282 41958
rect 1958 40572 1992 40864
rect 3016 40572 3050 40864
rect 4074 40572 4108 40864
rect 5132 40572 5166 40864
rect 6190 40572 6224 40864
rect 7248 40572 7282 40864
rect 8472 41674 8506 41966
rect 9530 41674 9564 41966
rect 10588 41674 10622 41966
rect 11646 41674 11680 41966
rect 12704 41674 12738 41966
rect 13762 41674 13796 41966
rect 1958 39478 1992 39770
rect 3016 39478 3050 39770
rect 4074 39478 4108 39770
rect 5132 39478 5166 39770
rect 6190 39478 6224 39770
rect 8472 40580 8506 40872
rect 9530 40580 9564 40872
rect 10588 40580 10622 40872
rect 11646 40580 11680 40872
rect 12704 40580 12738 40872
rect 13762 40580 13796 40872
rect 14978 41682 15012 41974
rect 16036 41682 16070 41974
rect 17094 41682 17128 41974
rect 18152 41682 18186 41974
rect 19210 41682 19244 41974
rect 20268 41682 20302 41974
rect 7248 39478 7282 39770
rect 8472 39486 8506 39778
rect 9530 39486 9564 39778
rect 10588 39486 10622 39778
rect 11646 39486 11680 39778
rect 12704 39486 12738 39778
rect 14978 40588 15012 40880
rect 16036 40588 16070 40880
rect 17094 40588 17128 40880
rect 18152 40588 18186 40880
rect 19210 40588 19244 40880
rect 20268 40588 20302 40880
rect 21468 41666 21502 41958
rect 22526 41666 22560 41958
rect 23584 41666 23618 41958
rect 24642 41666 24676 41958
rect 25700 41666 25734 41958
rect 26758 41666 26792 41958
rect 13762 39486 13796 39778
rect 14978 39494 15012 39786
rect 16036 39494 16070 39786
rect 17094 39494 17128 39786
rect 18152 39494 18186 39786
rect 19210 39494 19244 39786
rect 21468 40572 21502 40864
rect 22526 40572 22560 40864
rect 23584 40572 23618 40864
rect 24642 40572 24676 40864
rect 25700 40572 25734 40864
rect 26758 40572 26792 40864
rect 27990 41682 28024 41974
rect 29048 41682 29082 41974
rect 30106 41682 30140 41974
rect 31164 41682 31198 41974
rect 32222 41682 32256 41974
rect 33280 41682 33314 41974
rect 20268 39494 20302 39786
rect 21468 39478 21502 39770
rect 22526 39478 22560 39770
rect 23584 39478 23618 39770
rect 24642 39478 24676 39770
rect 25700 39478 25734 39770
rect 27990 40588 28024 40880
rect 29048 40588 29082 40880
rect 30106 40588 30140 40880
rect 31164 40588 31198 40880
rect 32222 40588 32256 40880
rect 33280 40588 33314 40880
rect 34500 41688 34534 41980
rect 35558 41688 35592 41980
rect 36616 41688 36650 41980
rect 37674 41688 37708 41980
rect 38732 41688 38766 41980
rect 39790 41688 39824 41980
rect 26758 39478 26792 39770
rect 27990 39494 28024 39786
rect 29048 39494 29082 39786
rect 30106 39494 30140 39786
rect 31164 39494 31198 39786
rect 32222 39494 32256 39786
rect 34500 40594 34534 40886
rect 35558 40594 35592 40886
rect 36616 40594 36650 40886
rect 37674 40594 37708 40886
rect 38732 40594 38766 40886
rect 39790 40594 39824 40886
rect 40990 41688 41024 41980
rect 42048 41688 42082 41980
rect 43106 41688 43140 41980
rect 44164 41688 44198 41980
rect 45222 41688 45256 41980
rect 46280 41688 46314 41980
rect 33280 39494 33314 39786
rect 34500 39500 34534 39792
rect 35558 39500 35592 39792
rect 36616 39500 36650 39792
rect 37674 39500 37708 39792
rect 38732 39500 38766 39792
rect 40990 40594 41024 40886
rect 42048 40594 42082 40886
rect 43106 40594 43140 40886
rect 44164 40594 44198 40886
rect 45222 40594 45256 40886
rect 46280 40594 46314 40886
rect 47578 41710 47612 42002
rect 48636 41710 48670 42002
rect 49694 41710 49728 42002
rect 50752 41710 50786 42002
rect 51810 41710 51844 42002
rect 52868 41710 52902 42002
rect 39790 39500 39824 39792
rect 40990 39500 41024 39792
rect 42048 39500 42082 39792
rect 43106 39500 43140 39792
rect 44164 39500 44198 39792
rect 45222 39500 45256 39792
rect 47578 40616 47612 40908
rect 48636 40616 48670 40908
rect 49694 40616 49728 40908
rect 50752 40616 50786 40908
rect 51810 40616 51844 40908
rect 52868 40616 52902 40908
rect 54092 41724 54126 42016
rect 55150 41724 55184 42016
rect 56208 41724 56242 42016
rect 57266 41724 57300 42016
rect 58324 41724 58358 42016
rect 59382 41724 59416 42016
rect 46280 39500 46314 39792
rect 47578 39522 47612 39814
rect 48636 39522 48670 39814
rect 49694 39522 49728 39814
rect 50752 39522 50786 39814
rect 51810 39522 51844 39814
rect 54092 40630 54126 40922
rect 55150 40630 55184 40922
rect 56208 40630 56242 40922
rect 57266 40630 57300 40922
rect 58324 40630 58358 40922
rect 59382 40630 59416 40922
rect 52868 39522 52902 39814
rect 54092 39536 54126 39828
rect 55150 39536 55184 39828
rect 56208 39536 56242 39828
rect 57266 39536 57300 39828
rect 58324 39536 58358 39828
rect 59382 39536 59416 39828
rect 1958 38384 1992 38676
rect 3016 38384 3050 38676
rect 4074 38384 4108 38676
rect 5132 38384 5166 38676
rect 6190 38384 6224 38676
rect 7248 38384 7282 38676
rect 8472 38392 8506 38684
rect 9530 38392 9564 38684
rect 10588 38392 10622 38684
rect 11646 38392 11680 38684
rect 12704 38392 12738 38684
rect 13762 38392 13796 38684
rect 14978 38400 15012 38692
rect 16036 38400 16070 38692
rect 17094 38400 17128 38692
rect 18152 38400 18186 38692
rect 19210 38400 19244 38692
rect 20268 38400 20302 38692
rect 21468 38384 21502 38676
rect 22526 38384 22560 38676
rect 23584 38384 23618 38676
rect 24642 38384 24676 38676
rect 25700 38384 25734 38676
rect 26758 38384 26792 38676
rect 27990 38400 28024 38692
rect 29048 38400 29082 38692
rect 30106 38400 30140 38692
rect 31164 38400 31198 38692
rect 32222 38400 32256 38692
rect 33280 38400 33314 38692
rect 34500 38406 34534 38698
rect 35558 38406 35592 38698
rect 36616 38406 36650 38698
rect 37674 38406 37708 38698
rect 38732 38406 38766 38698
rect 39790 38406 39824 38698
rect 40990 38406 41024 38698
rect 42048 38406 42082 38698
rect 43106 38406 43140 38698
rect 44164 38406 44198 38698
rect 45222 38406 45256 38698
rect 46280 38406 46314 38698
rect 47578 38428 47612 38720
rect 48636 38428 48670 38720
rect 49694 38428 49728 38720
rect 50752 38428 50786 38720
rect 51810 38428 51844 38720
rect 52868 38428 52902 38720
rect 54092 38442 54126 38734
rect 55150 38442 55184 38734
rect 56208 38442 56242 38734
rect 57266 38442 57300 38734
rect 58324 38442 58358 38734
rect 59382 38442 59416 38734
rect 1958 36944 1992 37236
rect 3016 36944 3050 37236
rect 4074 36944 4108 37236
rect 5132 36944 5166 37236
rect 6190 36944 6224 37236
rect 7248 36944 7282 37236
rect 8472 36952 8506 37244
rect 9530 36952 9564 37244
rect 10588 36952 10622 37244
rect 11646 36952 11680 37244
rect 12704 36952 12738 37244
rect 13762 36952 13796 37244
rect 14978 36960 15012 37252
rect 16036 36960 16070 37252
rect 17094 36960 17128 37252
rect 18152 36960 18186 37252
rect 19210 36960 19244 37252
rect 20268 36960 20302 37252
rect 21468 36944 21502 37236
rect 22526 36944 22560 37236
rect 23584 36944 23618 37236
rect 24642 36944 24676 37236
rect 25700 36944 25734 37236
rect 26758 36944 26792 37236
rect 27990 36960 28024 37252
rect 29048 36960 29082 37252
rect 30106 36960 30140 37252
rect 31164 36960 31198 37252
rect 32222 36960 32256 37252
rect 33280 36960 33314 37252
rect 34500 36966 34534 37258
rect 35558 36966 35592 37258
rect 36616 36966 36650 37258
rect 37674 36966 37708 37258
rect 38732 36966 38766 37258
rect 39790 36966 39824 37258
rect 40990 36966 41024 37258
rect 42048 36966 42082 37258
rect 43106 36966 43140 37258
rect 44164 36966 44198 37258
rect 45222 36966 45256 37258
rect 46280 36966 46314 37258
rect 47578 36988 47612 37280
rect 48636 36988 48670 37280
rect 49694 36988 49728 37280
rect 50752 36988 50786 37280
rect 51810 36988 51844 37280
rect 52868 36988 52902 37280
rect 54092 37002 54126 37294
rect 55150 37002 55184 37294
rect 56208 37002 56242 37294
rect 57266 37002 57300 37294
rect 58324 37002 58358 37294
rect 59382 37002 59416 37294
rect 1958 35850 1992 36142
rect 3016 35850 3050 36142
rect 4074 35850 4108 36142
rect 5132 35850 5166 36142
rect 6190 35850 6224 36142
rect 7248 35850 7282 36142
rect 1958 34756 1992 35048
rect 3016 34756 3050 35048
rect 4074 34756 4108 35048
rect 5132 34756 5166 35048
rect 6190 34756 6224 35048
rect 7248 34756 7282 35048
rect 8472 35858 8506 36150
rect 9530 35858 9564 36150
rect 10588 35858 10622 36150
rect 11646 35858 11680 36150
rect 12704 35858 12738 36150
rect 13762 35858 13796 36150
rect 1958 33662 1992 33954
rect 3016 33662 3050 33954
rect 4074 33662 4108 33954
rect 5132 33662 5166 33954
rect 6190 33662 6224 33954
rect 8472 34764 8506 35056
rect 9530 34764 9564 35056
rect 10588 34764 10622 35056
rect 11646 34764 11680 35056
rect 12704 34764 12738 35056
rect 13762 34764 13796 35056
rect 14978 35866 15012 36158
rect 16036 35866 16070 36158
rect 17094 35866 17128 36158
rect 18152 35866 18186 36158
rect 19210 35866 19244 36158
rect 20268 35866 20302 36158
rect 7248 33662 7282 33954
rect 8472 33670 8506 33962
rect 9530 33670 9564 33962
rect 10588 33670 10622 33962
rect 11646 33670 11680 33962
rect 12704 33670 12738 33962
rect 14978 34772 15012 35064
rect 16036 34772 16070 35064
rect 17094 34772 17128 35064
rect 18152 34772 18186 35064
rect 19210 34772 19244 35064
rect 20268 34772 20302 35064
rect 21468 35850 21502 36142
rect 22526 35850 22560 36142
rect 23584 35850 23618 36142
rect 24642 35850 24676 36142
rect 25700 35850 25734 36142
rect 26758 35850 26792 36142
rect 13762 33670 13796 33962
rect 14978 33678 15012 33970
rect 16036 33678 16070 33970
rect 17094 33678 17128 33970
rect 18152 33678 18186 33970
rect 19210 33678 19244 33970
rect 21468 34756 21502 35048
rect 22526 34756 22560 35048
rect 23584 34756 23618 35048
rect 24642 34756 24676 35048
rect 25700 34756 25734 35048
rect 26758 34756 26792 35048
rect 27990 35866 28024 36158
rect 29048 35866 29082 36158
rect 30106 35866 30140 36158
rect 31164 35866 31198 36158
rect 32222 35866 32256 36158
rect 33280 35866 33314 36158
rect 20268 33678 20302 33970
rect 21468 33662 21502 33954
rect 22526 33662 22560 33954
rect 23584 33662 23618 33954
rect 24642 33662 24676 33954
rect 25700 33662 25734 33954
rect 27990 34772 28024 35064
rect 29048 34772 29082 35064
rect 30106 34772 30140 35064
rect 31164 34772 31198 35064
rect 32222 34772 32256 35064
rect 33280 34772 33314 35064
rect 34500 35872 34534 36164
rect 35558 35872 35592 36164
rect 36616 35872 36650 36164
rect 37674 35872 37708 36164
rect 38732 35872 38766 36164
rect 39790 35872 39824 36164
rect 26758 33662 26792 33954
rect 27990 33678 28024 33970
rect 29048 33678 29082 33970
rect 30106 33678 30140 33970
rect 31164 33678 31198 33970
rect 32222 33678 32256 33970
rect 34500 34778 34534 35070
rect 35558 34778 35592 35070
rect 36616 34778 36650 35070
rect 37674 34778 37708 35070
rect 38732 34778 38766 35070
rect 39790 34778 39824 35070
rect 40990 35872 41024 36164
rect 42048 35872 42082 36164
rect 43106 35872 43140 36164
rect 44164 35872 44198 36164
rect 45222 35872 45256 36164
rect 46280 35872 46314 36164
rect 33280 33678 33314 33970
rect 34500 33684 34534 33976
rect 35558 33684 35592 33976
rect 36616 33684 36650 33976
rect 37674 33684 37708 33976
rect 38732 33684 38766 33976
rect 40990 34778 41024 35070
rect 42048 34778 42082 35070
rect 43106 34778 43140 35070
rect 44164 34778 44198 35070
rect 45222 34778 45256 35070
rect 46280 34778 46314 35070
rect 47578 35894 47612 36186
rect 48636 35894 48670 36186
rect 49694 35894 49728 36186
rect 50752 35894 50786 36186
rect 51810 35894 51844 36186
rect 52868 35894 52902 36186
rect 39790 33684 39824 33976
rect 40990 33684 41024 33976
rect 42048 33684 42082 33976
rect 43106 33684 43140 33976
rect 44164 33684 44198 33976
rect 45222 33684 45256 33976
rect 47578 34800 47612 35092
rect 48636 34800 48670 35092
rect 49694 34800 49728 35092
rect 50752 34800 50786 35092
rect 51810 34800 51844 35092
rect 52868 34800 52902 35092
rect 54092 35908 54126 36200
rect 55150 35908 55184 36200
rect 56208 35908 56242 36200
rect 57266 35908 57300 36200
rect 58324 35908 58358 36200
rect 59382 35908 59416 36200
rect 62508 42936 62542 43108
rect 63166 42936 63200 43108
rect 63824 42936 63858 43108
rect 64482 42936 64516 43108
rect 65140 42936 65174 43108
rect 65798 42936 65832 43108
rect 66302 42938 66336 43110
rect 66960 42938 66994 43110
rect 67618 42938 67652 43110
rect 68276 42938 68310 43110
rect 68934 42938 68968 43110
rect 69592 42938 69626 43110
rect 70110 42952 70144 43124
rect 70768 42952 70802 43124
rect 71426 42952 71460 43124
rect 72084 42952 72118 43124
rect 72742 42952 72776 43124
rect 73400 42952 73434 43124
rect 62508 42242 62542 42414
rect 63166 42242 63200 42414
rect 63824 42242 63858 42414
rect 64482 42242 64516 42414
rect 65140 42242 65174 42414
rect 65798 42242 65832 42414
rect 62508 41548 62542 41720
rect 63166 41548 63200 41720
rect 63824 41548 63858 41720
rect 64482 41548 64516 41720
rect 65140 41548 65174 41720
rect 65798 41548 65832 41720
rect 62508 40854 62542 41026
rect 63166 40854 63200 41026
rect 63824 40854 63858 41026
rect 64482 40854 64516 41026
rect 65140 40854 65174 41026
rect 65798 40854 65832 41026
rect 66302 42244 66336 42416
rect 66960 42244 66994 42416
rect 67618 42244 67652 42416
rect 68276 42244 68310 42416
rect 68934 42244 68968 42416
rect 69592 42244 69626 42416
rect 66302 41550 66336 41722
rect 66960 41550 66994 41722
rect 67618 41550 67652 41722
rect 68276 41550 68310 41722
rect 68934 41550 68968 41722
rect 69592 41550 69626 41722
rect 66302 40856 66336 41028
rect 66960 40856 66994 41028
rect 67618 40856 67652 41028
rect 68276 40856 68310 41028
rect 68934 40856 68968 41028
rect 69592 40856 69626 41028
rect 70110 42258 70144 42430
rect 70768 42258 70802 42430
rect 71426 42258 71460 42430
rect 72084 42258 72118 42430
rect 72742 42258 72776 42430
rect 73400 42258 73434 42430
rect 70110 41564 70144 41736
rect 70768 41564 70802 41736
rect 71426 41564 71460 41736
rect 72084 41564 72118 41736
rect 72742 41564 72776 41736
rect 73400 41564 73434 41736
rect 70110 40870 70144 41042
rect 70768 40870 70802 41042
rect 71426 40870 71460 41042
rect 72084 40870 72118 41042
rect 72742 40870 72776 41042
rect 73400 40870 73434 41042
rect 62508 40160 62542 40332
rect 63166 40160 63200 40332
rect 63824 40160 63858 40332
rect 64482 40160 64516 40332
rect 65140 40160 65174 40332
rect 65798 40160 65832 40332
rect 66302 40162 66336 40334
rect 66960 40162 66994 40334
rect 67618 40162 67652 40334
rect 68276 40162 68310 40334
rect 68934 40162 68968 40334
rect 69592 40162 69626 40334
rect 70110 40176 70144 40348
rect 70768 40176 70802 40348
rect 71426 40176 71460 40348
rect 72084 40176 72118 40348
rect 72742 40176 72776 40348
rect 73400 40176 73434 40348
rect 46280 33684 46314 33976
rect 47578 33706 47612 33998
rect 48636 33706 48670 33998
rect 49694 33706 49728 33998
rect 50752 33706 50786 33998
rect 51810 33706 51844 33998
rect 54092 34814 54126 35106
rect 55150 34814 55184 35106
rect 56208 34814 56242 35106
rect 57266 34814 57300 35106
rect 58324 34814 58358 35106
rect 59382 34814 59416 35106
rect 77170 38922 77204 39094
rect 77828 38922 77862 39094
rect 78486 38922 78520 39094
rect 79144 38922 79178 39094
rect 79802 38922 79836 39094
rect 77170 38228 77204 38400
rect 77828 38228 77862 38400
rect 78486 38228 78520 38400
rect 79144 38228 79178 38400
rect 79802 38228 79836 38400
rect 77170 37534 77204 37706
rect 77828 37534 77862 37706
rect 78486 37534 78520 37706
rect 79144 37534 79178 37706
rect 79802 37534 79836 37706
rect 77170 36840 77204 37012
rect 77828 36840 77862 37012
rect 78486 36840 78520 37012
rect 79144 36840 79178 37012
rect 79802 36840 79836 37012
rect 77170 36146 77204 36318
rect 77828 36146 77862 36318
rect 78486 36146 78520 36318
rect 79144 36146 79178 36318
rect 79802 36146 79836 36318
rect 77170 35452 77204 35624
rect 77828 35452 77862 35624
rect 78486 35452 78520 35624
rect 79144 35452 79178 35624
rect 79802 35452 79836 35624
rect 80496 38916 80530 39088
rect 81154 38916 81188 39088
rect 81812 38916 81846 39088
rect 82470 38916 82504 39088
rect 83128 38916 83162 39088
rect 80496 38222 80530 38394
rect 81154 38222 81188 38394
rect 81812 38222 81846 38394
rect 82470 38222 82504 38394
rect 83128 38222 83162 38394
rect 80496 37528 80530 37700
rect 81154 37528 81188 37700
rect 81812 37528 81846 37700
rect 82470 37528 82504 37700
rect 83128 37528 83162 37700
rect 80496 36834 80530 37006
rect 81154 36834 81188 37006
rect 81812 36834 81846 37006
rect 82470 36834 82504 37006
rect 83128 36834 83162 37006
rect 80496 36140 80530 36312
rect 81154 36140 81188 36312
rect 81812 36140 81846 36312
rect 82470 36140 82504 36312
rect 83128 36140 83162 36312
rect 80496 35446 80530 35618
rect 81154 35446 81188 35618
rect 81812 35446 81846 35618
rect 82470 35446 82504 35618
rect 83128 35446 83162 35618
rect 83806 38916 83840 39088
rect 84464 38916 84498 39088
rect 85122 38916 85156 39088
rect 85780 38916 85814 39088
rect 86438 38916 86472 39088
rect 83806 38222 83840 38394
rect 84464 38222 84498 38394
rect 85122 38222 85156 38394
rect 85780 38222 85814 38394
rect 86438 38222 86472 38394
rect 83806 37528 83840 37700
rect 84464 37528 84498 37700
rect 85122 37528 85156 37700
rect 85780 37528 85814 37700
rect 86438 37528 86472 37700
rect 83806 36834 83840 37006
rect 84464 36834 84498 37006
rect 85122 36834 85156 37006
rect 85780 36834 85814 37006
rect 86438 36834 86472 37006
rect 83806 36140 83840 36312
rect 84464 36140 84498 36312
rect 85122 36140 85156 36312
rect 85780 36140 85814 36312
rect 86438 36140 86472 36312
rect 83806 35446 83840 35618
rect 84464 35446 84498 35618
rect 85122 35446 85156 35618
rect 85780 35446 85814 35618
rect 86438 35446 86472 35618
rect 52868 33706 52902 33998
rect 54092 33720 54126 34012
rect 55150 33720 55184 34012
rect 56208 33720 56242 34012
rect 57266 33720 57300 34012
rect 58324 33720 58358 34012
rect 59382 33720 59416 34012
rect 1958 32568 1992 32860
rect 3016 32568 3050 32860
rect 4074 32568 4108 32860
rect 5132 32568 5166 32860
rect 6190 32568 6224 32860
rect 7248 32568 7282 32860
rect 8472 32576 8506 32868
rect 9530 32576 9564 32868
rect 10588 32576 10622 32868
rect 11646 32576 11680 32868
rect 12704 32576 12738 32868
rect 13762 32576 13796 32868
rect 14978 32584 15012 32876
rect 16036 32584 16070 32876
rect 17094 32584 17128 32876
rect 18152 32584 18186 32876
rect 19210 32584 19244 32876
rect 20268 32584 20302 32876
rect 21468 32568 21502 32860
rect 22526 32568 22560 32860
rect 23584 32568 23618 32860
rect 24642 32568 24676 32860
rect 25700 32568 25734 32860
rect 26758 32568 26792 32860
rect 27990 32584 28024 32876
rect 29048 32584 29082 32876
rect 30106 32584 30140 32876
rect 31164 32584 31198 32876
rect 32222 32584 32256 32876
rect 33280 32584 33314 32876
rect 34500 32590 34534 32882
rect 35558 32590 35592 32882
rect 36616 32590 36650 32882
rect 37674 32590 37708 32882
rect 38732 32590 38766 32882
rect 39790 32590 39824 32882
rect 40990 32590 41024 32882
rect 42048 32590 42082 32882
rect 43106 32590 43140 32882
rect 44164 32590 44198 32882
rect 45222 32590 45256 32882
rect 46280 32590 46314 32882
rect 47578 32612 47612 32904
rect 48636 32612 48670 32904
rect 49694 32612 49728 32904
rect 50752 32612 50786 32904
rect 51810 32612 51844 32904
rect 52868 32612 52902 32904
rect 54092 32626 54126 32918
rect 55150 32626 55184 32918
rect 56208 32626 56242 32918
rect 57266 32626 57300 32918
rect 58324 32626 58358 32918
rect 59382 32626 59416 32918
rect 1958 31110 1992 31402
rect 3016 31110 3050 31402
rect 4074 31110 4108 31402
rect 5132 31110 5166 31402
rect 6190 31110 6224 31402
rect 7248 31110 7282 31402
rect 8472 31118 8506 31410
rect 9530 31118 9564 31410
rect 10588 31118 10622 31410
rect 11646 31118 11680 31410
rect 12704 31118 12738 31410
rect 13762 31118 13796 31410
rect 14978 31126 15012 31418
rect 16036 31126 16070 31418
rect 17094 31126 17128 31418
rect 18152 31126 18186 31418
rect 19210 31126 19244 31418
rect 20268 31126 20302 31418
rect 21468 31110 21502 31402
rect 22526 31110 22560 31402
rect 23584 31110 23618 31402
rect 24642 31110 24676 31402
rect 25700 31110 25734 31402
rect 26758 31110 26792 31402
rect 27990 31126 28024 31418
rect 29048 31126 29082 31418
rect 30106 31126 30140 31418
rect 31164 31126 31198 31418
rect 32222 31126 32256 31418
rect 33280 31126 33314 31418
rect 34500 31132 34534 31424
rect 35558 31132 35592 31424
rect 36616 31132 36650 31424
rect 37674 31132 37708 31424
rect 38732 31132 38766 31424
rect 39790 31132 39824 31424
rect 40990 31132 41024 31424
rect 42048 31132 42082 31424
rect 43106 31132 43140 31424
rect 44164 31132 44198 31424
rect 45222 31132 45256 31424
rect 46280 31132 46314 31424
rect 47578 31154 47612 31446
rect 48636 31154 48670 31446
rect 49694 31154 49728 31446
rect 50752 31154 50786 31446
rect 51810 31154 51844 31446
rect 52868 31154 52902 31446
rect 54092 31168 54126 31460
rect 55150 31168 55184 31460
rect 56208 31168 56242 31460
rect 57266 31168 57300 31460
rect 58324 31168 58358 31460
rect 59382 31168 59416 31460
rect 1958 30016 1992 30308
rect 3016 30016 3050 30308
rect 4074 30016 4108 30308
rect 5132 30016 5166 30308
rect 6190 30016 6224 30308
rect 7248 30016 7282 30308
rect 1958 28922 1992 29214
rect 3016 28922 3050 29214
rect 4074 28922 4108 29214
rect 5132 28922 5166 29214
rect 6190 28922 6224 29214
rect 7248 28922 7282 29214
rect 8472 30024 8506 30316
rect 9530 30024 9564 30316
rect 10588 30024 10622 30316
rect 11646 30024 11680 30316
rect 12704 30024 12738 30316
rect 13762 30024 13796 30316
rect 1958 27828 1992 28120
rect 3016 27828 3050 28120
rect 4074 27828 4108 28120
rect 5132 27828 5166 28120
rect 6190 27828 6224 28120
rect 8472 28930 8506 29222
rect 9530 28930 9564 29222
rect 10588 28930 10622 29222
rect 11646 28930 11680 29222
rect 12704 28930 12738 29222
rect 13762 28930 13796 29222
rect 14978 30032 15012 30324
rect 16036 30032 16070 30324
rect 17094 30032 17128 30324
rect 18152 30032 18186 30324
rect 19210 30032 19244 30324
rect 20268 30032 20302 30324
rect 7248 27828 7282 28120
rect 8472 27836 8506 28128
rect 9530 27836 9564 28128
rect 10588 27836 10622 28128
rect 11646 27836 11680 28128
rect 12704 27836 12738 28128
rect 14978 28938 15012 29230
rect 16036 28938 16070 29230
rect 17094 28938 17128 29230
rect 18152 28938 18186 29230
rect 19210 28938 19244 29230
rect 20268 28938 20302 29230
rect 21468 30016 21502 30308
rect 22526 30016 22560 30308
rect 23584 30016 23618 30308
rect 24642 30016 24676 30308
rect 25700 30016 25734 30308
rect 26758 30016 26792 30308
rect 13762 27836 13796 28128
rect 14978 27844 15012 28136
rect 16036 27844 16070 28136
rect 17094 27844 17128 28136
rect 18152 27844 18186 28136
rect 19210 27844 19244 28136
rect 21468 28922 21502 29214
rect 22526 28922 22560 29214
rect 23584 28922 23618 29214
rect 24642 28922 24676 29214
rect 25700 28922 25734 29214
rect 26758 28922 26792 29214
rect 27990 30032 28024 30324
rect 29048 30032 29082 30324
rect 30106 30032 30140 30324
rect 31164 30032 31198 30324
rect 32222 30032 32256 30324
rect 33280 30032 33314 30324
rect 20268 27844 20302 28136
rect 21468 27828 21502 28120
rect 22526 27828 22560 28120
rect 23584 27828 23618 28120
rect 24642 27828 24676 28120
rect 25700 27828 25734 28120
rect 27990 28938 28024 29230
rect 29048 28938 29082 29230
rect 30106 28938 30140 29230
rect 31164 28938 31198 29230
rect 32222 28938 32256 29230
rect 33280 28938 33314 29230
rect 34500 30038 34534 30330
rect 35558 30038 35592 30330
rect 36616 30038 36650 30330
rect 37674 30038 37708 30330
rect 38732 30038 38766 30330
rect 39790 30038 39824 30330
rect 26758 27828 26792 28120
rect 27990 27844 28024 28136
rect 29048 27844 29082 28136
rect 30106 27844 30140 28136
rect 31164 27844 31198 28136
rect 32222 27844 32256 28136
rect 34500 28944 34534 29236
rect 35558 28944 35592 29236
rect 36616 28944 36650 29236
rect 37674 28944 37708 29236
rect 38732 28944 38766 29236
rect 39790 28944 39824 29236
rect 40990 30038 41024 30330
rect 42048 30038 42082 30330
rect 43106 30038 43140 30330
rect 44164 30038 44198 30330
rect 45222 30038 45256 30330
rect 46280 30038 46314 30330
rect 33280 27844 33314 28136
rect 34500 27850 34534 28142
rect 35558 27850 35592 28142
rect 36616 27850 36650 28142
rect 37674 27850 37708 28142
rect 38732 27850 38766 28142
rect 40990 28944 41024 29236
rect 42048 28944 42082 29236
rect 43106 28944 43140 29236
rect 44164 28944 44198 29236
rect 45222 28944 45256 29236
rect 46280 28944 46314 29236
rect 47578 30060 47612 30352
rect 48636 30060 48670 30352
rect 49694 30060 49728 30352
rect 50752 30060 50786 30352
rect 51810 30060 51844 30352
rect 52868 30060 52902 30352
rect 39790 27850 39824 28142
rect 40990 27850 41024 28142
rect 42048 27850 42082 28142
rect 43106 27850 43140 28142
rect 44164 27850 44198 28142
rect 45222 27850 45256 28142
rect 47578 28966 47612 29258
rect 48636 28966 48670 29258
rect 49694 28966 49728 29258
rect 50752 28966 50786 29258
rect 51810 28966 51844 29258
rect 52868 28966 52902 29258
rect 54092 30074 54126 30366
rect 55150 30074 55184 30366
rect 56208 30074 56242 30366
rect 57266 30074 57300 30366
rect 58324 30074 58358 30366
rect 59382 30074 59416 30366
rect 46280 27850 46314 28142
rect 47578 27872 47612 28164
rect 48636 27872 48670 28164
rect 49694 27872 49728 28164
rect 50752 27872 50786 28164
rect 51810 27872 51844 28164
rect 54092 28980 54126 29272
rect 55150 28980 55184 29272
rect 56208 28980 56242 29272
rect 57266 28980 57300 29272
rect 58324 28980 58358 29272
rect 59382 28980 59416 29272
rect 52868 27872 52902 28164
rect 54092 27886 54126 28178
rect 55150 27886 55184 28178
rect 56208 27886 56242 28178
rect 57266 27886 57300 28178
rect 58324 27886 58358 28178
rect 59382 27886 59416 28178
rect 1958 26734 1992 27026
rect 3016 26734 3050 27026
rect 4074 26734 4108 27026
rect 5132 26734 5166 27026
rect 6190 26734 6224 27026
rect 7248 26734 7282 27026
rect 8472 26742 8506 27034
rect 9530 26742 9564 27034
rect 10588 26742 10622 27034
rect 11646 26742 11680 27034
rect 12704 26742 12738 27034
rect 13762 26742 13796 27034
rect 14978 26750 15012 27042
rect 16036 26750 16070 27042
rect 17094 26750 17128 27042
rect 18152 26750 18186 27042
rect 19210 26750 19244 27042
rect 20268 26750 20302 27042
rect 21468 26734 21502 27026
rect 22526 26734 22560 27026
rect 23584 26734 23618 27026
rect 24642 26734 24676 27026
rect 25700 26734 25734 27026
rect 26758 26734 26792 27026
rect 27990 26750 28024 27042
rect 29048 26750 29082 27042
rect 30106 26750 30140 27042
rect 31164 26750 31198 27042
rect 32222 26750 32256 27042
rect 33280 26750 33314 27042
rect 34500 26756 34534 27048
rect 35558 26756 35592 27048
rect 36616 26756 36650 27048
rect 37674 26756 37708 27048
rect 38732 26756 38766 27048
rect 39790 26756 39824 27048
rect 40990 26756 41024 27048
rect 42048 26756 42082 27048
rect 43106 26756 43140 27048
rect 44164 26756 44198 27048
rect 45222 26756 45256 27048
rect 46280 26756 46314 27048
rect 47578 26778 47612 27070
rect 48636 26778 48670 27070
rect 49694 26778 49728 27070
rect 50752 26778 50786 27070
rect 51810 26778 51844 27070
rect 52868 26778 52902 27070
rect 54092 26792 54126 27084
rect 55150 26792 55184 27084
rect 56208 26792 56242 27084
rect 57266 26792 57300 27084
rect 58324 26792 58358 27084
rect 59382 26792 59416 27084
rect 1958 25274 1992 25566
rect 3016 25274 3050 25566
rect 4074 25274 4108 25566
rect 5132 25274 5166 25566
rect 6190 25274 6224 25566
rect 7248 25274 7282 25566
rect 8472 25282 8506 25574
rect 9530 25282 9564 25574
rect 10588 25282 10622 25574
rect 11646 25282 11680 25574
rect 12704 25282 12738 25574
rect 13762 25282 13796 25574
rect 14978 25290 15012 25582
rect 16036 25290 16070 25582
rect 17094 25290 17128 25582
rect 18152 25290 18186 25582
rect 19210 25290 19244 25582
rect 20268 25290 20302 25582
rect 21468 25274 21502 25566
rect 22526 25274 22560 25566
rect 23584 25274 23618 25566
rect 24642 25274 24676 25566
rect 25700 25274 25734 25566
rect 26758 25274 26792 25566
rect 27990 25290 28024 25582
rect 29048 25290 29082 25582
rect 30106 25290 30140 25582
rect 31164 25290 31198 25582
rect 32222 25290 32256 25582
rect 33280 25290 33314 25582
rect 34500 25296 34534 25588
rect 35558 25296 35592 25588
rect 36616 25296 36650 25588
rect 37674 25296 37708 25588
rect 38732 25296 38766 25588
rect 39790 25296 39824 25588
rect 40990 25296 41024 25588
rect 42048 25296 42082 25588
rect 43106 25296 43140 25588
rect 44164 25296 44198 25588
rect 45222 25296 45256 25588
rect 46280 25296 46314 25588
rect 47578 25318 47612 25610
rect 48636 25318 48670 25610
rect 49694 25318 49728 25610
rect 50752 25318 50786 25610
rect 51810 25318 51844 25610
rect 52868 25318 52902 25610
rect 54092 25332 54126 25624
rect 55150 25332 55184 25624
rect 56208 25332 56242 25624
rect 57266 25332 57300 25624
rect 58324 25332 58358 25624
rect 59382 25332 59416 25624
rect 1958 24180 1992 24472
rect 3016 24180 3050 24472
rect 4074 24180 4108 24472
rect 5132 24180 5166 24472
rect 6190 24180 6224 24472
rect 7248 24180 7282 24472
rect 1958 23086 1992 23378
rect 3016 23086 3050 23378
rect 4074 23086 4108 23378
rect 5132 23086 5166 23378
rect 6190 23086 6224 23378
rect 7248 23086 7282 23378
rect 8472 24188 8506 24480
rect 9530 24188 9564 24480
rect 10588 24188 10622 24480
rect 11646 24188 11680 24480
rect 12704 24188 12738 24480
rect 13762 24188 13796 24480
rect 1958 21992 1992 22284
rect 3016 21992 3050 22284
rect 4074 21992 4108 22284
rect 5132 21992 5166 22284
rect 6190 21992 6224 22284
rect 8472 23094 8506 23386
rect 9530 23094 9564 23386
rect 10588 23094 10622 23386
rect 11646 23094 11680 23386
rect 12704 23094 12738 23386
rect 13762 23094 13796 23386
rect 14978 24196 15012 24488
rect 16036 24196 16070 24488
rect 17094 24196 17128 24488
rect 18152 24196 18186 24488
rect 19210 24196 19244 24488
rect 20268 24196 20302 24488
rect 7248 21992 7282 22284
rect 8472 22000 8506 22292
rect 9530 22000 9564 22292
rect 10588 22000 10622 22292
rect 11646 22000 11680 22292
rect 12704 22000 12738 22292
rect 14978 23102 15012 23394
rect 16036 23102 16070 23394
rect 17094 23102 17128 23394
rect 18152 23102 18186 23394
rect 19210 23102 19244 23394
rect 20268 23102 20302 23394
rect 21468 24180 21502 24472
rect 22526 24180 22560 24472
rect 23584 24180 23618 24472
rect 24642 24180 24676 24472
rect 25700 24180 25734 24472
rect 26758 24180 26792 24472
rect 13762 22000 13796 22292
rect 14978 22008 15012 22300
rect 16036 22008 16070 22300
rect 17094 22008 17128 22300
rect 18152 22008 18186 22300
rect 19210 22008 19244 22300
rect 21468 23086 21502 23378
rect 22526 23086 22560 23378
rect 23584 23086 23618 23378
rect 24642 23086 24676 23378
rect 25700 23086 25734 23378
rect 26758 23086 26792 23378
rect 27990 24196 28024 24488
rect 29048 24196 29082 24488
rect 30106 24196 30140 24488
rect 31164 24196 31198 24488
rect 32222 24196 32256 24488
rect 33280 24196 33314 24488
rect 20268 22008 20302 22300
rect 21468 21992 21502 22284
rect 22526 21992 22560 22284
rect 23584 21992 23618 22284
rect 24642 21992 24676 22284
rect 25700 21992 25734 22284
rect 27990 23102 28024 23394
rect 29048 23102 29082 23394
rect 30106 23102 30140 23394
rect 31164 23102 31198 23394
rect 32222 23102 32256 23394
rect 33280 23102 33314 23394
rect 34500 24202 34534 24494
rect 35558 24202 35592 24494
rect 36616 24202 36650 24494
rect 37674 24202 37708 24494
rect 38732 24202 38766 24494
rect 39790 24202 39824 24494
rect 26758 21992 26792 22284
rect 27990 22008 28024 22300
rect 29048 22008 29082 22300
rect 30106 22008 30140 22300
rect 31164 22008 31198 22300
rect 32222 22008 32256 22300
rect 34500 23108 34534 23400
rect 35558 23108 35592 23400
rect 36616 23108 36650 23400
rect 37674 23108 37708 23400
rect 38732 23108 38766 23400
rect 39790 23108 39824 23400
rect 40990 24202 41024 24494
rect 42048 24202 42082 24494
rect 43106 24202 43140 24494
rect 44164 24202 44198 24494
rect 45222 24202 45256 24494
rect 46280 24202 46314 24494
rect 33280 22008 33314 22300
rect 34500 22014 34534 22306
rect 35558 22014 35592 22306
rect 36616 22014 36650 22306
rect 37674 22014 37708 22306
rect 38732 22014 38766 22306
rect 40990 23108 41024 23400
rect 42048 23108 42082 23400
rect 43106 23108 43140 23400
rect 44164 23108 44198 23400
rect 45222 23108 45256 23400
rect 46280 23108 46314 23400
rect 47578 24224 47612 24516
rect 48636 24224 48670 24516
rect 49694 24224 49728 24516
rect 50752 24224 50786 24516
rect 51810 24224 51844 24516
rect 52868 24224 52902 24516
rect 39790 22014 39824 22306
rect 40990 22014 41024 22306
rect 42048 22014 42082 22306
rect 43106 22014 43140 22306
rect 44164 22014 44198 22306
rect 45222 22014 45256 22306
rect 47578 23130 47612 23422
rect 48636 23130 48670 23422
rect 49694 23130 49728 23422
rect 50752 23130 50786 23422
rect 51810 23130 51844 23422
rect 52868 23130 52902 23422
rect 54092 24238 54126 24530
rect 55150 24238 55184 24530
rect 56208 24238 56242 24530
rect 57266 24238 57300 24530
rect 58324 24238 58358 24530
rect 59382 24238 59416 24530
rect 46280 22014 46314 22306
rect 47578 22036 47612 22328
rect 48636 22036 48670 22328
rect 49694 22036 49728 22328
rect 50752 22036 50786 22328
rect 51810 22036 51844 22328
rect 54092 23144 54126 23436
rect 55150 23144 55184 23436
rect 56208 23144 56242 23436
rect 57266 23144 57300 23436
rect 58324 23144 58358 23436
rect 59382 23144 59416 23436
rect 52868 22036 52902 22328
rect 54092 22050 54126 22342
rect 55150 22050 55184 22342
rect 56208 22050 56242 22342
rect 57266 22050 57300 22342
rect 58324 22050 58358 22342
rect 59382 22050 59416 22342
rect 1958 20898 1992 21190
rect 3016 20898 3050 21190
rect 4074 20898 4108 21190
rect 5132 20898 5166 21190
rect 6190 20898 6224 21190
rect 7248 20898 7282 21190
rect 8472 20906 8506 21198
rect 9530 20906 9564 21198
rect 10588 20906 10622 21198
rect 11646 20906 11680 21198
rect 12704 20906 12738 21198
rect 13762 20906 13796 21198
rect 14978 20914 15012 21206
rect 16036 20914 16070 21206
rect 17094 20914 17128 21206
rect 18152 20914 18186 21206
rect 19210 20914 19244 21206
rect 20268 20914 20302 21206
rect 21468 20898 21502 21190
rect 22526 20898 22560 21190
rect 23584 20898 23618 21190
rect 24642 20898 24676 21190
rect 25700 20898 25734 21190
rect 26758 20898 26792 21190
rect 27990 20914 28024 21206
rect 29048 20914 29082 21206
rect 30106 20914 30140 21206
rect 31164 20914 31198 21206
rect 32222 20914 32256 21206
rect 33280 20914 33314 21206
rect 34500 20920 34534 21212
rect 35558 20920 35592 21212
rect 36616 20920 36650 21212
rect 37674 20920 37708 21212
rect 38732 20920 38766 21212
rect 39790 20920 39824 21212
rect 40990 20920 41024 21212
rect 42048 20920 42082 21212
rect 43106 20920 43140 21212
rect 44164 20920 44198 21212
rect 45222 20920 45256 21212
rect 46280 20920 46314 21212
rect 47578 20942 47612 21234
rect 48636 20942 48670 21234
rect 49694 20942 49728 21234
rect 50752 20942 50786 21234
rect 51810 20942 51844 21234
rect 52868 20942 52902 21234
rect 54092 20956 54126 21248
rect 55150 20956 55184 21248
rect 56208 20956 56242 21248
rect 57266 20956 57300 21248
rect 58324 20956 58358 21248
rect 59382 20956 59416 21248
rect 1958 19410 1992 19702
rect 3016 19410 3050 19702
rect 4074 19410 4108 19702
rect 5132 19410 5166 19702
rect 6190 19410 6224 19702
rect 7248 19410 7282 19702
rect 8472 19418 8506 19710
rect 9530 19418 9564 19710
rect 10588 19418 10622 19710
rect 11646 19418 11680 19710
rect 12704 19418 12738 19710
rect 13762 19418 13796 19710
rect 14978 19426 15012 19718
rect 16036 19426 16070 19718
rect 17094 19426 17128 19718
rect 18152 19426 18186 19718
rect 19210 19426 19244 19718
rect 20268 19426 20302 19718
rect 21468 19410 21502 19702
rect 22526 19410 22560 19702
rect 23584 19410 23618 19702
rect 24642 19410 24676 19702
rect 25700 19410 25734 19702
rect 26758 19410 26792 19702
rect 27990 19426 28024 19718
rect 29048 19426 29082 19718
rect 30106 19426 30140 19718
rect 31164 19426 31198 19718
rect 32222 19426 32256 19718
rect 33280 19426 33314 19718
rect 34500 19432 34534 19724
rect 35558 19432 35592 19724
rect 36616 19432 36650 19724
rect 37674 19432 37708 19724
rect 38732 19432 38766 19724
rect 39790 19432 39824 19724
rect 40990 19432 41024 19724
rect 42048 19432 42082 19724
rect 43106 19432 43140 19724
rect 44164 19432 44198 19724
rect 45222 19432 45256 19724
rect 46280 19432 46314 19724
rect 47578 19454 47612 19746
rect 48636 19454 48670 19746
rect 49694 19454 49728 19746
rect 50752 19454 50786 19746
rect 51810 19454 51844 19746
rect 52868 19454 52902 19746
rect 54092 19468 54126 19760
rect 55150 19468 55184 19760
rect 56208 19468 56242 19760
rect 57266 19468 57300 19760
rect 58324 19468 58358 19760
rect 59382 19468 59416 19760
rect 1958 18316 1992 18608
rect 3016 18316 3050 18608
rect 4074 18316 4108 18608
rect 5132 18316 5166 18608
rect 6190 18316 6224 18608
rect 7248 18316 7282 18608
rect 1958 17222 1992 17514
rect 3016 17222 3050 17514
rect 4074 17222 4108 17514
rect 5132 17222 5166 17514
rect 6190 17222 6224 17514
rect 7248 17222 7282 17514
rect 8472 18324 8506 18616
rect 9530 18324 9564 18616
rect 10588 18324 10622 18616
rect 11646 18324 11680 18616
rect 12704 18324 12738 18616
rect 13762 18324 13796 18616
rect 1958 16128 1992 16420
rect 3016 16128 3050 16420
rect 4074 16128 4108 16420
rect 5132 16128 5166 16420
rect 6190 16128 6224 16420
rect 8472 17230 8506 17522
rect 9530 17230 9564 17522
rect 10588 17230 10622 17522
rect 11646 17230 11680 17522
rect 12704 17230 12738 17522
rect 13762 17230 13796 17522
rect 14978 18332 15012 18624
rect 16036 18332 16070 18624
rect 17094 18332 17128 18624
rect 18152 18332 18186 18624
rect 19210 18332 19244 18624
rect 20268 18332 20302 18624
rect 7248 16128 7282 16420
rect 8472 16136 8506 16428
rect 9530 16136 9564 16428
rect 10588 16136 10622 16428
rect 11646 16136 11680 16428
rect 12704 16136 12738 16428
rect 14978 17238 15012 17530
rect 16036 17238 16070 17530
rect 17094 17238 17128 17530
rect 18152 17238 18186 17530
rect 19210 17238 19244 17530
rect 20268 17238 20302 17530
rect 21468 18316 21502 18608
rect 22526 18316 22560 18608
rect 23584 18316 23618 18608
rect 24642 18316 24676 18608
rect 25700 18316 25734 18608
rect 26758 18316 26792 18608
rect 13762 16136 13796 16428
rect 14978 16144 15012 16436
rect 16036 16144 16070 16436
rect 17094 16144 17128 16436
rect 18152 16144 18186 16436
rect 19210 16144 19244 16436
rect 21468 17222 21502 17514
rect 22526 17222 22560 17514
rect 23584 17222 23618 17514
rect 24642 17222 24676 17514
rect 25700 17222 25734 17514
rect 26758 17222 26792 17514
rect 27990 18332 28024 18624
rect 29048 18332 29082 18624
rect 30106 18332 30140 18624
rect 31164 18332 31198 18624
rect 32222 18332 32256 18624
rect 33280 18332 33314 18624
rect 20268 16144 20302 16436
rect 21468 16128 21502 16420
rect 22526 16128 22560 16420
rect 23584 16128 23618 16420
rect 24642 16128 24676 16420
rect 25700 16128 25734 16420
rect 27990 17238 28024 17530
rect 29048 17238 29082 17530
rect 30106 17238 30140 17530
rect 31164 17238 31198 17530
rect 32222 17238 32256 17530
rect 33280 17238 33314 17530
rect 34500 18338 34534 18630
rect 35558 18338 35592 18630
rect 36616 18338 36650 18630
rect 37674 18338 37708 18630
rect 38732 18338 38766 18630
rect 39790 18338 39824 18630
rect 26758 16128 26792 16420
rect 27990 16144 28024 16436
rect 29048 16144 29082 16436
rect 30106 16144 30140 16436
rect 31164 16144 31198 16436
rect 32222 16144 32256 16436
rect 34500 17244 34534 17536
rect 35558 17244 35592 17536
rect 36616 17244 36650 17536
rect 37674 17244 37708 17536
rect 38732 17244 38766 17536
rect 39790 17244 39824 17536
rect 40990 18338 41024 18630
rect 42048 18338 42082 18630
rect 43106 18338 43140 18630
rect 44164 18338 44198 18630
rect 45222 18338 45256 18630
rect 46280 18338 46314 18630
rect 33280 16144 33314 16436
rect 34500 16150 34534 16442
rect 35558 16150 35592 16442
rect 36616 16150 36650 16442
rect 37674 16150 37708 16442
rect 38732 16150 38766 16442
rect 40990 17244 41024 17536
rect 42048 17244 42082 17536
rect 43106 17244 43140 17536
rect 44164 17244 44198 17536
rect 45222 17244 45256 17536
rect 46280 17244 46314 17536
rect 47578 18360 47612 18652
rect 48636 18360 48670 18652
rect 49694 18360 49728 18652
rect 50752 18360 50786 18652
rect 51810 18360 51844 18652
rect 52868 18360 52902 18652
rect 39790 16150 39824 16442
rect 40990 16150 41024 16442
rect 42048 16150 42082 16442
rect 43106 16150 43140 16442
rect 44164 16150 44198 16442
rect 45222 16150 45256 16442
rect 47578 17266 47612 17558
rect 48636 17266 48670 17558
rect 49694 17266 49728 17558
rect 50752 17266 50786 17558
rect 51810 17266 51844 17558
rect 52868 17266 52902 17558
rect 54092 18374 54126 18666
rect 55150 18374 55184 18666
rect 56208 18374 56242 18666
rect 57266 18374 57300 18666
rect 58324 18374 58358 18666
rect 59382 18374 59416 18666
rect 46280 16150 46314 16442
rect 47578 16172 47612 16464
rect 48636 16172 48670 16464
rect 49694 16172 49728 16464
rect 50752 16172 50786 16464
rect 51810 16172 51844 16464
rect 54092 17280 54126 17572
rect 55150 17280 55184 17572
rect 56208 17280 56242 17572
rect 57266 17280 57300 17572
rect 58324 17280 58358 17572
rect 59382 17280 59416 17572
rect 52868 16172 52902 16464
rect 54092 16186 54126 16478
rect 55150 16186 55184 16478
rect 56208 16186 56242 16478
rect 57266 16186 57300 16478
rect 58324 16186 58358 16478
rect 59382 16186 59416 16478
rect 1958 15034 1992 15326
rect 3016 15034 3050 15326
rect 4074 15034 4108 15326
rect 5132 15034 5166 15326
rect 6190 15034 6224 15326
rect 7248 15034 7282 15326
rect 8472 15042 8506 15334
rect 9530 15042 9564 15334
rect 10588 15042 10622 15334
rect 11646 15042 11680 15334
rect 12704 15042 12738 15334
rect 13762 15042 13796 15334
rect 14978 15050 15012 15342
rect 16036 15050 16070 15342
rect 17094 15050 17128 15342
rect 18152 15050 18186 15342
rect 19210 15050 19244 15342
rect 20268 15050 20302 15342
rect 21468 15034 21502 15326
rect 22526 15034 22560 15326
rect 23584 15034 23618 15326
rect 24642 15034 24676 15326
rect 25700 15034 25734 15326
rect 26758 15034 26792 15326
rect 27990 15050 28024 15342
rect 29048 15050 29082 15342
rect 30106 15050 30140 15342
rect 31164 15050 31198 15342
rect 32222 15050 32256 15342
rect 33280 15050 33314 15342
rect 34500 15056 34534 15348
rect 35558 15056 35592 15348
rect 36616 15056 36650 15348
rect 37674 15056 37708 15348
rect 38732 15056 38766 15348
rect 39790 15056 39824 15348
rect 40990 15056 41024 15348
rect 42048 15056 42082 15348
rect 43106 15056 43140 15348
rect 44164 15056 44198 15348
rect 45222 15056 45256 15348
rect 46280 15056 46314 15348
rect 47578 15078 47612 15370
rect 48636 15078 48670 15370
rect 49694 15078 49728 15370
rect 50752 15078 50786 15370
rect 51810 15078 51844 15370
rect 52868 15078 52902 15370
rect 54092 15092 54126 15384
rect 55150 15092 55184 15384
rect 56208 15092 56242 15384
rect 57266 15092 57300 15384
rect 58324 15092 58358 15384
rect 59382 15092 59416 15384
rect 1968 13554 2002 13846
rect 3026 13554 3060 13846
rect 4084 13554 4118 13846
rect 5142 13554 5176 13846
rect 6200 13554 6234 13846
rect 7258 13554 7292 13846
rect 8482 13562 8516 13854
rect 9540 13562 9574 13854
rect 10598 13562 10632 13854
rect 11656 13562 11690 13854
rect 12714 13562 12748 13854
rect 13772 13562 13806 13854
rect 14988 13570 15022 13862
rect 16046 13570 16080 13862
rect 17104 13570 17138 13862
rect 18162 13570 18196 13862
rect 19220 13570 19254 13862
rect 20278 13570 20312 13862
rect 21478 13554 21512 13846
rect 22536 13554 22570 13846
rect 23594 13554 23628 13846
rect 24652 13554 24686 13846
rect 25710 13554 25744 13846
rect 26768 13554 26802 13846
rect 28000 13570 28034 13862
rect 29058 13570 29092 13862
rect 30116 13570 30150 13862
rect 31174 13570 31208 13862
rect 32232 13570 32266 13862
rect 33290 13570 33324 13862
rect 34510 13576 34544 13868
rect 35568 13576 35602 13868
rect 36626 13576 36660 13868
rect 37684 13576 37718 13868
rect 38742 13576 38776 13868
rect 39800 13576 39834 13868
rect 41000 13576 41034 13868
rect 42058 13576 42092 13868
rect 43116 13576 43150 13868
rect 44174 13576 44208 13868
rect 45232 13576 45266 13868
rect 46290 13576 46324 13868
rect 47588 13598 47622 13890
rect 48646 13598 48680 13890
rect 49704 13598 49738 13890
rect 50762 13598 50796 13890
rect 51820 13598 51854 13890
rect 52878 13598 52912 13890
rect 54102 13612 54136 13904
rect 55160 13612 55194 13904
rect 56218 13612 56252 13904
rect 57276 13612 57310 13904
rect 58334 13612 58368 13904
rect 59392 13612 59426 13904
rect 1968 12460 2002 12752
rect 3026 12460 3060 12752
rect 4084 12460 4118 12752
rect 5142 12460 5176 12752
rect 6200 12460 6234 12752
rect 7258 12460 7292 12752
rect 1968 11366 2002 11658
rect 3026 11366 3060 11658
rect 4084 11366 4118 11658
rect 5142 11366 5176 11658
rect 6200 11366 6234 11658
rect 7258 11366 7292 11658
rect 8482 12468 8516 12760
rect 9540 12468 9574 12760
rect 10598 12468 10632 12760
rect 11656 12468 11690 12760
rect 12714 12468 12748 12760
rect 13772 12468 13806 12760
rect 1968 10272 2002 10564
rect 3026 10272 3060 10564
rect 4084 10272 4118 10564
rect 5142 10272 5176 10564
rect 6200 10272 6234 10564
rect 8482 11374 8516 11666
rect 9540 11374 9574 11666
rect 10598 11374 10632 11666
rect 11656 11374 11690 11666
rect 12714 11374 12748 11666
rect 13772 11374 13806 11666
rect 14988 12476 15022 12768
rect 16046 12476 16080 12768
rect 17104 12476 17138 12768
rect 18162 12476 18196 12768
rect 19220 12476 19254 12768
rect 20278 12476 20312 12768
rect 7258 10272 7292 10564
rect 8482 10280 8516 10572
rect 9540 10280 9574 10572
rect 10598 10280 10632 10572
rect 11656 10280 11690 10572
rect 12714 10280 12748 10572
rect 14988 11382 15022 11674
rect 16046 11382 16080 11674
rect 17104 11382 17138 11674
rect 18162 11382 18196 11674
rect 19220 11382 19254 11674
rect 20278 11382 20312 11674
rect 21478 12460 21512 12752
rect 22536 12460 22570 12752
rect 23594 12460 23628 12752
rect 24652 12460 24686 12752
rect 25710 12460 25744 12752
rect 26768 12460 26802 12752
rect 13772 10280 13806 10572
rect 14988 10288 15022 10580
rect 16046 10288 16080 10580
rect 17104 10288 17138 10580
rect 18162 10288 18196 10580
rect 19220 10288 19254 10580
rect 21478 11366 21512 11658
rect 22536 11366 22570 11658
rect 23594 11366 23628 11658
rect 24652 11366 24686 11658
rect 25710 11366 25744 11658
rect 26768 11366 26802 11658
rect 28000 12476 28034 12768
rect 29058 12476 29092 12768
rect 30116 12476 30150 12768
rect 31174 12476 31208 12768
rect 32232 12476 32266 12768
rect 33290 12476 33324 12768
rect 20278 10288 20312 10580
rect 21478 10272 21512 10564
rect 22536 10272 22570 10564
rect 23594 10272 23628 10564
rect 24652 10272 24686 10564
rect 25710 10272 25744 10564
rect 28000 11382 28034 11674
rect 29058 11382 29092 11674
rect 30116 11382 30150 11674
rect 31174 11382 31208 11674
rect 32232 11382 32266 11674
rect 33290 11382 33324 11674
rect 34510 12482 34544 12774
rect 35568 12482 35602 12774
rect 36626 12482 36660 12774
rect 37684 12482 37718 12774
rect 38742 12482 38776 12774
rect 39800 12482 39834 12774
rect 26768 10272 26802 10564
rect 28000 10288 28034 10580
rect 29058 10288 29092 10580
rect 30116 10288 30150 10580
rect 31174 10288 31208 10580
rect 32232 10288 32266 10580
rect 34510 11388 34544 11680
rect 35568 11388 35602 11680
rect 36626 11388 36660 11680
rect 37684 11388 37718 11680
rect 38742 11388 38776 11680
rect 39800 11388 39834 11680
rect 41000 12482 41034 12774
rect 42058 12482 42092 12774
rect 43116 12482 43150 12774
rect 44174 12482 44208 12774
rect 45232 12482 45266 12774
rect 46290 12482 46324 12774
rect 33290 10288 33324 10580
rect 34510 10294 34544 10586
rect 35568 10294 35602 10586
rect 36626 10294 36660 10586
rect 37684 10294 37718 10586
rect 38742 10294 38776 10586
rect 41000 11388 41034 11680
rect 42058 11388 42092 11680
rect 43116 11388 43150 11680
rect 44174 11388 44208 11680
rect 45232 11388 45266 11680
rect 46290 11388 46324 11680
rect 47588 12504 47622 12796
rect 48646 12504 48680 12796
rect 49704 12504 49738 12796
rect 50762 12504 50796 12796
rect 51820 12504 51854 12796
rect 52878 12504 52912 12796
rect 39800 10294 39834 10586
rect 41000 10294 41034 10586
rect 42058 10294 42092 10586
rect 43116 10294 43150 10586
rect 44174 10294 44208 10586
rect 45232 10294 45266 10586
rect 47588 11410 47622 11702
rect 48646 11410 48680 11702
rect 49704 11410 49738 11702
rect 50762 11410 50796 11702
rect 51820 11410 51854 11702
rect 52878 11410 52912 11702
rect 54102 12518 54136 12810
rect 55160 12518 55194 12810
rect 56218 12518 56252 12810
rect 57276 12518 57310 12810
rect 58334 12518 58368 12810
rect 59392 12518 59426 12810
rect 46290 10294 46324 10586
rect 47588 10316 47622 10608
rect 48646 10316 48680 10608
rect 49704 10316 49738 10608
rect 50762 10316 50796 10608
rect 51820 10316 51854 10608
rect 54102 11424 54136 11716
rect 55160 11424 55194 11716
rect 56218 11424 56252 11716
rect 57276 11424 57310 11716
rect 58334 11424 58368 11716
rect 59392 11424 59426 11716
rect 52878 10316 52912 10608
rect 54102 10330 54136 10622
rect 55160 10330 55194 10622
rect 56218 10330 56252 10622
rect 57276 10330 57310 10622
rect 58334 10330 58368 10622
rect 59392 10330 59426 10622
rect 1968 9178 2002 9470
rect 3026 9178 3060 9470
rect 4084 9178 4118 9470
rect 5142 9178 5176 9470
rect 6200 9178 6234 9470
rect 7258 9178 7292 9470
rect 8482 9186 8516 9478
rect 9540 9186 9574 9478
rect 10598 9186 10632 9478
rect 11656 9186 11690 9478
rect 12714 9186 12748 9478
rect 13772 9186 13806 9478
rect 14988 9194 15022 9486
rect 16046 9194 16080 9486
rect 17104 9194 17138 9486
rect 18162 9194 18196 9486
rect 19220 9194 19254 9486
rect 20278 9194 20312 9486
rect 21478 9178 21512 9470
rect 22536 9178 22570 9470
rect 23594 9178 23628 9470
rect 24652 9178 24686 9470
rect 25710 9178 25744 9470
rect 26768 9178 26802 9470
rect 28000 9194 28034 9486
rect 29058 9194 29092 9486
rect 30116 9194 30150 9486
rect 31174 9194 31208 9486
rect 32232 9194 32266 9486
rect 33290 9194 33324 9486
rect 34510 9200 34544 9492
rect 35568 9200 35602 9492
rect 36626 9200 36660 9492
rect 37684 9200 37718 9492
rect 38742 9200 38776 9492
rect 39800 9200 39834 9492
rect 41000 9200 41034 9492
rect 42058 9200 42092 9492
rect 43116 9200 43150 9492
rect 44174 9200 44208 9492
rect 45232 9200 45266 9492
rect 46290 9200 46324 9492
rect 47588 9222 47622 9514
rect 48646 9222 48680 9514
rect 49704 9222 49738 9514
rect 50762 9222 50796 9514
rect 51820 9222 51854 9514
rect 52878 9222 52912 9514
rect 54102 9236 54136 9528
rect 55160 9236 55194 9528
rect 56218 9236 56252 9528
rect 57276 9236 57310 9528
rect 58334 9236 58368 9528
rect 59392 9236 59426 9528
rect 1986 7646 2020 7938
rect 3044 7646 3078 7938
rect 4102 7646 4136 7938
rect 5160 7646 5194 7938
rect 6218 7646 6252 7938
rect 7276 7646 7310 7938
rect 8500 7654 8534 7946
rect 9558 7654 9592 7946
rect 10616 7654 10650 7946
rect 11674 7654 11708 7946
rect 12732 7654 12766 7946
rect 13790 7654 13824 7946
rect 15006 7662 15040 7954
rect 16064 7662 16098 7954
rect 17122 7662 17156 7954
rect 18180 7662 18214 7954
rect 19238 7662 19272 7954
rect 20296 7662 20330 7954
rect 21496 7646 21530 7938
rect 22554 7646 22588 7938
rect 23612 7646 23646 7938
rect 24670 7646 24704 7938
rect 25728 7646 25762 7938
rect 26786 7646 26820 7938
rect 28018 7662 28052 7954
rect 29076 7662 29110 7954
rect 30134 7662 30168 7954
rect 31192 7662 31226 7954
rect 32250 7662 32284 7954
rect 33308 7662 33342 7954
rect 34528 7668 34562 7960
rect 35586 7668 35620 7960
rect 36644 7668 36678 7960
rect 37702 7668 37736 7960
rect 38760 7668 38794 7960
rect 39818 7668 39852 7960
rect 41018 7668 41052 7960
rect 42076 7668 42110 7960
rect 43134 7668 43168 7960
rect 44192 7668 44226 7960
rect 45250 7668 45284 7960
rect 46308 7668 46342 7960
rect 47606 7690 47640 7982
rect 48664 7690 48698 7982
rect 49722 7690 49756 7982
rect 50780 7690 50814 7982
rect 51838 7690 51872 7982
rect 52896 7690 52930 7982
rect 54120 7704 54154 7996
rect 55178 7704 55212 7996
rect 56236 7704 56270 7996
rect 57294 7704 57328 7996
rect 58352 7704 58386 7996
rect 59410 7704 59444 7996
rect 1986 6552 2020 6844
rect 3044 6552 3078 6844
rect 4102 6552 4136 6844
rect 5160 6552 5194 6844
rect 6218 6552 6252 6844
rect 7276 6552 7310 6844
rect 1986 5458 2020 5750
rect 3044 5458 3078 5750
rect 4102 5458 4136 5750
rect 5160 5458 5194 5750
rect 6218 5458 6252 5750
rect 7276 5458 7310 5750
rect 8500 6560 8534 6852
rect 9558 6560 9592 6852
rect 10616 6560 10650 6852
rect 11674 6560 11708 6852
rect 12732 6560 12766 6852
rect 13790 6560 13824 6852
rect 1986 4364 2020 4656
rect 3044 4364 3078 4656
rect 4102 4364 4136 4656
rect 5160 4364 5194 4656
rect 6218 4364 6252 4656
rect 8500 5466 8534 5758
rect 9558 5466 9592 5758
rect 10616 5466 10650 5758
rect 11674 5466 11708 5758
rect 12732 5466 12766 5758
rect 13790 5466 13824 5758
rect 15006 6568 15040 6860
rect 16064 6568 16098 6860
rect 17122 6568 17156 6860
rect 18180 6568 18214 6860
rect 19238 6568 19272 6860
rect 20296 6568 20330 6860
rect 7276 4364 7310 4656
rect 8500 4372 8534 4664
rect 9558 4372 9592 4664
rect 10616 4372 10650 4664
rect 11674 4372 11708 4664
rect 12732 4372 12766 4664
rect 15006 5474 15040 5766
rect 16064 5474 16098 5766
rect 17122 5474 17156 5766
rect 18180 5474 18214 5766
rect 19238 5474 19272 5766
rect 20296 5474 20330 5766
rect 21496 6552 21530 6844
rect 22554 6552 22588 6844
rect 23612 6552 23646 6844
rect 24670 6552 24704 6844
rect 25728 6552 25762 6844
rect 26786 6552 26820 6844
rect 13790 4372 13824 4664
rect 15006 4380 15040 4672
rect 16064 4380 16098 4672
rect 17122 4380 17156 4672
rect 18180 4380 18214 4672
rect 19238 4380 19272 4672
rect 21496 5458 21530 5750
rect 22554 5458 22588 5750
rect 23612 5458 23646 5750
rect 24670 5458 24704 5750
rect 25728 5458 25762 5750
rect 26786 5458 26820 5750
rect 28018 6568 28052 6860
rect 29076 6568 29110 6860
rect 30134 6568 30168 6860
rect 31192 6568 31226 6860
rect 32250 6568 32284 6860
rect 33308 6568 33342 6860
rect 20296 4380 20330 4672
rect 21496 4364 21530 4656
rect 22554 4364 22588 4656
rect 23612 4364 23646 4656
rect 24670 4364 24704 4656
rect 25728 4364 25762 4656
rect 28018 5474 28052 5766
rect 29076 5474 29110 5766
rect 30134 5474 30168 5766
rect 31192 5474 31226 5766
rect 32250 5474 32284 5766
rect 33308 5474 33342 5766
rect 34528 6574 34562 6866
rect 35586 6574 35620 6866
rect 36644 6574 36678 6866
rect 37702 6574 37736 6866
rect 38760 6574 38794 6866
rect 39818 6574 39852 6866
rect 26786 4364 26820 4656
rect 28018 4380 28052 4672
rect 29076 4380 29110 4672
rect 30134 4380 30168 4672
rect 31192 4380 31226 4672
rect 32250 4380 32284 4672
rect 34528 5480 34562 5772
rect 35586 5480 35620 5772
rect 36644 5480 36678 5772
rect 37702 5480 37736 5772
rect 38760 5480 38794 5772
rect 39818 5480 39852 5772
rect 41018 6574 41052 6866
rect 42076 6574 42110 6866
rect 43134 6574 43168 6866
rect 44192 6574 44226 6866
rect 45250 6574 45284 6866
rect 46308 6574 46342 6866
rect 33308 4380 33342 4672
rect 34528 4386 34562 4678
rect 35586 4386 35620 4678
rect 36644 4386 36678 4678
rect 37702 4386 37736 4678
rect 38760 4386 38794 4678
rect 41018 5480 41052 5772
rect 42076 5480 42110 5772
rect 43134 5480 43168 5772
rect 44192 5480 44226 5772
rect 45250 5480 45284 5772
rect 46308 5480 46342 5772
rect 47606 6596 47640 6888
rect 48664 6596 48698 6888
rect 49722 6596 49756 6888
rect 50780 6596 50814 6888
rect 51838 6596 51872 6888
rect 52896 6596 52930 6888
rect 39818 4386 39852 4678
rect 41018 4386 41052 4678
rect 42076 4386 42110 4678
rect 43134 4386 43168 4678
rect 44192 4386 44226 4678
rect 45250 4386 45284 4678
rect 47606 5502 47640 5794
rect 48664 5502 48698 5794
rect 49722 5502 49756 5794
rect 50780 5502 50814 5794
rect 51838 5502 51872 5794
rect 52896 5502 52930 5794
rect 54120 6610 54154 6902
rect 55178 6610 55212 6902
rect 56236 6610 56270 6902
rect 57294 6610 57328 6902
rect 58352 6610 58386 6902
rect 59410 6610 59444 6902
rect 46308 4386 46342 4678
rect 47606 4408 47640 4700
rect 48664 4408 48698 4700
rect 49722 4408 49756 4700
rect 50780 4408 50814 4700
rect 51838 4408 51872 4700
rect 54120 5516 54154 5808
rect 55178 5516 55212 5808
rect 56236 5516 56270 5808
rect 57294 5516 57328 5808
rect 58352 5516 58386 5808
rect 59410 5516 59444 5808
rect 52896 4408 52930 4700
rect 54120 4422 54154 4714
rect 55178 4422 55212 4714
rect 56236 4422 56270 4714
rect 57294 4422 57328 4714
rect 58352 4422 58386 4714
rect 59410 4422 59444 4714
rect 1986 3270 2020 3562
rect 3044 3270 3078 3562
rect 4102 3270 4136 3562
rect 5160 3270 5194 3562
rect 6218 3270 6252 3562
rect 7276 3270 7310 3562
rect 8500 3278 8534 3570
rect 9558 3278 9592 3570
rect 10616 3278 10650 3570
rect 11674 3278 11708 3570
rect 12732 3278 12766 3570
rect 13790 3278 13824 3570
rect 15006 3286 15040 3578
rect 16064 3286 16098 3578
rect 17122 3286 17156 3578
rect 18180 3286 18214 3578
rect 19238 3286 19272 3578
rect 20296 3286 20330 3578
rect 21496 3270 21530 3562
rect 22554 3270 22588 3562
rect 23612 3270 23646 3562
rect 24670 3270 24704 3562
rect 25728 3270 25762 3562
rect 26786 3270 26820 3562
rect 28018 3286 28052 3578
rect 29076 3286 29110 3578
rect 30134 3286 30168 3578
rect 31192 3286 31226 3578
rect 32250 3286 32284 3578
rect 33308 3286 33342 3578
rect 34528 3292 34562 3584
rect 35586 3292 35620 3584
rect 36644 3292 36678 3584
rect 37702 3292 37736 3584
rect 38760 3292 38794 3584
rect 39818 3292 39852 3584
rect 41018 3292 41052 3584
rect 42076 3292 42110 3584
rect 43134 3292 43168 3584
rect 44192 3292 44226 3584
rect 45250 3292 45284 3584
rect 46308 3292 46342 3584
rect 47606 3314 47640 3606
rect 48664 3314 48698 3606
rect 49722 3314 49756 3606
rect 50780 3314 50814 3606
rect 51838 3314 51872 3606
rect 52896 3314 52930 3606
rect 54120 3328 54154 3620
rect 55178 3328 55212 3620
rect 56236 3328 56270 3620
rect 57294 3328 57328 3620
rect 58352 3328 58386 3620
rect 59410 3328 59444 3620
rect 62112 25276 62146 25568
rect 63170 25276 63204 25568
rect 64228 25276 64262 25568
rect 65286 25276 65320 25568
rect 66344 25276 66378 25568
rect 67402 25276 67436 25568
rect 68574 25274 68608 25566
rect 69632 25274 69666 25566
rect 70690 25274 70724 25566
rect 71748 25274 71782 25566
rect 72806 25274 72840 25566
rect 73864 25274 73898 25566
rect 75268 25248 75302 25540
rect 76326 25248 76360 25540
rect 77384 25248 77418 25540
rect 78442 25248 78476 25540
rect 79500 25248 79534 25540
rect 80558 25248 80592 25540
rect 81730 25246 81764 25538
rect 82788 25246 82822 25538
rect 83846 25246 83880 25538
rect 84904 25246 84938 25538
rect 85962 25246 85996 25538
rect 87020 25246 87054 25538
rect 88502 25240 88536 25532
rect 62112 24182 62146 24474
rect 63170 24182 63204 24474
rect 64228 24182 64262 24474
rect 65286 24182 65320 24474
rect 66344 24182 66378 24474
rect 89560 25240 89594 25532
rect 90618 25240 90652 25532
rect 91676 25240 91710 25532
rect 92734 25240 92768 25532
rect 93792 25240 93826 25532
rect 94964 25238 94998 25530
rect 67402 24182 67436 24474
rect 62112 23088 62146 23380
rect 63170 23088 63204 23380
rect 64228 23088 64262 23380
rect 65286 23088 65320 23380
rect 66344 23088 66378 23380
rect 67402 23088 67436 23380
rect 68574 24180 68608 24472
rect 69632 24180 69666 24472
rect 70690 24180 70724 24472
rect 71748 24180 71782 24472
rect 72806 24180 72840 24472
rect 96022 25238 96056 25530
rect 97080 25238 97114 25530
rect 98138 25238 98172 25530
rect 99196 25238 99230 25530
rect 100254 25238 100288 25530
rect 73864 24180 73898 24472
rect 62112 21994 62146 22286
rect 63170 21994 63204 22286
rect 64228 21994 64262 22286
rect 65286 21994 65320 22286
rect 66344 21994 66378 22286
rect 68574 23086 68608 23378
rect 69632 23086 69666 23378
rect 70690 23086 70724 23378
rect 71748 23086 71782 23378
rect 72806 23086 72840 23378
rect 73864 23086 73898 23378
rect 75268 24154 75302 24446
rect 76326 24154 76360 24446
rect 77384 24154 77418 24446
rect 78442 24154 78476 24446
rect 79500 24154 79534 24446
rect 80558 24154 80592 24446
rect 67402 21994 67436 22286
rect 68574 21992 68608 22284
rect 69632 21992 69666 22284
rect 70690 21992 70724 22284
rect 71748 21992 71782 22284
rect 72806 21992 72840 22284
rect 75268 23060 75302 23352
rect 76326 23060 76360 23352
rect 77384 23060 77418 23352
rect 78442 23060 78476 23352
rect 79500 23060 79534 23352
rect 80558 23060 80592 23352
rect 81730 24152 81764 24444
rect 82788 24152 82822 24444
rect 83846 24152 83880 24444
rect 84904 24152 84938 24444
rect 85962 24152 85996 24444
rect 87020 24152 87054 24444
rect 73864 21992 73898 22284
rect 75268 21966 75302 22258
rect 76326 21966 76360 22258
rect 77384 21966 77418 22258
rect 78442 21966 78476 22258
rect 79500 21966 79534 22258
rect 81730 23058 81764 23350
rect 82788 23058 82822 23350
rect 83846 23058 83880 23350
rect 84904 23058 84938 23350
rect 85962 23058 85996 23350
rect 87020 23058 87054 23350
rect 88502 24146 88536 24438
rect 89560 24146 89594 24438
rect 90618 24146 90652 24438
rect 91676 24146 91710 24438
rect 92734 24146 92768 24438
rect 93792 24146 93826 24438
rect 80558 21966 80592 22258
rect 81730 21964 81764 22256
rect 82788 21964 82822 22256
rect 83846 21964 83880 22256
rect 84904 21964 84938 22256
rect 85962 21964 85996 22256
rect 88502 23052 88536 23344
rect 89560 23052 89594 23344
rect 90618 23052 90652 23344
rect 91676 23052 91710 23344
rect 92734 23052 92768 23344
rect 93792 23052 93826 23344
rect 94964 24144 94998 24436
rect 96022 24144 96056 24436
rect 97080 24144 97114 24436
rect 98138 24144 98172 24436
rect 99196 24144 99230 24436
rect 100254 24144 100288 24436
rect 87020 21964 87054 22256
rect 88502 21958 88536 22250
rect 62112 20900 62146 21192
rect 63170 20900 63204 21192
rect 64228 20900 64262 21192
rect 65286 20900 65320 21192
rect 66344 20900 66378 21192
rect 89560 21958 89594 22250
rect 90618 21958 90652 22250
rect 91676 21958 91710 22250
rect 92734 21958 92768 22250
rect 94964 23050 94998 23342
rect 96022 23050 96056 23342
rect 97080 23050 97114 23342
rect 98138 23050 98172 23342
rect 99196 23050 99230 23342
rect 100254 23050 100288 23342
rect 93792 21958 93826 22250
rect 94964 21956 94998 22248
rect 67402 20900 67436 21192
rect 68574 20898 68608 21190
rect 69632 20898 69666 21190
rect 70690 20898 70724 21190
rect 71748 20898 71782 21190
rect 72806 20898 72840 21190
rect 96022 21956 96056 22248
rect 97080 21956 97114 22248
rect 98138 21956 98172 22248
rect 99196 21956 99230 22248
rect 100254 21956 100288 22248
rect 73864 20898 73898 21190
rect 75268 20872 75302 21164
rect 76326 20872 76360 21164
rect 77384 20872 77418 21164
rect 78442 20872 78476 21164
rect 79500 20872 79534 21164
rect 80558 20872 80592 21164
rect 81730 20870 81764 21162
rect 82788 20870 82822 21162
rect 83846 20870 83880 21162
rect 84904 20870 84938 21162
rect 85962 20870 85996 21162
rect 87020 20870 87054 21162
rect 88502 20864 88536 21156
rect 89560 20864 89594 21156
rect 90618 20864 90652 21156
rect 91676 20864 91710 21156
rect 92734 20864 92768 21156
rect 93792 20864 93826 21156
rect 94964 20862 94998 21154
rect 96022 20862 96056 21154
rect 97080 20862 97114 21154
rect 98138 20862 98172 21154
rect 99196 20862 99230 21154
rect 100254 20862 100288 21154
rect 62118 19438 62152 19730
rect 63176 19438 63210 19730
rect 64234 19438 64268 19730
rect 65292 19438 65326 19730
rect 66350 19438 66384 19730
rect 67408 19438 67442 19730
rect 68582 19450 68616 19742
rect 69640 19450 69674 19742
rect 70698 19450 70732 19742
rect 71756 19450 71790 19742
rect 72814 19450 72848 19742
rect 73872 19450 73906 19742
rect 75274 19410 75308 19702
rect 76332 19410 76366 19702
rect 77390 19410 77424 19702
rect 78448 19410 78482 19702
rect 79506 19410 79540 19702
rect 80564 19410 80598 19702
rect 81738 19422 81772 19714
rect 82796 19422 82830 19714
rect 83854 19422 83888 19714
rect 84912 19422 84946 19714
rect 85970 19422 86004 19714
rect 87028 19422 87062 19714
rect 88508 19402 88542 19694
rect 89566 19402 89600 19694
rect 90624 19402 90658 19694
rect 91682 19402 91716 19694
rect 92740 19402 92774 19694
rect 93798 19402 93832 19694
rect 94972 19414 95006 19706
rect 96030 19414 96064 19706
rect 97088 19414 97122 19706
rect 98146 19414 98180 19706
rect 99204 19414 99238 19706
rect 100262 19414 100296 19706
rect 62118 18344 62152 18636
rect 63176 18344 63210 18636
rect 64234 18344 64268 18636
rect 65292 18344 65326 18636
rect 66350 18344 66384 18636
rect 67408 18344 67442 18636
rect 62118 17250 62152 17542
rect 63176 17250 63210 17542
rect 64234 17250 64268 17542
rect 65292 17250 65326 17542
rect 66350 17250 66384 17542
rect 67408 17250 67442 17542
rect 68582 18356 68616 18648
rect 69640 18356 69674 18648
rect 70698 18356 70732 18648
rect 71756 18356 71790 18648
rect 72814 18356 72848 18648
rect 73872 18356 73906 18648
rect 62118 16156 62152 16448
rect 63176 16156 63210 16448
rect 64234 16156 64268 16448
rect 65292 16156 65326 16448
rect 66350 16156 66384 16448
rect 68582 17262 68616 17554
rect 69640 17262 69674 17554
rect 70698 17262 70732 17554
rect 71756 17262 71790 17554
rect 72814 17262 72848 17554
rect 73872 17262 73906 17554
rect 75274 18316 75308 18608
rect 76332 18316 76366 18608
rect 77390 18316 77424 18608
rect 78448 18316 78482 18608
rect 79506 18316 79540 18608
rect 80564 18316 80598 18608
rect 67408 16156 67442 16448
rect 68582 16168 68616 16460
rect 69640 16168 69674 16460
rect 70698 16168 70732 16460
rect 71756 16168 71790 16460
rect 72814 16168 72848 16460
rect 75274 17222 75308 17514
rect 76332 17222 76366 17514
rect 77390 17222 77424 17514
rect 78448 17222 78482 17514
rect 79506 17222 79540 17514
rect 80564 17222 80598 17514
rect 81738 18328 81772 18620
rect 82796 18328 82830 18620
rect 83854 18328 83888 18620
rect 84912 18328 84946 18620
rect 85970 18328 86004 18620
rect 87028 18328 87062 18620
rect 73872 16168 73906 16460
rect 75274 16128 75308 16420
rect 76332 16128 76366 16420
rect 77390 16128 77424 16420
rect 78448 16128 78482 16420
rect 79506 16128 79540 16420
rect 81738 17234 81772 17526
rect 82796 17234 82830 17526
rect 83854 17234 83888 17526
rect 84912 17234 84946 17526
rect 85970 17234 86004 17526
rect 87028 17234 87062 17526
rect 88508 18308 88542 18600
rect 89566 18308 89600 18600
rect 90624 18308 90658 18600
rect 91682 18308 91716 18600
rect 92740 18308 92774 18600
rect 93798 18308 93832 18600
rect 80564 16128 80598 16420
rect 81738 16140 81772 16432
rect 82796 16140 82830 16432
rect 83854 16140 83888 16432
rect 84912 16140 84946 16432
rect 85970 16140 86004 16432
rect 88508 17214 88542 17506
rect 89566 17214 89600 17506
rect 90624 17214 90658 17506
rect 91682 17214 91716 17506
rect 92740 17214 92774 17506
rect 93798 17214 93832 17506
rect 94972 18320 95006 18612
rect 96030 18320 96064 18612
rect 97088 18320 97122 18612
rect 98146 18320 98180 18612
rect 99204 18320 99238 18612
rect 100262 18320 100296 18612
rect 87028 16140 87062 16432
rect 88508 16120 88542 16412
rect 89566 16120 89600 16412
rect 90624 16120 90658 16412
rect 91682 16120 91716 16412
rect 92740 16120 92774 16412
rect 94972 17226 95006 17518
rect 96030 17226 96064 17518
rect 97088 17226 97122 17518
rect 98146 17226 98180 17518
rect 99204 17226 99238 17518
rect 100262 17226 100296 17518
rect 93798 16120 93832 16412
rect 94972 16132 95006 16424
rect 96030 16132 96064 16424
rect 97088 16132 97122 16424
rect 98146 16132 98180 16424
rect 99204 16132 99238 16424
rect 100262 16132 100296 16424
rect 62118 15062 62152 15354
rect 63176 15062 63210 15354
rect 64234 15062 64268 15354
rect 65292 15062 65326 15354
rect 66350 15062 66384 15354
rect 67408 15062 67442 15354
rect 68582 15074 68616 15366
rect 69640 15074 69674 15366
rect 70698 15074 70732 15366
rect 71756 15074 71790 15366
rect 72814 15074 72848 15366
rect 73872 15074 73906 15366
rect 75274 15034 75308 15326
rect 76332 15034 76366 15326
rect 77390 15034 77424 15326
rect 78448 15034 78482 15326
rect 79506 15034 79540 15326
rect 80564 15034 80598 15326
rect 81738 15046 81772 15338
rect 82796 15046 82830 15338
rect 83854 15046 83888 15338
rect 84912 15046 84946 15338
rect 85970 15046 86004 15338
rect 87028 15046 87062 15338
rect 88508 15026 88542 15318
rect 89566 15026 89600 15318
rect 90624 15026 90658 15318
rect 91682 15026 91716 15318
rect 92740 15026 92774 15318
rect 93798 15026 93832 15318
rect 94972 15038 95006 15330
rect 96030 15038 96064 15330
rect 97088 15038 97122 15330
rect 98146 15038 98180 15330
rect 99204 15038 99238 15330
rect 100262 15038 100296 15330
rect 62118 13580 62152 13872
rect 63176 13580 63210 13872
rect 64234 13580 64268 13872
rect 65292 13580 65326 13872
rect 66350 13580 66384 13872
rect 67408 13580 67442 13872
rect 68586 13578 68620 13870
rect 69644 13578 69678 13870
rect 70702 13578 70736 13870
rect 71760 13578 71794 13870
rect 72818 13578 72852 13870
rect 73876 13578 73910 13870
rect 75274 13552 75308 13844
rect 76332 13552 76366 13844
rect 77390 13552 77424 13844
rect 78448 13552 78482 13844
rect 79506 13552 79540 13844
rect 80564 13552 80598 13844
rect 81742 13550 81776 13842
rect 82800 13550 82834 13842
rect 83858 13550 83892 13842
rect 84916 13550 84950 13842
rect 85974 13550 86008 13842
rect 87032 13550 87066 13842
rect 88508 13544 88542 13836
rect 62118 12486 62152 12778
rect 63176 12486 63210 12778
rect 64234 12486 64268 12778
rect 65292 12486 65326 12778
rect 66350 12486 66384 12778
rect 89566 13544 89600 13836
rect 90624 13544 90658 13836
rect 91682 13544 91716 13836
rect 92740 13544 92774 13836
rect 93798 13544 93832 13836
rect 94976 13542 95010 13834
rect 67408 12486 67442 12778
rect 62118 11392 62152 11684
rect 63176 11392 63210 11684
rect 64234 11392 64268 11684
rect 65292 11392 65326 11684
rect 66350 11392 66384 11684
rect 67408 11392 67442 11684
rect 68586 12484 68620 12776
rect 69644 12484 69678 12776
rect 70702 12484 70736 12776
rect 71760 12484 71794 12776
rect 72818 12484 72852 12776
rect 96034 13542 96068 13834
rect 97092 13542 97126 13834
rect 98150 13542 98184 13834
rect 99208 13542 99242 13834
rect 100266 13542 100300 13834
rect 73876 12484 73910 12776
rect 62118 10298 62152 10590
rect 63176 10298 63210 10590
rect 64234 10298 64268 10590
rect 65292 10298 65326 10590
rect 66350 10298 66384 10590
rect 68586 11390 68620 11682
rect 69644 11390 69678 11682
rect 70702 11390 70736 11682
rect 71760 11390 71794 11682
rect 72818 11390 72852 11682
rect 73876 11390 73910 11682
rect 75274 12458 75308 12750
rect 76332 12458 76366 12750
rect 77390 12458 77424 12750
rect 78448 12458 78482 12750
rect 79506 12458 79540 12750
rect 80564 12458 80598 12750
rect 67408 10298 67442 10590
rect 68586 10296 68620 10588
rect 69644 10296 69678 10588
rect 70702 10296 70736 10588
rect 71760 10296 71794 10588
rect 72818 10296 72852 10588
rect 75274 11364 75308 11656
rect 76332 11364 76366 11656
rect 77390 11364 77424 11656
rect 78448 11364 78482 11656
rect 79506 11364 79540 11656
rect 80564 11364 80598 11656
rect 81742 12456 81776 12748
rect 82800 12456 82834 12748
rect 83858 12456 83892 12748
rect 84916 12456 84950 12748
rect 85974 12456 86008 12748
rect 87032 12456 87066 12748
rect 73876 10296 73910 10588
rect 75274 10270 75308 10562
rect 76332 10270 76366 10562
rect 77390 10270 77424 10562
rect 78448 10270 78482 10562
rect 79506 10270 79540 10562
rect 81742 11362 81776 11654
rect 82800 11362 82834 11654
rect 83858 11362 83892 11654
rect 84916 11362 84950 11654
rect 85974 11362 86008 11654
rect 87032 11362 87066 11654
rect 88508 12450 88542 12742
rect 89566 12450 89600 12742
rect 90624 12450 90658 12742
rect 91682 12450 91716 12742
rect 92740 12450 92774 12742
rect 93798 12450 93832 12742
rect 80564 10270 80598 10562
rect 81742 10268 81776 10560
rect 82800 10268 82834 10560
rect 83858 10268 83892 10560
rect 84916 10268 84950 10560
rect 85974 10268 86008 10560
rect 88508 11356 88542 11648
rect 89566 11356 89600 11648
rect 90624 11356 90658 11648
rect 91682 11356 91716 11648
rect 92740 11356 92774 11648
rect 93798 11356 93832 11648
rect 94976 12448 95010 12740
rect 96034 12448 96068 12740
rect 97092 12448 97126 12740
rect 98150 12448 98184 12740
rect 99208 12448 99242 12740
rect 100266 12448 100300 12740
rect 87032 10268 87066 10560
rect 88508 10262 88542 10554
rect 62118 9204 62152 9496
rect 63176 9204 63210 9496
rect 64234 9204 64268 9496
rect 65292 9204 65326 9496
rect 66350 9204 66384 9496
rect 89566 10262 89600 10554
rect 90624 10262 90658 10554
rect 91682 10262 91716 10554
rect 92740 10262 92774 10554
rect 94976 11354 95010 11646
rect 96034 11354 96068 11646
rect 97092 11354 97126 11646
rect 98150 11354 98184 11646
rect 99208 11354 99242 11646
rect 100266 11354 100300 11646
rect 93798 10262 93832 10554
rect 94976 10260 95010 10552
rect 67408 9204 67442 9496
rect 68586 9202 68620 9494
rect 69644 9202 69678 9494
rect 70702 9202 70736 9494
rect 71760 9202 71794 9494
rect 72818 9202 72852 9494
rect 96034 10260 96068 10552
rect 97092 10260 97126 10552
rect 98150 10260 98184 10552
rect 99208 10260 99242 10552
rect 100266 10260 100300 10552
rect 73876 9202 73910 9494
rect 75274 9176 75308 9468
rect 76332 9176 76366 9468
rect 77390 9176 77424 9468
rect 78448 9176 78482 9468
rect 79506 9176 79540 9468
rect 80564 9176 80598 9468
rect 81742 9174 81776 9466
rect 82800 9174 82834 9466
rect 83858 9174 83892 9466
rect 84916 9174 84950 9466
rect 85974 9174 86008 9466
rect 87032 9174 87066 9466
rect 88508 9168 88542 9460
rect 89566 9168 89600 9460
rect 90624 9168 90658 9460
rect 91682 9168 91716 9460
rect 92740 9168 92774 9460
rect 93798 9168 93832 9460
rect 94976 9166 95010 9458
rect 62118 7722 62152 8014
rect 63176 7722 63210 8014
rect 64234 7722 64268 8014
rect 65292 7722 65326 8014
rect 66350 7722 66384 8014
rect 96034 9166 96068 9458
rect 97092 9166 97126 9458
rect 98150 9166 98184 9458
rect 99208 9166 99242 9458
rect 100266 9166 100300 9458
rect 67408 7722 67442 8014
rect 68590 7720 68624 8012
rect 69648 7720 69682 8012
rect 70706 7720 70740 8012
rect 71764 7720 71798 8012
rect 72822 7720 72856 8012
rect 73880 7720 73914 8012
rect 75274 7694 75308 7986
rect 76332 7694 76366 7986
rect 77390 7694 77424 7986
rect 78448 7694 78482 7986
rect 79506 7694 79540 7986
rect 80564 7694 80598 7986
rect 81746 7692 81780 7984
rect 82804 7692 82838 7984
rect 83862 7692 83896 7984
rect 84920 7692 84954 7984
rect 85978 7692 86012 7984
rect 87036 7692 87070 7984
rect 88508 7686 88542 7978
rect 62118 6628 62152 6920
rect 63176 6628 63210 6920
rect 64234 6628 64268 6920
rect 65292 6628 65326 6920
rect 66350 6628 66384 6920
rect 89566 7686 89600 7978
rect 90624 7686 90658 7978
rect 91682 7686 91716 7978
rect 92740 7686 92774 7978
rect 93798 7686 93832 7978
rect 94980 7684 95014 7976
rect 67408 6628 67442 6920
rect 62118 5534 62152 5826
rect 63176 5534 63210 5826
rect 64234 5534 64268 5826
rect 65292 5534 65326 5826
rect 66350 5534 66384 5826
rect 67408 5534 67442 5826
rect 68590 6626 68624 6918
rect 69648 6626 69682 6918
rect 70706 6626 70740 6918
rect 71764 6626 71798 6918
rect 72822 6626 72856 6918
rect 96038 7684 96072 7976
rect 97096 7684 97130 7976
rect 98154 7684 98188 7976
rect 99212 7684 99246 7976
rect 100270 7684 100304 7976
rect 73880 6626 73914 6918
rect 62118 4440 62152 4732
rect 63176 4440 63210 4732
rect 64234 4440 64268 4732
rect 65292 4440 65326 4732
rect 66350 4440 66384 4732
rect 68590 5532 68624 5824
rect 69648 5532 69682 5824
rect 70706 5532 70740 5824
rect 71764 5532 71798 5824
rect 72822 5532 72856 5824
rect 73880 5532 73914 5824
rect 75274 6600 75308 6892
rect 76332 6600 76366 6892
rect 77390 6600 77424 6892
rect 78448 6600 78482 6892
rect 79506 6600 79540 6892
rect 80564 6600 80598 6892
rect 67408 4440 67442 4732
rect 68590 4438 68624 4730
rect 69648 4438 69682 4730
rect 70706 4438 70740 4730
rect 71764 4438 71798 4730
rect 72822 4438 72856 4730
rect 75274 5506 75308 5798
rect 76332 5506 76366 5798
rect 77390 5506 77424 5798
rect 78448 5506 78482 5798
rect 79506 5506 79540 5798
rect 80564 5506 80598 5798
rect 81746 6598 81780 6890
rect 82804 6598 82838 6890
rect 83862 6598 83896 6890
rect 84920 6598 84954 6890
rect 85978 6598 86012 6890
rect 87036 6598 87070 6890
rect 73880 4438 73914 4730
rect 75274 4412 75308 4704
rect 76332 4412 76366 4704
rect 77390 4412 77424 4704
rect 78448 4412 78482 4704
rect 79506 4412 79540 4704
rect 81746 5504 81780 5796
rect 82804 5504 82838 5796
rect 83862 5504 83896 5796
rect 84920 5504 84954 5796
rect 85978 5504 86012 5796
rect 87036 5504 87070 5796
rect 88508 6592 88542 6884
rect 89566 6592 89600 6884
rect 90624 6592 90658 6884
rect 91682 6592 91716 6884
rect 92740 6592 92774 6884
rect 93798 6592 93832 6884
rect 80564 4412 80598 4704
rect 81746 4410 81780 4702
rect 82804 4410 82838 4702
rect 83862 4410 83896 4702
rect 84920 4410 84954 4702
rect 85978 4410 86012 4702
rect 88508 5498 88542 5790
rect 89566 5498 89600 5790
rect 90624 5498 90658 5790
rect 91682 5498 91716 5790
rect 92740 5498 92774 5790
rect 93798 5498 93832 5790
rect 94980 6590 95014 6882
rect 96038 6590 96072 6882
rect 97096 6590 97130 6882
rect 98154 6590 98188 6882
rect 99212 6590 99246 6882
rect 100270 6590 100304 6882
rect 87036 4410 87070 4702
rect 88508 4404 88542 4696
rect 62118 3346 62152 3638
rect 63176 3346 63210 3638
rect 64234 3346 64268 3638
rect 65292 3346 65326 3638
rect 66350 3346 66384 3638
rect 89566 4404 89600 4696
rect 90624 4404 90658 4696
rect 91682 4404 91716 4696
rect 92740 4404 92774 4696
rect 94980 5496 95014 5788
rect 96038 5496 96072 5788
rect 97096 5496 97130 5788
rect 98154 5496 98188 5788
rect 99212 5496 99246 5788
rect 100270 5496 100304 5788
rect 93798 4404 93832 4696
rect 94980 4402 95014 4694
rect 67408 3346 67442 3638
rect 68590 3344 68624 3636
rect 69648 3344 69682 3636
rect 70706 3344 70740 3636
rect 71764 3344 71798 3636
rect 72822 3344 72856 3636
rect 96038 4402 96072 4694
rect 97096 4402 97130 4694
rect 98154 4402 98188 4694
rect 99212 4402 99246 4694
rect 100270 4402 100304 4694
rect 73880 3344 73914 3636
rect 75274 3318 75308 3610
rect 76332 3318 76366 3610
rect 77390 3318 77424 3610
rect 78448 3318 78482 3610
rect 79506 3318 79540 3610
rect 80564 3318 80598 3610
rect 81746 3316 81780 3608
rect 82804 3316 82838 3608
rect 83862 3316 83896 3608
rect 84920 3316 84954 3608
rect 85978 3316 86012 3608
rect 87036 3316 87070 3608
rect 88508 3310 88542 3602
rect 89566 3310 89600 3602
rect 90624 3310 90658 3602
rect 91682 3310 91716 3602
rect 92740 3310 92774 3602
rect 93798 3310 93832 3602
rect 94980 3308 95014 3600
rect 96038 3308 96072 3600
rect 97096 3308 97130 3600
rect 98154 3308 98188 3600
rect 99212 3308 99246 3600
rect 100270 3308 100304 3600
<< mvpdiffc >>
rect 42410 73194 42582 73228
rect 43104 73194 43276 73228
rect 43798 73194 43970 73228
rect 44492 73194 44664 73228
rect 45186 73194 45358 73228
rect 46418 73192 46590 73226
rect 47112 73192 47284 73226
rect 47806 73192 47978 73226
rect 48500 73192 48672 73226
rect 49194 73192 49366 73226
rect 50430 73192 50602 73226
rect 51124 73192 51296 73226
rect 51818 73192 51990 73226
rect 52512 73192 52684 73226
rect 53206 73192 53378 73226
rect 54440 73192 54612 73226
rect 55134 73192 55306 73226
rect 55828 73192 56000 73226
rect 56522 73192 56694 73226
rect 57216 73192 57388 73226
rect 42410 72536 42582 72570
rect 43104 72536 43276 72570
rect 43798 72536 43970 72570
rect 44492 72536 44664 72570
rect 45186 72536 45358 72570
rect 71338 73868 71372 74040
rect 71996 73868 72030 74040
rect 72654 73868 72688 74040
rect 73312 73868 73346 74040
rect 73970 73868 74004 74040
rect 75202 73848 75236 74020
rect 75860 73848 75894 74020
rect 76518 73848 76552 74020
rect 77176 73848 77210 74020
rect 77834 73848 77868 74020
rect 79052 73862 79086 74034
rect 79710 73862 79744 74034
rect 80368 73862 80402 74034
rect 81026 73862 81060 74034
rect 81684 73862 81718 74034
rect 46418 72534 46590 72568
rect 47112 72534 47284 72568
rect 47806 72534 47978 72568
rect 48500 72534 48672 72568
rect 49194 72534 49366 72568
rect 50430 72534 50602 72568
rect 51124 72534 51296 72568
rect 51818 72534 51990 72568
rect 52512 72534 52684 72568
rect 53206 72534 53378 72568
rect 54440 72534 54612 72568
rect 55134 72534 55306 72568
rect 55828 72534 56000 72568
rect 56522 72534 56694 72568
rect 57216 72534 57388 72568
rect 42410 71878 42582 71912
rect 43104 71878 43276 71912
rect 43798 71878 43970 71912
rect 44492 71878 44664 71912
rect 45186 71878 45358 71912
rect 46418 71876 46590 71910
rect 47112 71876 47284 71910
rect 47806 71876 47978 71910
rect 48500 71876 48672 71910
rect 49194 71876 49366 71910
rect 50430 71876 50602 71910
rect 51124 71876 51296 71910
rect 51818 71876 51990 71910
rect 52512 71876 52684 71910
rect 53206 71876 53378 71910
rect 54440 71876 54612 71910
rect 55134 71876 55306 71910
rect 55828 71876 56000 71910
rect 56522 71876 56694 71910
rect 57216 71876 57388 71910
rect 42410 71220 42582 71254
rect 43104 71220 43276 71254
rect 43798 71220 43970 71254
rect 44492 71220 44664 71254
rect 45186 71220 45358 71254
rect 46418 71218 46590 71252
rect 47112 71218 47284 71252
rect 47806 71218 47978 71252
rect 48500 71218 48672 71252
rect 49194 71218 49366 71252
rect 50430 71218 50602 71252
rect 51124 71218 51296 71252
rect 51818 71218 51990 71252
rect 52512 71218 52684 71252
rect 53206 71218 53378 71252
rect 54440 71218 54612 71252
rect 55134 71218 55306 71252
rect 55828 71218 56000 71252
rect 56522 71218 56694 71252
rect 57216 71218 57388 71252
rect 42410 70562 42582 70596
rect 43104 70562 43276 70596
rect 43798 70562 43970 70596
rect 44492 70562 44664 70596
rect 45186 70562 45358 70596
rect 46418 70560 46590 70594
rect 47112 70560 47284 70594
rect 47806 70560 47978 70594
rect 48500 70560 48672 70594
rect 49194 70560 49366 70594
rect 50430 70560 50602 70594
rect 51124 70560 51296 70594
rect 51818 70560 51990 70594
rect 52512 70560 52684 70594
rect 53206 70560 53378 70594
rect 54440 70560 54612 70594
rect 55134 70560 55306 70594
rect 55828 70560 56000 70594
rect 56522 70560 56694 70594
rect 57216 70560 57388 70594
rect 42410 69904 42582 69938
rect 43104 69904 43276 69938
rect 43798 69904 43970 69938
rect 44492 69904 44664 69938
rect 45186 69904 45358 69938
rect 46418 69902 46590 69936
rect 47112 69902 47284 69936
rect 47806 69902 47978 69936
rect 48500 69902 48672 69936
rect 49194 69902 49366 69936
rect 50430 69902 50602 69936
rect 51124 69902 51296 69936
rect 51818 69902 51990 69936
rect 52512 69902 52684 69936
rect 53206 69902 53378 69936
rect 54440 69902 54612 69936
rect 55134 69902 55306 69936
rect 55828 69902 56000 69936
rect 56522 69902 56694 69936
rect 57216 69902 57388 69936
rect 42402 68996 42574 69030
rect 43096 68996 43268 69030
rect 43790 68996 43962 69030
rect 44484 68996 44656 69030
rect 45178 68996 45350 69030
rect 46396 68996 46568 69030
rect 47090 68996 47262 69030
rect 47784 68996 47956 69030
rect 48478 68996 48650 69030
rect 49172 68996 49344 69030
rect 50418 68996 50590 69030
rect 51112 68996 51284 69030
rect 51806 68996 51978 69030
rect 52500 68996 52672 69030
rect 53194 68996 53366 69030
rect 54440 68996 54612 69030
rect 55134 68996 55306 69030
rect 55828 68996 56000 69030
rect 56522 68996 56694 69030
rect 57216 68996 57388 69030
rect 71310 72954 71344 73126
rect 71968 72954 72002 73126
rect 72626 72954 72660 73126
rect 73284 72954 73318 73126
rect 73942 72954 73976 73126
rect 71310 72260 71344 72432
rect 71968 72260 72002 72432
rect 72626 72260 72660 72432
rect 73284 72260 73318 72432
rect 73942 72260 73976 72432
rect 71310 71566 71344 71738
rect 71968 71566 72002 71738
rect 72626 71566 72660 71738
rect 73284 71566 73318 71738
rect 73942 71566 73976 71738
rect 71310 70872 71344 71044
rect 71968 70872 72002 71044
rect 72626 70872 72660 71044
rect 73284 70872 73318 71044
rect 73942 70872 73976 71044
rect 71310 70178 71344 70350
rect 71968 70178 72002 70350
rect 72626 70178 72660 70350
rect 73284 70178 73318 70350
rect 73942 70178 73976 70350
rect 75174 72934 75208 73106
rect 75832 72934 75866 73106
rect 76490 72934 76524 73106
rect 77148 72934 77182 73106
rect 77806 72934 77840 73106
rect 75174 72240 75208 72412
rect 75832 72240 75866 72412
rect 76490 72240 76524 72412
rect 77148 72240 77182 72412
rect 77806 72240 77840 72412
rect 75174 71546 75208 71718
rect 75832 71546 75866 71718
rect 76490 71546 76524 71718
rect 77148 71546 77182 71718
rect 77806 71546 77840 71718
rect 75174 70852 75208 71024
rect 75832 70852 75866 71024
rect 76490 70852 76524 71024
rect 77148 70852 77182 71024
rect 77806 70852 77840 71024
rect 75174 70158 75208 70330
rect 75832 70158 75866 70330
rect 76490 70158 76524 70330
rect 77148 70158 77182 70330
rect 77806 70158 77840 70330
rect 79024 72948 79058 73120
rect 79682 72948 79716 73120
rect 80340 72948 80374 73120
rect 80998 72948 81032 73120
rect 81656 72948 81690 73120
rect 79024 72254 79058 72426
rect 79682 72254 79716 72426
rect 80340 72254 80374 72426
rect 80998 72254 81032 72426
rect 81656 72254 81690 72426
rect 79024 71560 79058 71732
rect 79682 71560 79716 71732
rect 80340 71560 80374 71732
rect 80998 71560 81032 71732
rect 81656 71560 81690 71732
rect 79024 70866 79058 71038
rect 79682 70866 79716 71038
rect 80340 70866 80374 71038
rect 80998 70866 81032 71038
rect 81656 70866 81690 71038
rect 79024 70172 79058 70344
rect 79682 70172 79716 70344
rect 80340 70172 80374 70344
rect 80998 70172 81032 70344
rect 81656 70172 81690 70344
rect 42402 68338 42574 68372
rect 43096 68338 43268 68372
rect 43790 68338 43962 68372
rect 44484 68338 44656 68372
rect 45178 68338 45350 68372
rect 46396 68338 46568 68372
rect 47090 68338 47262 68372
rect 47784 68338 47956 68372
rect 48478 68338 48650 68372
rect 49172 68338 49344 68372
rect 50418 68338 50590 68372
rect 51112 68338 51284 68372
rect 51806 68338 51978 68372
rect 52500 68338 52672 68372
rect 53194 68338 53366 68372
rect 54440 68338 54612 68372
rect 55134 68338 55306 68372
rect 55828 68338 56000 68372
rect 56522 68338 56694 68372
rect 57216 68338 57388 68372
rect 42402 67680 42574 67714
rect 43096 67680 43268 67714
rect 43790 67680 43962 67714
rect 44484 67680 44656 67714
rect 45178 67680 45350 67714
rect 46396 67680 46568 67714
rect 47090 67680 47262 67714
rect 47784 67680 47956 67714
rect 48478 67680 48650 67714
rect 49172 67680 49344 67714
rect 50418 67680 50590 67714
rect 51112 67680 51284 67714
rect 51806 67680 51978 67714
rect 52500 67680 52672 67714
rect 53194 67680 53366 67714
rect 54440 67680 54612 67714
rect 55134 67680 55306 67714
rect 55828 67680 56000 67714
rect 56522 67680 56694 67714
rect 57216 67680 57388 67714
rect 42402 67022 42574 67056
rect 43096 67022 43268 67056
rect 43790 67022 43962 67056
rect 44484 67022 44656 67056
rect 45178 67022 45350 67056
rect 46396 67022 46568 67056
rect 47090 67022 47262 67056
rect 47784 67022 47956 67056
rect 48478 67022 48650 67056
rect 49172 67022 49344 67056
rect 50418 67022 50590 67056
rect 51112 67022 51284 67056
rect 51806 67022 51978 67056
rect 52500 67022 52672 67056
rect 53194 67022 53366 67056
rect 54440 67022 54612 67056
rect 55134 67022 55306 67056
rect 55828 67022 56000 67056
rect 56522 67022 56694 67056
rect 57216 67022 57388 67056
rect 42402 66364 42574 66398
rect 43096 66364 43268 66398
rect 43790 66364 43962 66398
rect 44484 66364 44656 66398
rect 45178 66364 45350 66398
rect 46396 66364 46568 66398
rect 47090 66364 47262 66398
rect 47784 66364 47956 66398
rect 48478 66364 48650 66398
rect 49172 66364 49344 66398
rect 50418 66364 50590 66398
rect 51112 66364 51284 66398
rect 51806 66364 51978 66398
rect 52500 66364 52672 66398
rect 53194 66364 53366 66398
rect 54440 66364 54612 66398
rect 55134 66364 55306 66398
rect 55828 66364 56000 66398
rect 56522 66364 56694 66398
rect 57216 66364 57388 66398
rect 71306 69178 71340 69350
rect 71964 69178 71998 69350
rect 72622 69178 72656 69350
rect 73280 69178 73314 69350
rect 73938 69178 73972 69350
rect 71306 68484 71340 68656
rect 71964 68484 71998 68656
rect 72622 68484 72656 68656
rect 73280 68484 73314 68656
rect 73938 68484 73972 68656
rect 71306 67790 71340 67962
rect 71964 67790 71998 67962
rect 72622 67790 72656 67962
rect 73280 67790 73314 67962
rect 73938 67790 73972 67962
rect 71306 67096 71340 67268
rect 71964 67096 71998 67268
rect 72622 67096 72656 67268
rect 73280 67096 73314 67268
rect 73938 67096 73972 67268
rect 966 65536 1138 65570
rect 1660 65536 1832 65570
rect 2354 65536 2526 65570
rect 3634 65532 3806 65566
rect 4328 65532 4500 65566
rect 5022 65532 5194 65566
rect 6308 65538 6480 65572
rect 7002 65538 7174 65572
rect 7696 65538 7868 65572
rect 8954 65538 9126 65572
rect 9648 65538 9820 65572
rect 10342 65538 10514 65572
rect 11608 65532 11780 65566
rect 966 64878 1138 64912
rect 1660 64878 1832 64912
rect 2354 64878 2526 64912
rect 12302 65532 12474 65566
rect 12996 65532 13168 65566
rect 14262 65538 14434 65572
rect 14956 65538 15128 65572
rect 15650 65538 15822 65572
rect 16888 65542 17060 65576
rect 17582 65542 17754 65576
rect 18276 65542 18448 65576
rect 19572 65586 19744 65620
rect 20266 65586 20438 65620
rect 3634 64874 3806 64908
rect 4328 64874 4500 64908
rect 5022 64874 5194 64908
rect 6308 64880 6480 64914
rect 7002 64880 7174 64914
rect 7696 64880 7868 64914
rect 8954 64880 9126 64914
rect 9648 64880 9820 64914
rect 10342 64880 10514 64914
rect 966 64220 1138 64254
rect 1660 64220 1832 64254
rect 2354 64220 2526 64254
rect 11608 64874 11780 64908
rect 12302 64874 12474 64908
rect 12996 64874 13168 64908
rect 14262 64880 14434 64914
rect 14956 64880 15128 64914
rect 15650 64880 15822 64914
rect 16888 64884 17060 64918
rect 17582 64884 17754 64918
rect 18276 64884 18448 64918
rect 19572 64928 19744 64962
rect 20266 64928 20438 64962
rect 3634 64216 3806 64250
rect 4328 64216 4500 64250
rect 5022 64216 5194 64250
rect 6308 64222 6480 64256
rect 7002 64222 7174 64256
rect 7696 64222 7868 64256
rect 8954 64222 9126 64256
rect 9648 64222 9820 64256
rect 10342 64222 10514 64256
rect 966 63562 1138 63596
rect 1660 63562 1832 63596
rect 2354 63562 2526 63596
rect 11608 64216 11780 64250
rect 12302 64216 12474 64250
rect 12996 64216 13168 64250
rect 14262 64222 14434 64256
rect 14956 64222 15128 64256
rect 15650 64222 15822 64256
rect 16888 64226 17060 64260
rect 17582 64226 17754 64260
rect 18276 64226 18448 64260
rect 19572 64270 19744 64304
rect 20266 64270 20438 64304
rect 3634 63558 3806 63592
rect 4328 63558 4500 63592
rect 5022 63558 5194 63592
rect 6308 63564 6480 63598
rect 7002 63564 7174 63598
rect 7696 63564 7868 63598
rect 8954 63564 9126 63598
rect 9648 63564 9820 63598
rect 10342 63564 10514 63598
rect 966 62904 1138 62938
rect 1660 62904 1832 62938
rect 2354 62904 2526 62938
rect 11608 63558 11780 63592
rect 12302 63558 12474 63592
rect 12996 63558 13168 63592
rect 14262 63564 14434 63598
rect 14956 63564 15128 63598
rect 15650 63564 15822 63598
rect 16888 63568 17060 63602
rect 17582 63568 17754 63602
rect 18276 63568 18448 63602
rect 19572 63612 19744 63646
rect 20266 63612 20438 63646
rect 3634 62900 3806 62934
rect 4328 62900 4500 62934
rect 5022 62900 5194 62934
rect 6308 62906 6480 62940
rect 7002 62906 7174 62940
rect 7696 62906 7868 62940
rect 8954 62906 9126 62940
rect 9648 62906 9820 62940
rect 10342 62906 10514 62940
rect 966 62246 1138 62280
rect 1660 62246 1832 62280
rect 2354 62246 2526 62280
rect 11608 62900 11780 62934
rect 12302 62900 12474 62934
rect 12996 62900 13168 62934
rect 14262 62906 14434 62940
rect 14956 62906 15128 62940
rect 15650 62906 15822 62940
rect 16888 62910 17060 62944
rect 17582 62910 17754 62944
rect 18276 62910 18448 62944
rect 19572 62954 19744 62988
rect 20266 62954 20438 62988
rect 3634 62242 3806 62276
rect 4328 62242 4500 62276
rect 5022 62242 5194 62276
rect 6308 62248 6480 62282
rect 7002 62248 7174 62282
rect 7696 62248 7868 62282
rect 8954 62248 9126 62282
rect 9648 62248 9820 62282
rect 10342 62248 10514 62282
rect 966 61588 1138 61622
rect 1660 61588 1832 61622
rect 2354 61588 2526 61622
rect 11608 62242 11780 62276
rect 12302 62242 12474 62276
rect 12996 62242 13168 62276
rect 14262 62248 14434 62282
rect 14956 62248 15128 62282
rect 15650 62248 15822 62282
rect 16888 62252 17060 62286
rect 17582 62252 17754 62286
rect 18276 62252 18448 62286
rect 19572 62296 19744 62330
rect 20266 62296 20438 62330
rect 3634 61584 3806 61618
rect 4328 61584 4500 61618
rect 5022 61584 5194 61618
rect 6308 61590 6480 61624
rect 7002 61590 7174 61624
rect 7696 61590 7868 61624
rect 8954 61590 9126 61624
rect 9648 61590 9820 61624
rect 10342 61590 10514 61624
rect 966 60930 1138 60964
rect 1660 60930 1832 60964
rect 2354 60930 2526 60964
rect 11608 61584 11780 61618
rect 12302 61584 12474 61618
rect 12996 61584 13168 61618
rect 14262 61590 14434 61624
rect 14956 61590 15128 61624
rect 15650 61590 15822 61624
rect 16888 61594 17060 61628
rect 17582 61594 17754 61628
rect 18276 61594 18448 61628
rect 19572 61638 19744 61672
rect 20266 61638 20438 61672
rect 3634 60926 3806 60960
rect 4328 60926 4500 60960
rect 5022 60926 5194 60960
rect 6308 60932 6480 60966
rect 7002 60932 7174 60966
rect 7696 60932 7868 60966
rect 8954 60932 9126 60966
rect 9648 60932 9820 60966
rect 10342 60932 10514 60966
rect 966 60272 1138 60306
rect 1660 60272 1832 60306
rect 11608 60926 11780 60960
rect 12302 60926 12474 60960
rect 12996 60926 13168 60960
rect 14262 60932 14434 60966
rect 14956 60932 15128 60966
rect 15650 60932 15822 60966
rect 16888 60936 17060 60970
rect 17582 60936 17754 60970
rect 18276 60936 18448 60970
rect 19572 60980 19744 61014
rect 20266 60980 20438 61014
rect 2354 60272 2526 60306
rect 3634 60268 3806 60302
rect 4328 60268 4500 60302
rect 5022 60268 5194 60302
rect 6308 60274 6480 60308
rect 7002 60274 7174 60308
rect 7696 60274 7868 60308
rect 8954 60274 9126 60308
rect 9648 60274 9820 60308
rect 10342 60274 10514 60308
rect 11608 60268 11780 60302
rect 12302 60268 12474 60302
rect 12996 60268 13168 60302
rect 14262 60274 14434 60308
rect 14956 60274 15128 60308
rect 15650 60274 15822 60308
rect 16888 60278 17060 60312
rect 17582 60278 17754 60312
rect 18276 60278 18448 60312
rect 19572 60322 19744 60356
rect 20266 60322 20438 60356
rect 938 59268 1110 59302
rect 1632 59268 1804 59302
rect 2326 59268 2498 59302
rect 3606 59264 3778 59298
rect 4300 59264 4472 59298
rect 4994 59264 5166 59298
rect 6280 59270 6452 59304
rect 6974 59270 7146 59304
rect 7668 59270 7840 59304
rect 8926 59270 9098 59304
rect 9620 59270 9792 59304
rect 10314 59270 10486 59304
rect 11580 59264 11752 59298
rect 938 58610 1110 58644
rect 1632 58610 1804 58644
rect 2326 58610 2498 58644
rect 12274 59264 12446 59298
rect 12968 59264 13140 59298
rect 14234 59270 14406 59304
rect 14928 59270 15100 59304
rect 15622 59270 15794 59304
rect 16860 59274 17032 59308
rect 17554 59274 17726 59308
rect 18248 59274 18420 59308
rect 19544 59318 19716 59352
rect 20238 59318 20410 59352
rect 3606 58606 3778 58640
rect 4300 58606 4472 58640
rect 4994 58606 5166 58640
rect 6280 58612 6452 58646
rect 6974 58612 7146 58646
rect 7668 58612 7840 58646
rect 8926 58612 9098 58646
rect 9620 58612 9792 58646
rect 10314 58612 10486 58646
rect 938 57952 1110 57986
rect 1632 57952 1804 57986
rect 2326 57952 2498 57986
rect 11580 58606 11752 58640
rect 12274 58606 12446 58640
rect 12968 58606 13140 58640
rect 14234 58612 14406 58646
rect 14928 58612 15100 58646
rect 15622 58612 15794 58646
rect 16860 58616 17032 58650
rect 17554 58616 17726 58650
rect 18248 58616 18420 58650
rect 19544 58660 19716 58694
rect 20238 58660 20410 58694
rect 3606 57948 3778 57982
rect 4300 57948 4472 57982
rect 4994 57948 5166 57982
rect 6280 57954 6452 57988
rect 6974 57954 7146 57988
rect 7668 57954 7840 57988
rect 8926 57954 9098 57988
rect 9620 57954 9792 57988
rect 10314 57954 10486 57988
rect 938 57294 1110 57328
rect 1632 57294 1804 57328
rect 2326 57294 2498 57328
rect 11580 57948 11752 57982
rect 12274 57948 12446 57982
rect 12968 57948 13140 57982
rect 14234 57954 14406 57988
rect 14928 57954 15100 57988
rect 15622 57954 15794 57988
rect 16860 57958 17032 57992
rect 17554 57958 17726 57992
rect 18248 57958 18420 57992
rect 19544 58002 19716 58036
rect 20238 58002 20410 58036
rect 3606 57290 3778 57324
rect 4300 57290 4472 57324
rect 4994 57290 5166 57324
rect 6280 57296 6452 57330
rect 6974 57296 7146 57330
rect 7668 57296 7840 57330
rect 8926 57296 9098 57330
rect 9620 57296 9792 57330
rect 10314 57296 10486 57330
rect 938 56636 1110 56670
rect 1632 56636 1804 56670
rect 2326 56636 2498 56670
rect 11580 57290 11752 57324
rect 12274 57290 12446 57324
rect 12968 57290 13140 57324
rect 14234 57296 14406 57330
rect 14928 57296 15100 57330
rect 15622 57296 15794 57330
rect 16860 57300 17032 57334
rect 17554 57300 17726 57334
rect 18248 57300 18420 57334
rect 19544 57344 19716 57378
rect 20238 57344 20410 57378
rect 3606 56632 3778 56666
rect 4300 56632 4472 56666
rect 4994 56632 5166 56666
rect 6280 56638 6452 56672
rect 6974 56638 7146 56672
rect 7668 56638 7840 56672
rect 8926 56638 9098 56672
rect 9620 56638 9792 56672
rect 10314 56638 10486 56672
rect 938 55978 1110 56012
rect 1632 55978 1804 56012
rect 2326 55978 2498 56012
rect 11580 56632 11752 56666
rect 12274 56632 12446 56666
rect 12968 56632 13140 56666
rect 14234 56638 14406 56672
rect 14928 56638 15100 56672
rect 15622 56638 15794 56672
rect 16860 56642 17032 56676
rect 17554 56642 17726 56676
rect 18248 56642 18420 56676
rect 19544 56686 19716 56720
rect 20238 56686 20410 56720
rect 3606 55974 3778 56008
rect 4300 55974 4472 56008
rect 4994 55974 5166 56008
rect 6280 55980 6452 56014
rect 6974 55980 7146 56014
rect 7668 55980 7840 56014
rect 8926 55980 9098 56014
rect 9620 55980 9792 56014
rect 10314 55980 10486 56014
rect 938 55320 1110 55354
rect 1632 55320 1804 55354
rect 2326 55320 2498 55354
rect 11580 55974 11752 56008
rect 12274 55974 12446 56008
rect 12968 55974 13140 56008
rect 14234 55980 14406 56014
rect 14928 55980 15100 56014
rect 15622 55980 15794 56014
rect 16860 55984 17032 56018
rect 17554 55984 17726 56018
rect 18248 55984 18420 56018
rect 19544 56028 19716 56062
rect 20238 56028 20410 56062
rect 3606 55316 3778 55350
rect 4300 55316 4472 55350
rect 4994 55316 5166 55350
rect 6280 55322 6452 55356
rect 6974 55322 7146 55356
rect 7668 55322 7840 55356
rect 8926 55322 9098 55356
rect 9620 55322 9792 55356
rect 10314 55322 10486 55356
rect 938 54662 1110 54696
rect 1632 54662 1804 54696
rect 2326 54662 2498 54696
rect 11580 55316 11752 55350
rect 12274 55316 12446 55350
rect 12968 55316 13140 55350
rect 14234 55322 14406 55356
rect 14928 55322 15100 55356
rect 15622 55322 15794 55356
rect 16860 55326 17032 55360
rect 17554 55326 17726 55360
rect 18248 55326 18420 55360
rect 19544 55370 19716 55404
rect 20238 55370 20410 55404
rect 3606 54658 3778 54692
rect 4300 54658 4472 54692
rect 4994 54658 5166 54692
rect 6280 54664 6452 54698
rect 6974 54664 7146 54698
rect 7668 54664 7840 54698
rect 8926 54664 9098 54698
rect 9620 54664 9792 54698
rect 10314 54664 10486 54698
rect 938 54004 1110 54038
rect 1632 54004 1804 54038
rect 11580 54658 11752 54692
rect 12274 54658 12446 54692
rect 12968 54658 13140 54692
rect 14234 54664 14406 54698
rect 14928 54664 15100 54698
rect 15622 54664 15794 54698
rect 16860 54668 17032 54702
rect 17554 54668 17726 54702
rect 18248 54668 18420 54702
rect 19544 54712 19716 54746
rect 20238 54712 20410 54746
rect 2326 54004 2498 54038
rect 3606 54000 3778 54034
rect 4300 54000 4472 54034
rect 4994 54000 5166 54034
rect 6280 54006 6452 54040
rect 6974 54006 7146 54040
rect 7668 54006 7840 54040
rect 8926 54006 9098 54040
rect 9620 54006 9792 54040
rect 10314 54006 10486 54040
rect 11580 54000 11752 54034
rect 12274 54000 12446 54034
rect 12968 54000 13140 54034
rect 14234 54006 14406 54040
rect 14928 54006 15100 54040
rect 15622 54006 15794 54040
rect 16860 54010 17032 54044
rect 17554 54010 17726 54044
rect 18248 54010 18420 54044
rect 19544 54054 19716 54088
rect 20238 54054 20410 54088
rect 938 52902 1110 52936
rect 1632 52902 1804 52936
rect 2326 52902 2498 52936
rect 3606 52898 3778 52932
rect 4300 52898 4472 52932
rect 4994 52898 5166 52932
rect 6280 52904 6452 52938
rect 6974 52904 7146 52938
rect 7668 52904 7840 52938
rect 8926 52904 9098 52938
rect 9620 52904 9792 52938
rect 10314 52904 10486 52938
rect 11580 52898 11752 52932
rect 938 52244 1110 52278
rect 1632 52244 1804 52278
rect 2326 52244 2498 52278
rect 12274 52898 12446 52932
rect 12968 52898 13140 52932
rect 14234 52904 14406 52938
rect 14928 52904 15100 52938
rect 15622 52904 15794 52938
rect 16860 52908 17032 52942
rect 17554 52908 17726 52942
rect 18248 52908 18420 52942
rect 19544 52952 19716 52986
rect 20238 52952 20410 52986
rect 3606 52240 3778 52274
rect 4300 52240 4472 52274
rect 4994 52240 5166 52274
rect 6280 52246 6452 52280
rect 6974 52246 7146 52280
rect 7668 52246 7840 52280
rect 8926 52246 9098 52280
rect 9620 52246 9792 52280
rect 10314 52246 10486 52280
rect 938 51586 1110 51620
rect 1632 51586 1804 51620
rect 2326 51586 2498 51620
rect 11580 52240 11752 52274
rect 12274 52240 12446 52274
rect 12968 52240 13140 52274
rect 14234 52246 14406 52280
rect 14928 52246 15100 52280
rect 15622 52246 15794 52280
rect 16860 52250 17032 52284
rect 17554 52250 17726 52284
rect 18248 52250 18420 52284
rect 19544 52294 19716 52328
rect 20238 52294 20410 52328
rect 3606 51582 3778 51616
rect 4300 51582 4472 51616
rect 4994 51582 5166 51616
rect 6280 51588 6452 51622
rect 6974 51588 7146 51622
rect 7668 51588 7840 51622
rect 8926 51588 9098 51622
rect 9620 51588 9792 51622
rect 10314 51588 10486 51622
rect 938 50928 1110 50962
rect 1632 50928 1804 50962
rect 2326 50928 2498 50962
rect 11580 51582 11752 51616
rect 12274 51582 12446 51616
rect 12968 51582 13140 51616
rect 14234 51588 14406 51622
rect 14928 51588 15100 51622
rect 15622 51588 15794 51622
rect 16860 51592 17032 51626
rect 17554 51592 17726 51626
rect 18248 51592 18420 51626
rect 19544 51636 19716 51670
rect 20238 51636 20410 51670
rect 3606 50924 3778 50958
rect 4300 50924 4472 50958
rect 4994 50924 5166 50958
rect 6280 50930 6452 50964
rect 6974 50930 7146 50964
rect 7668 50930 7840 50964
rect 8926 50930 9098 50964
rect 9620 50930 9792 50964
rect 10314 50930 10486 50964
rect 938 50270 1110 50304
rect 1632 50270 1804 50304
rect 2326 50270 2498 50304
rect 11580 50924 11752 50958
rect 12274 50924 12446 50958
rect 12968 50924 13140 50958
rect 14234 50930 14406 50964
rect 14928 50930 15100 50964
rect 15622 50930 15794 50964
rect 16860 50934 17032 50968
rect 17554 50934 17726 50968
rect 18248 50934 18420 50968
rect 19544 50978 19716 51012
rect 20238 50978 20410 51012
rect 3606 50266 3778 50300
rect 4300 50266 4472 50300
rect 4994 50266 5166 50300
rect 6280 50272 6452 50306
rect 6974 50272 7146 50306
rect 7668 50272 7840 50306
rect 8926 50272 9098 50306
rect 9620 50272 9792 50306
rect 10314 50272 10486 50306
rect 938 49612 1110 49646
rect 1632 49612 1804 49646
rect 2326 49612 2498 49646
rect 11580 50266 11752 50300
rect 12274 50266 12446 50300
rect 12968 50266 13140 50300
rect 14234 50272 14406 50306
rect 14928 50272 15100 50306
rect 15622 50272 15794 50306
rect 16860 50276 17032 50310
rect 17554 50276 17726 50310
rect 18248 50276 18420 50310
rect 19544 50320 19716 50354
rect 20238 50320 20410 50354
rect 3606 49608 3778 49642
rect 4300 49608 4472 49642
rect 4994 49608 5166 49642
rect 6280 49614 6452 49648
rect 6974 49614 7146 49648
rect 7668 49614 7840 49648
rect 8926 49614 9098 49648
rect 9620 49614 9792 49648
rect 10314 49614 10486 49648
rect 938 48954 1110 48988
rect 1632 48954 1804 48988
rect 2326 48954 2498 48988
rect 11580 49608 11752 49642
rect 12274 49608 12446 49642
rect 12968 49608 13140 49642
rect 14234 49614 14406 49648
rect 14928 49614 15100 49648
rect 15622 49614 15794 49648
rect 16860 49618 17032 49652
rect 17554 49618 17726 49652
rect 18248 49618 18420 49652
rect 19544 49662 19716 49696
rect 20238 49662 20410 49696
rect 3606 48950 3778 48984
rect 4300 48950 4472 48984
rect 4994 48950 5166 48984
rect 6280 48956 6452 48990
rect 6974 48956 7146 48990
rect 7668 48956 7840 48990
rect 8926 48956 9098 48990
rect 9620 48956 9792 48990
rect 10314 48956 10486 48990
rect 938 48296 1110 48330
rect 1632 48296 1804 48330
rect 2326 48296 2498 48330
rect 11580 48950 11752 48984
rect 12274 48950 12446 48984
rect 12968 48950 13140 48984
rect 14234 48956 14406 48990
rect 14928 48956 15100 48990
rect 15622 48956 15794 48990
rect 16860 48960 17032 48994
rect 17554 48960 17726 48994
rect 18248 48960 18420 48994
rect 19544 49004 19716 49038
rect 20238 49004 20410 49038
rect 3606 48292 3778 48326
rect 4300 48292 4472 48326
rect 4994 48292 5166 48326
rect 6280 48298 6452 48332
rect 6974 48298 7146 48332
rect 7668 48298 7840 48332
rect 8926 48298 9098 48332
rect 9620 48298 9792 48332
rect 10314 48298 10486 48332
rect 938 47638 1110 47672
rect 1632 47638 1804 47672
rect 11580 48292 11752 48326
rect 12274 48292 12446 48326
rect 12968 48292 13140 48326
rect 14234 48298 14406 48332
rect 14928 48298 15100 48332
rect 15622 48298 15794 48332
rect 16860 48302 17032 48336
rect 17554 48302 17726 48336
rect 18248 48302 18420 48336
rect 19544 48346 19716 48380
rect 20238 48346 20410 48380
rect 2326 47638 2498 47672
rect 3606 47634 3778 47668
rect 4300 47634 4472 47668
rect 4994 47634 5166 47668
rect 6280 47640 6452 47674
rect 6974 47640 7146 47674
rect 7668 47640 7840 47674
rect 8926 47640 9098 47674
rect 9620 47640 9792 47674
rect 10314 47640 10486 47674
rect 11580 47634 11752 47668
rect 12274 47634 12446 47668
rect 12968 47634 13140 47668
rect 14234 47640 14406 47674
rect 14928 47640 15100 47674
rect 15622 47640 15794 47674
rect 16860 47644 17032 47678
rect 17554 47644 17726 47678
rect 18248 47644 18420 47678
rect 19544 47688 19716 47722
rect 20238 47688 20410 47722
rect 42402 65706 42574 65740
rect 43096 65706 43268 65740
rect 43790 65706 43962 65740
rect 44484 65706 44656 65740
rect 45178 65706 45350 65740
rect 46396 65706 46568 65740
rect 47090 65706 47262 65740
rect 47784 65706 47956 65740
rect 48478 65706 48650 65740
rect 49172 65706 49344 65740
rect 50418 65706 50590 65740
rect 51112 65706 51284 65740
rect 51806 65706 51978 65740
rect 52500 65706 52672 65740
rect 53194 65706 53366 65740
rect 54440 65706 54612 65740
rect 55134 65706 55306 65740
rect 55828 65706 56000 65740
rect 56522 65706 56694 65740
rect 57216 65706 57388 65740
rect 71306 66402 71340 66574
rect 71964 66402 71998 66574
rect 72622 66402 72656 66574
rect 73280 66402 73314 66574
rect 73938 66402 73972 66574
rect 75170 69158 75204 69330
rect 75828 69158 75862 69330
rect 76486 69158 76520 69330
rect 77144 69158 77178 69330
rect 77802 69158 77836 69330
rect 75170 68464 75204 68636
rect 75828 68464 75862 68636
rect 76486 68464 76520 68636
rect 77144 68464 77178 68636
rect 77802 68464 77836 68636
rect 75170 67770 75204 67942
rect 75828 67770 75862 67942
rect 76486 67770 76520 67942
rect 77144 67770 77178 67942
rect 77802 67770 77836 67942
rect 75170 67076 75204 67248
rect 75828 67076 75862 67248
rect 76486 67076 76520 67248
rect 77144 67076 77178 67248
rect 77802 67076 77836 67248
rect 75170 66382 75204 66554
rect 75828 66382 75862 66554
rect 76486 66382 76520 66554
rect 77144 66382 77178 66554
rect 77802 66382 77836 66554
rect 79020 69172 79054 69344
rect 79678 69172 79712 69344
rect 80336 69172 80370 69344
rect 80994 69172 81028 69344
rect 81652 69172 81686 69344
rect 79020 68478 79054 68650
rect 79678 68478 79712 68650
rect 80336 68478 80370 68650
rect 80994 68478 81028 68650
rect 81652 68478 81686 68650
rect 79020 67784 79054 67956
rect 79678 67784 79712 67956
rect 80336 67784 80370 67956
rect 80994 67784 81028 67956
rect 81652 67784 81686 67956
rect 79020 67090 79054 67262
rect 79678 67090 79712 67262
rect 80336 67090 80370 67262
rect 80994 67090 81028 67262
rect 81652 67090 81686 67262
rect 79020 66396 79054 66568
rect 79678 66396 79712 66568
rect 80336 66396 80370 66568
rect 80994 66396 81028 66568
rect 81652 66396 81686 66568
rect 42390 64522 42562 64556
rect 43084 64522 43256 64556
rect 43778 64522 43950 64556
rect 44472 64522 44644 64556
rect 45166 64522 45338 64556
rect 46398 64520 46570 64554
rect 47092 64520 47264 64554
rect 47786 64520 47958 64554
rect 48480 64520 48652 64554
rect 49174 64520 49346 64554
rect 50410 64520 50582 64554
rect 51104 64520 51276 64554
rect 51798 64520 51970 64554
rect 52492 64520 52664 64554
rect 53186 64520 53358 64554
rect 54420 64520 54592 64554
rect 55114 64520 55286 64554
rect 55808 64520 55980 64554
rect 56502 64520 56674 64554
rect 57196 64520 57368 64554
rect 42390 63864 42562 63898
rect 43084 63864 43256 63898
rect 43778 63864 43950 63898
rect 44472 63864 44644 63898
rect 45166 63864 45338 63898
rect 46398 63862 46570 63896
rect 47092 63862 47264 63896
rect 47786 63862 47958 63896
rect 48480 63862 48652 63896
rect 49174 63862 49346 63896
rect 50410 63862 50582 63896
rect 51104 63862 51276 63896
rect 51798 63862 51970 63896
rect 52492 63862 52664 63896
rect 53186 63862 53358 63896
rect 54420 63862 54592 63896
rect 55114 63862 55286 63896
rect 55808 63862 55980 63896
rect 56502 63862 56674 63896
rect 57196 63862 57368 63896
rect 42390 63206 42562 63240
rect 43084 63206 43256 63240
rect 43778 63206 43950 63240
rect 44472 63206 44644 63240
rect 45166 63206 45338 63240
rect 46398 63204 46570 63238
rect 47092 63204 47264 63238
rect 47786 63204 47958 63238
rect 48480 63204 48652 63238
rect 49174 63204 49346 63238
rect 50410 63204 50582 63238
rect 51104 63204 51276 63238
rect 51798 63204 51970 63238
rect 52492 63204 52664 63238
rect 53186 63204 53358 63238
rect 54420 63204 54592 63238
rect 55114 63204 55286 63238
rect 55808 63204 55980 63238
rect 56502 63204 56674 63238
rect 57196 63204 57368 63238
rect 42390 62548 42562 62582
rect 43084 62548 43256 62582
rect 43778 62548 43950 62582
rect 44472 62548 44644 62582
rect 45166 62548 45338 62582
rect 46398 62546 46570 62580
rect 47092 62546 47264 62580
rect 47786 62546 47958 62580
rect 48480 62546 48652 62580
rect 49174 62546 49346 62580
rect 50410 62546 50582 62580
rect 51104 62546 51276 62580
rect 51798 62546 51970 62580
rect 52492 62546 52664 62580
rect 53186 62546 53358 62580
rect 54420 62546 54592 62580
rect 55114 62546 55286 62580
rect 55808 62546 55980 62580
rect 56502 62546 56674 62580
rect 57196 62546 57368 62580
rect 42390 61890 42562 61924
rect 43084 61890 43256 61924
rect 43778 61890 43950 61924
rect 44472 61890 44644 61924
rect 45166 61890 45338 61924
rect 71306 65408 71340 65580
rect 71964 65408 71998 65580
rect 72622 65408 72656 65580
rect 73280 65408 73314 65580
rect 73938 65408 73972 65580
rect 71306 64714 71340 64886
rect 71964 64714 71998 64886
rect 72622 64714 72656 64886
rect 73280 64714 73314 64886
rect 73938 64714 73972 64886
rect 71306 64020 71340 64192
rect 71964 64020 71998 64192
rect 72622 64020 72656 64192
rect 73280 64020 73314 64192
rect 73938 64020 73972 64192
rect 71306 63326 71340 63498
rect 71964 63326 71998 63498
rect 72622 63326 72656 63498
rect 73280 63326 73314 63498
rect 73938 63326 73972 63498
rect 46398 61888 46570 61922
rect 47092 61888 47264 61922
rect 47786 61888 47958 61922
rect 48480 61888 48652 61922
rect 49174 61888 49346 61922
rect 50410 61888 50582 61922
rect 51104 61888 51276 61922
rect 51798 61888 51970 61922
rect 52492 61888 52664 61922
rect 53186 61888 53358 61922
rect 54420 61888 54592 61922
rect 55114 61888 55286 61922
rect 55808 61888 55980 61922
rect 56502 61888 56674 61922
rect 57196 61888 57368 61922
rect 42390 61232 42562 61266
rect 43084 61232 43256 61266
rect 43778 61232 43950 61266
rect 44472 61232 44644 61266
rect 71306 62632 71340 62804
rect 71964 62632 71998 62804
rect 72622 62632 72656 62804
rect 73280 62632 73314 62804
rect 73938 62632 73972 62804
rect 75170 65388 75204 65560
rect 75828 65388 75862 65560
rect 76486 65388 76520 65560
rect 77144 65388 77178 65560
rect 77802 65388 77836 65560
rect 75170 64694 75204 64866
rect 75828 64694 75862 64866
rect 76486 64694 76520 64866
rect 77144 64694 77178 64866
rect 77802 64694 77836 64866
rect 75170 64000 75204 64172
rect 75828 64000 75862 64172
rect 76486 64000 76520 64172
rect 77144 64000 77178 64172
rect 77802 64000 77836 64172
rect 75170 63306 75204 63478
rect 75828 63306 75862 63478
rect 76486 63306 76520 63478
rect 77144 63306 77178 63478
rect 77802 63306 77836 63478
rect 75170 62612 75204 62784
rect 75828 62612 75862 62784
rect 76486 62612 76520 62784
rect 77144 62612 77178 62784
rect 77802 62612 77836 62784
rect 79020 65402 79054 65574
rect 79678 65402 79712 65574
rect 80336 65402 80370 65574
rect 80994 65402 81028 65574
rect 81652 65402 81686 65574
rect 79020 64708 79054 64880
rect 79678 64708 79712 64880
rect 80336 64708 80370 64880
rect 80994 64708 81028 64880
rect 81652 64708 81686 64880
rect 79020 64014 79054 64186
rect 79678 64014 79712 64186
rect 80336 64014 80370 64186
rect 80994 64014 81028 64186
rect 81652 64014 81686 64186
rect 79020 63320 79054 63492
rect 79678 63320 79712 63492
rect 80336 63320 80370 63492
rect 80994 63320 81028 63492
rect 81652 63320 81686 63492
rect 79020 62626 79054 62798
rect 79678 62626 79712 62798
rect 80336 62626 80370 62798
rect 80994 62626 81028 62798
rect 81652 62626 81686 62798
rect 45166 61232 45338 61266
rect 46398 61230 46570 61264
rect 47092 61230 47264 61264
rect 47786 61230 47958 61264
rect 48480 61230 48652 61264
rect 49174 61230 49346 61264
rect 50410 61230 50582 61264
rect 51104 61230 51276 61264
rect 51798 61230 51970 61264
rect 52492 61230 52664 61264
rect 53186 61230 53358 61264
rect 54420 61230 54592 61264
rect 55114 61230 55286 61264
rect 55808 61230 55980 61264
rect 56502 61230 56674 61264
rect 57196 61230 57368 61264
rect 42382 60324 42554 60358
rect 43076 60324 43248 60358
rect 43770 60324 43942 60358
rect 44464 60324 44636 60358
rect 45158 60324 45330 60358
rect 46376 60324 46548 60358
rect 47070 60324 47242 60358
rect 47764 60324 47936 60358
rect 48458 60324 48630 60358
rect 49152 60324 49324 60358
rect 50398 60324 50570 60358
rect 51092 60324 51264 60358
rect 51786 60324 51958 60358
rect 52480 60324 52652 60358
rect 53174 60324 53346 60358
rect 54420 60324 54592 60358
rect 55114 60324 55286 60358
rect 55808 60324 55980 60358
rect 56502 60324 56674 60358
rect 57196 60324 57368 60358
rect 42382 59666 42554 59700
rect 43076 59666 43248 59700
rect 43770 59666 43942 59700
rect 44464 59666 44636 59700
rect 45158 59666 45330 59700
rect 46376 59666 46548 59700
rect 47070 59666 47242 59700
rect 47764 59666 47936 59700
rect 48458 59666 48630 59700
rect 49152 59666 49324 59700
rect 50398 59666 50570 59700
rect 51092 59666 51264 59700
rect 51786 59666 51958 59700
rect 52480 59666 52652 59700
rect 53174 59666 53346 59700
rect 54420 59666 54592 59700
rect 55114 59666 55286 59700
rect 55808 59666 55980 59700
rect 56502 59666 56674 59700
rect 57196 59666 57368 59700
rect 42382 59008 42554 59042
rect 43076 59008 43248 59042
rect 43770 59008 43942 59042
rect 44464 59008 44636 59042
rect 45158 59008 45330 59042
rect 46376 59008 46548 59042
rect 47070 59008 47242 59042
rect 47764 59008 47936 59042
rect 48458 59008 48630 59042
rect 49152 59008 49324 59042
rect 50398 59008 50570 59042
rect 51092 59008 51264 59042
rect 51786 59008 51958 59042
rect 52480 59008 52652 59042
rect 53174 59008 53346 59042
rect 54420 59008 54592 59042
rect 55114 59008 55286 59042
rect 55808 59008 55980 59042
rect 56502 59008 56674 59042
rect 57196 59008 57368 59042
rect 42382 58350 42554 58384
rect 43076 58350 43248 58384
rect 43770 58350 43942 58384
rect 44464 58350 44636 58384
rect 45158 58350 45330 58384
rect 46376 58350 46548 58384
rect 47070 58350 47242 58384
rect 47764 58350 47936 58384
rect 48458 58350 48630 58384
rect 49152 58350 49324 58384
rect 50398 58350 50570 58384
rect 51092 58350 51264 58384
rect 51786 58350 51958 58384
rect 52480 58350 52652 58384
rect 53174 58350 53346 58384
rect 54420 58350 54592 58384
rect 55114 58350 55286 58384
rect 55808 58350 55980 58384
rect 56502 58350 56674 58384
rect 57196 58350 57368 58384
rect 42382 57692 42554 57726
rect 43076 57692 43248 57726
rect 43770 57692 43942 57726
rect 44464 57692 44636 57726
rect 45158 57692 45330 57726
rect 46376 57692 46548 57726
rect 47070 57692 47242 57726
rect 47764 57692 47936 57726
rect 48458 57692 48630 57726
rect 49152 57692 49324 57726
rect 50398 57692 50570 57726
rect 51092 57692 51264 57726
rect 51786 57692 51958 57726
rect 52480 57692 52652 57726
rect 53174 57692 53346 57726
rect 54420 57692 54592 57726
rect 55114 57692 55286 57726
rect 55808 57692 55980 57726
rect 56502 57692 56674 57726
rect 57196 57692 57368 57726
rect 71306 61644 71340 61816
rect 71964 61644 71998 61816
rect 72622 61644 72656 61816
rect 73280 61644 73314 61816
rect 73938 61644 73972 61816
rect 71306 60950 71340 61122
rect 71964 60950 71998 61122
rect 72622 60950 72656 61122
rect 73280 60950 73314 61122
rect 73938 60950 73972 61122
rect 71306 60256 71340 60428
rect 71964 60256 71998 60428
rect 72622 60256 72656 60428
rect 73280 60256 73314 60428
rect 73938 60256 73972 60428
rect 71306 59562 71340 59734
rect 71964 59562 71998 59734
rect 72622 59562 72656 59734
rect 73280 59562 73314 59734
rect 73938 59562 73972 59734
rect 71306 58868 71340 59040
rect 71964 58868 71998 59040
rect 72622 58868 72656 59040
rect 73280 58868 73314 59040
rect 73938 58868 73972 59040
rect 75170 61624 75204 61796
rect 75828 61624 75862 61796
rect 76486 61624 76520 61796
rect 77144 61624 77178 61796
rect 77802 61624 77836 61796
rect 75170 60930 75204 61102
rect 75828 60930 75862 61102
rect 76486 60930 76520 61102
rect 77144 60930 77178 61102
rect 77802 60930 77836 61102
rect 75170 60236 75204 60408
rect 75828 60236 75862 60408
rect 76486 60236 76520 60408
rect 77144 60236 77178 60408
rect 77802 60236 77836 60408
rect 75170 59542 75204 59714
rect 75828 59542 75862 59714
rect 76486 59542 76520 59714
rect 77144 59542 77178 59714
rect 77802 59542 77836 59714
rect 75170 58848 75204 59020
rect 75828 58848 75862 59020
rect 76486 58848 76520 59020
rect 77144 58848 77178 59020
rect 77802 58848 77836 59020
rect 79020 61638 79054 61810
rect 79678 61638 79712 61810
rect 80336 61638 80370 61810
rect 80994 61638 81028 61810
rect 81652 61638 81686 61810
rect 79020 60944 79054 61116
rect 79678 60944 79712 61116
rect 80336 60944 80370 61116
rect 80994 60944 81028 61116
rect 81652 60944 81686 61116
rect 79020 60250 79054 60422
rect 79678 60250 79712 60422
rect 80336 60250 80370 60422
rect 80994 60250 81028 60422
rect 81652 60250 81686 60422
rect 79020 59556 79054 59728
rect 79678 59556 79712 59728
rect 80336 59556 80370 59728
rect 80994 59556 81028 59728
rect 81652 59556 81686 59728
rect 79020 58862 79054 59034
rect 79678 58862 79712 59034
rect 80336 58862 80370 59034
rect 80994 58862 81028 59034
rect 81652 58862 81686 59034
rect 42382 57034 42554 57068
rect 43076 57034 43248 57068
rect 43770 57034 43942 57068
rect 44464 57034 44636 57068
rect 45158 57034 45330 57068
rect 46376 57034 46548 57068
rect 47070 57034 47242 57068
rect 47764 57034 47936 57068
rect 48458 57034 48630 57068
rect 49152 57034 49324 57068
rect 50398 57034 50570 57068
rect 51092 57034 51264 57068
rect 51786 57034 51958 57068
rect 52480 57034 52652 57068
rect 53174 57034 53346 57068
rect 54420 57034 54592 57068
rect 55114 57034 55286 57068
rect 55808 57034 55980 57068
rect 56502 57034 56674 57068
rect 57196 57034 57368 57068
rect 42334 55934 42506 55968
rect 43028 55934 43200 55968
rect 43722 55934 43894 55968
rect 44416 55934 44588 55968
rect 45110 55934 45282 55968
rect 46342 55932 46514 55966
rect 47036 55932 47208 55966
rect 47730 55932 47902 55966
rect 48424 55932 48596 55966
rect 49118 55932 49290 55966
rect 50354 55932 50526 55966
rect 51048 55932 51220 55966
rect 51742 55932 51914 55966
rect 52436 55932 52608 55966
rect 53130 55932 53302 55966
rect 54364 55932 54536 55966
rect 55058 55932 55230 55966
rect 55752 55932 55924 55966
rect 56446 55932 56618 55966
rect 57140 55932 57312 55966
rect 42334 55276 42506 55310
rect 43028 55276 43200 55310
rect 43722 55276 43894 55310
rect 44416 55276 44588 55310
rect 45110 55276 45282 55310
rect 46342 55274 46514 55308
rect 47036 55274 47208 55308
rect 47730 55274 47902 55308
rect 48424 55274 48596 55308
rect 49118 55274 49290 55308
rect 50354 55274 50526 55308
rect 51048 55274 51220 55308
rect 51742 55274 51914 55308
rect 52436 55274 52608 55308
rect 53130 55274 53302 55308
rect 54364 55274 54536 55308
rect 55058 55274 55230 55308
rect 55752 55274 55924 55308
rect 56446 55274 56618 55308
rect 57140 55274 57312 55308
rect 42334 54618 42506 54652
rect 43028 54618 43200 54652
rect 43722 54618 43894 54652
rect 44416 54618 44588 54652
rect 45110 54618 45282 54652
rect 46342 54616 46514 54650
rect 47036 54616 47208 54650
rect 47730 54616 47902 54650
rect 48424 54616 48596 54650
rect 49118 54616 49290 54650
rect 50354 54616 50526 54650
rect 51048 54616 51220 54650
rect 51742 54616 51914 54650
rect 52436 54616 52608 54650
rect 53130 54616 53302 54650
rect 54364 54616 54536 54650
rect 55058 54616 55230 54650
rect 55752 54616 55924 54650
rect 56446 54616 56618 54650
rect 57140 54616 57312 54650
rect 42334 53960 42506 53994
rect 43028 53960 43200 53994
rect 43722 53960 43894 53994
rect 44416 53960 44588 53994
rect 45110 53960 45282 53994
rect 46342 53958 46514 53992
rect 47036 53958 47208 53992
rect 47730 53958 47902 53992
rect 48424 53958 48596 53992
rect 49118 53958 49290 53992
rect 50354 53958 50526 53992
rect 51048 53958 51220 53992
rect 51742 53958 51914 53992
rect 52436 53958 52608 53992
rect 53130 53958 53302 53992
rect 54364 53958 54536 53992
rect 55058 53958 55230 53992
rect 55752 53958 55924 53992
rect 56446 53958 56618 53992
rect 57140 53958 57312 53992
rect 42334 53302 42506 53336
rect 43028 53302 43200 53336
rect 43722 53302 43894 53336
rect 44416 53302 44588 53336
rect 45110 53302 45282 53336
rect 71306 57868 71340 58040
rect 71964 57868 71998 58040
rect 72622 57868 72656 58040
rect 73280 57868 73314 58040
rect 73938 57868 73972 58040
rect 71306 57174 71340 57346
rect 71964 57174 71998 57346
rect 72622 57174 72656 57346
rect 73280 57174 73314 57346
rect 73938 57174 73972 57346
rect 71306 56480 71340 56652
rect 71964 56480 71998 56652
rect 72622 56480 72656 56652
rect 73280 56480 73314 56652
rect 73938 56480 73972 56652
rect 71306 55786 71340 55958
rect 71964 55786 71998 55958
rect 72622 55786 72656 55958
rect 73280 55786 73314 55958
rect 73938 55786 73972 55958
rect 71306 55092 71340 55264
rect 71964 55092 71998 55264
rect 72622 55092 72656 55264
rect 73280 55092 73314 55264
rect 73938 55092 73972 55264
rect 75170 57848 75204 58020
rect 75828 57848 75862 58020
rect 76486 57848 76520 58020
rect 77144 57848 77178 58020
rect 77802 57848 77836 58020
rect 75170 57154 75204 57326
rect 75828 57154 75862 57326
rect 76486 57154 76520 57326
rect 77144 57154 77178 57326
rect 77802 57154 77836 57326
rect 75170 56460 75204 56632
rect 75828 56460 75862 56632
rect 76486 56460 76520 56632
rect 77144 56460 77178 56632
rect 77802 56460 77836 56632
rect 75170 55766 75204 55938
rect 75828 55766 75862 55938
rect 76486 55766 76520 55938
rect 77144 55766 77178 55938
rect 77802 55766 77836 55938
rect 75170 55072 75204 55244
rect 75828 55072 75862 55244
rect 76486 55072 76520 55244
rect 77144 55072 77178 55244
rect 77802 55072 77836 55244
rect 79020 57862 79054 58034
rect 79678 57862 79712 58034
rect 80336 57862 80370 58034
rect 80994 57862 81028 58034
rect 81652 57862 81686 58034
rect 79020 57168 79054 57340
rect 79678 57168 79712 57340
rect 80336 57168 80370 57340
rect 80994 57168 81028 57340
rect 81652 57168 81686 57340
rect 79020 56474 79054 56646
rect 79678 56474 79712 56646
rect 80336 56474 80370 56646
rect 80994 56474 81028 56646
rect 81652 56474 81686 56646
rect 79020 55780 79054 55952
rect 79678 55780 79712 55952
rect 80336 55780 80370 55952
rect 80994 55780 81028 55952
rect 81652 55780 81686 55952
rect 79020 55086 79054 55258
rect 79678 55086 79712 55258
rect 80336 55086 80370 55258
rect 80994 55086 81028 55258
rect 81652 55086 81686 55258
rect 46342 53300 46514 53334
rect 47036 53300 47208 53334
rect 47730 53300 47902 53334
rect 48424 53300 48596 53334
rect 49118 53300 49290 53334
rect 50354 53300 50526 53334
rect 51048 53300 51220 53334
rect 51742 53300 51914 53334
rect 52436 53300 52608 53334
rect 53130 53300 53302 53334
rect 54364 53300 54536 53334
rect 55058 53300 55230 53334
rect 55752 53300 55924 53334
rect 56446 53300 56618 53334
rect 57140 53300 57312 53334
rect 42334 52644 42506 52678
rect 43028 52644 43200 52678
rect 43722 52644 43894 52678
rect 44416 52644 44588 52678
rect 45110 52644 45282 52678
rect 46342 52642 46514 52676
rect 47036 52642 47208 52676
rect 47730 52642 47902 52676
rect 48424 52642 48596 52676
rect 49118 52642 49290 52676
rect 50354 52642 50526 52676
rect 51048 52642 51220 52676
rect 51742 52642 51914 52676
rect 52436 52642 52608 52676
rect 53130 52642 53302 52676
rect 54364 52642 54536 52676
rect 55058 52642 55230 52676
rect 55752 52642 55924 52676
rect 56446 52642 56618 52676
rect 57140 52642 57312 52676
rect 42326 51736 42498 51770
rect 43020 51736 43192 51770
rect 43714 51736 43886 51770
rect 44408 51736 44580 51770
rect 45102 51736 45274 51770
rect 46320 51736 46492 51770
rect 47014 51736 47186 51770
rect 47708 51736 47880 51770
rect 48402 51736 48574 51770
rect 49096 51736 49268 51770
rect 50342 51736 50514 51770
rect 51036 51736 51208 51770
rect 51730 51736 51902 51770
rect 52424 51736 52596 51770
rect 53118 51736 53290 51770
rect 54364 51736 54536 51770
rect 55058 51736 55230 51770
rect 55752 51736 55924 51770
rect 56446 51736 56618 51770
rect 57140 51736 57312 51770
rect 71310 54096 71344 54268
rect 71968 54096 72002 54268
rect 72626 54096 72660 54268
rect 73284 54096 73318 54268
rect 73942 54096 73976 54268
rect 71310 53402 71344 53574
rect 71968 53402 72002 53574
rect 72626 53402 72660 53574
rect 73284 53402 73318 53574
rect 73942 53402 73976 53574
rect 71310 52708 71344 52880
rect 71968 52708 72002 52880
rect 72626 52708 72660 52880
rect 73284 52708 73318 52880
rect 73942 52708 73976 52880
rect 71310 52014 71344 52186
rect 71968 52014 72002 52186
rect 72626 52014 72660 52186
rect 73284 52014 73318 52186
rect 73942 52014 73976 52186
rect 42326 51078 42498 51112
rect 43020 51078 43192 51112
rect 43714 51078 43886 51112
rect 44408 51078 44580 51112
rect 45102 51078 45274 51112
rect 46320 51078 46492 51112
rect 47014 51078 47186 51112
rect 47708 51078 47880 51112
rect 48402 51078 48574 51112
rect 49096 51078 49268 51112
rect 50342 51078 50514 51112
rect 51036 51078 51208 51112
rect 51730 51078 51902 51112
rect 52424 51078 52596 51112
rect 53118 51078 53290 51112
rect 54364 51078 54536 51112
rect 55058 51078 55230 51112
rect 55752 51078 55924 51112
rect 56446 51078 56618 51112
rect 57140 51078 57312 51112
rect 71310 51320 71344 51492
rect 71968 51320 72002 51492
rect 72626 51320 72660 51492
rect 73284 51320 73318 51492
rect 73942 51320 73976 51492
rect 75174 54076 75208 54248
rect 75832 54076 75866 54248
rect 76490 54076 76524 54248
rect 77148 54076 77182 54248
rect 77806 54076 77840 54248
rect 75174 53382 75208 53554
rect 75832 53382 75866 53554
rect 76490 53382 76524 53554
rect 77148 53382 77182 53554
rect 77806 53382 77840 53554
rect 75174 52688 75208 52860
rect 75832 52688 75866 52860
rect 76490 52688 76524 52860
rect 77148 52688 77182 52860
rect 77806 52688 77840 52860
rect 75174 51994 75208 52166
rect 75832 51994 75866 52166
rect 76490 51994 76524 52166
rect 77148 51994 77182 52166
rect 77806 51994 77840 52166
rect 75174 51300 75208 51472
rect 75832 51300 75866 51472
rect 76490 51300 76524 51472
rect 77148 51300 77182 51472
rect 77806 51300 77840 51472
rect 79024 54090 79058 54262
rect 79682 54090 79716 54262
rect 80340 54090 80374 54262
rect 80998 54090 81032 54262
rect 81656 54090 81690 54262
rect 79024 53396 79058 53568
rect 79682 53396 79716 53568
rect 80340 53396 80374 53568
rect 80998 53396 81032 53568
rect 81656 53396 81690 53568
rect 79024 52702 79058 52874
rect 79682 52702 79716 52874
rect 80340 52702 80374 52874
rect 80998 52702 81032 52874
rect 81656 52702 81690 52874
rect 79024 52008 79058 52180
rect 79682 52008 79716 52180
rect 80340 52008 80374 52180
rect 80998 52008 81032 52180
rect 81656 52008 81690 52180
rect 79024 51314 79058 51486
rect 79682 51314 79716 51486
rect 80340 51314 80374 51486
rect 80998 51314 81032 51486
rect 81656 51314 81690 51486
rect 83310 53909 83344 53943
rect 83310 53817 83344 53851
rect 83466 53913 83500 53947
rect 83466 53813 83500 53847
rect 83622 53909 83656 53943
rect 83736 53908 83770 53942
rect 83892 53942 83926 53976
rect 84048 53908 84082 53942
rect 84204 53916 84238 53950
rect 84502 53927 84536 53961
rect 84674 53916 84708 53950
rect 84846 53964 84880 53998
rect 83622 53817 83656 53851
rect 85002 53819 85036 53853
rect 85158 53969 85192 54003
rect 85158 53894 85192 53928
rect 86116 53965 86150 53999
rect 85158 53819 85192 53853
rect 85479 53836 85513 53870
rect 85656 53836 85690 53870
rect 85812 53849 85846 53883
rect 86116 53885 86150 53919
rect 85941 53819 85975 53853
rect 85941 53719 85975 53753
rect 86116 53803 86150 53837
rect 86116 53723 86150 53757
rect 86272 53965 86306 53999
rect 86272 53885 86306 53919
rect 86272 53803 86306 53837
rect 86272 53723 86306 53757
rect 42326 50420 42498 50454
rect 43020 50420 43192 50454
rect 43714 50420 43886 50454
rect 44408 50420 44580 50454
rect 45102 50420 45274 50454
rect 46320 50420 46492 50454
rect 47014 50420 47186 50454
rect 47708 50420 47880 50454
rect 48402 50420 48574 50454
rect 49096 50420 49268 50454
rect 50342 50420 50514 50454
rect 51036 50420 51208 50454
rect 51730 50420 51902 50454
rect 52424 50420 52596 50454
rect 53118 50420 53290 50454
rect 54364 50420 54536 50454
rect 55058 50420 55230 50454
rect 55752 50420 55924 50454
rect 56446 50420 56618 50454
rect 57140 50420 57312 50454
rect 42326 49762 42498 49796
rect 43020 49762 43192 49796
rect 43714 49762 43886 49796
rect 44408 49762 44580 49796
rect 45102 49762 45274 49796
rect 46320 49762 46492 49796
rect 47014 49762 47186 49796
rect 47708 49762 47880 49796
rect 48402 49762 48574 49796
rect 49096 49762 49268 49796
rect 50342 49762 50514 49796
rect 51036 49762 51208 49796
rect 51730 49762 51902 49796
rect 52424 49762 52596 49796
rect 53118 49762 53290 49796
rect 54364 49762 54536 49796
rect 55058 49762 55230 49796
rect 55752 49762 55924 49796
rect 56446 49762 56618 49796
rect 57140 49762 57312 49796
rect 42326 49104 42498 49138
rect 43020 49104 43192 49138
rect 43714 49104 43886 49138
rect 44408 49104 44580 49138
rect 45102 49104 45274 49138
rect 46320 49104 46492 49138
rect 47014 49104 47186 49138
rect 47708 49104 47880 49138
rect 48402 49104 48574 49138
rect 49096 49104 49268 49138
rect 50342 49104 50514 49138
rect 51036 49104 51208 49138
rect 51730 49104 51902 49138
rect 52424 49104 52596 49138
rect 53118 49104 53290 49138
rect 54364 49104 54536 49138
rect 55058 49104 55230 49138
rect 55752 49104 55924 49138
rect 56446 49104 56618 49138
rect 57140 49104 57312 49138
rect 42326 48446 42498 48480
rect 43020 48446 43192 48480
rect 43714 48446 43886 48480
rect 44408 48446 44580 48480
rect 45102 48446 45274 48480
rect 46320 48446 46492 48480
rect 47014 48446 47186 48480
rect 47708 48446 47880 48480
rect 48402 48446 48574 48480
rect 49096 48446 49268 48480
rect 50342 48446 50514 48480
rect 51036 48446 51208 48480
rect 51730 48446 51902 48480
rect 52424 48446 52596 48480
rect 53118 48446 53290 48480
rect 54364 48446 54536 48480
rect 55058 48446 55230 48480
rect 55752 48446 55924 48480
rect 56446 48446 56618 48480
rect 57140 48446 57312 48480
<< mvpsubdiff >>
rect 30576 58170 30928 58184
rect 22890 57656 30928 58170
rect 22890 55346 23242 57656
rect 28686 55970 29576 55990
rect 24274 55868 25162 55908
rect 24274 55766 24368 55868
rect 25098 55766 25162 55868
rect 28686 55872 28714 55970
rect 29532 55872 29576 55970
rect 28686 55848 29576 55872
rect 24274 55732 25162 55766
rect 22890 54924 22980 55346
rect 23102 54924 23242 55346
rect 22890 52204 23242 54924
rect 28692 54080 29582 54100
rect 24280 53978 25168 54018
rect 24280 53876 24374 53978
rect 25104 53876 25168 53978
rect 28692 53982 28720 54080
rect 29538 53982 29582 54080
rect 28692 53958 29582 53982
rect 24280 53842 25168 53876
rect 30576 52204 30928 57656
rect 22890 52138 30928 52204
rect 22890 52040 28736 52138
rect 29554 52040 30928 52138
rect 22890 52036 30928 52040
rect 22890 51934 24390 52036
rect 25120 51934 30928 52036
rect 22890 51718 30928 51934
rect 22890 51704 30900 51718
rect 23066 51690 30900 51704
rect 83272 53251 83303 53285
rect 83337 53251 83399 53285
rect 83433 53251 83495 53285
rect 83529 53251 83591 53285
rect 83625 53251 83687 53285
rect 83721 53251 83783 53285
rect 83817 53251 83879 53285
rect 83913 53251 83975 53285
rect 84009 53251 84071 53285
rect 84105 53251 84167 53285
rect 84201 53251 84263 53285
rect 84297 53251 84359 53285
rect 84393 53251 84455 53285
rect 84489 53251 84551 53285
rect 84585 53251 84647 53285
rect 84681 53251 84743 53285
rect 84777 53251 84839 53285
rect 84873 53251 84935 53285
rect 84969 53251 85031 53285
rect 85065 53251 85127 53285
rect 85161 53251 85223 53285
rect 85257 53251 85319 53285
rect 85353 53251 85415 53285
rect 85449 53251 85511 53285
rect 85545 53251 85607 53285
rect 85641 53251 85703 53285
rect 85737 53251 85799 53285
rect 85833 53251 85895 53285
rect 85929 53251 85991 53285
rect 86025 53251 86087 53285
rect 86121 53251 86183 53285
rect 86217 53251 86279 53285
rect 86313 53251 86344 53285
rect 0 45406 60208 45432
rect 0 45148 60238 45406
rect 0 44998 38946 45148
rect 0 44696 24240 44998
rect 25328 44696 38946 44998
rect 0 44424 38946 44696
rect 42360 44424 60238 45148
rect 0 44094 60238 44424
rect 48 41518 1702 44094
rect 48 40322 1326 41518
rect 1420 40322 1702 41518
rect 7794 41526 8002 41688
rect 48 35702 1702 40322
rect 7794 40330 7840 41526
rect 7934 40330 8002 41526
rect 14300 41534 14508 41696
rect 7794 39966 8002 40330
rect 14300 40338 14346 41534
rect 14440 40338 14508 41534
rect 20790 41518 20998 41680
rect 14300 39974 14508 40338
rect 20790 40322 20836 41518
rect 20930 40322 20998 41518
rect 27312 41534 27520 41696
rect 20790 39958 20998 40322
rect 27312 40338 27358 41534
rect 27452 40338 27520 41534
rect 33822 41540 34030 41702
rect 27312 39974 27520 40338
rect 33822 40344 33868 41540
rect 33962 40344 34030 41540
rect 40312 41540 40520 41702
rect 33822 39980 34030 40344
rect 40312 40344 40358 41540
rect 40452 40344 40520 41540
rect 46900 41562 47108 41724
rect 40312 39980 40520 40344
rect 46900 40366 46946 41562
rect 47040 40366 47108 41562
rect 53414 41576 53622 41738
rect 46900 40002 47108 40366
rect 53414 40380 53460 41576
rect 53554 40380 53622 41576
rect 59558 41952 60238 44094
rect 62020 43950 73948 44040
rect 62020 43808 68330 43950
rect 68980 43808 73948 43950
rect 62020 43744 73948 43808
rect 59530 41772 60238 41952
rect 53414 40016 53622 40380
rect 59530 40204 59572 41772
rect 59836 40204 60238 41772
rect 59530 40066 60238 40204
rect 48 34506 1326 35702
rect 1420 34506 1702 35702
rect 7794 35710 8002 35872
rect 48 29868 1702 34506
rect 7794 34514 7840 35710
rect 7934 34514 8002 35710
rect 14300 35718 14508 35880
rect 7794 34150 8002 34514
rect 14300 34522 14346 35718
rect 14440 34522 14508 35718
rect 20790 35702 20998 35864
rect 14300 34158 14508 34522
rect 20790 34506 20836 35702
rect 20930 34506 20998 35702
rect 27312 35718 27520 35880
rect 20790 34142 20998 34506
rect 27312 34522 27358 35718
rect 27452 34522 27520 35718
rect 33822 35724 34030 35886
rect 27312 34158 27520 34522
rect 33822 34528 33868 35724
rect 33962 34528 34030 35724
rect 40312 35724 40520 35886
rect 33822 34164 34030 34528
rect 40312 34528 40358 35724
rect 40452 34528 40520 35724
rect 46900 35746 47108 35908
rect 40312 34164 40520 34528
rect 46900 34550 46946 35746
rect 47040 34550 47108 35746
rect 53414 35760 53622 35922
rect 46900 34186 47108 34550
rect 53414 34564 53460 35760
rect 53554 34564 53622 35760
rect 59558 35834 60238 40066
rect 62072 42630 62406 43744
rect 73592 43002 73946 43744
rect 73592 42876 73950 43002
rect 62072 40876 62180 42630
rect 62328 40876 62406 42630
rect 65942 42632 66154 42702
rect 62072 39664 62406 40876
rect 65942 40878 65974 42632
rect 66122 40878 66154 42632
rect 69750 42646 69962 42716
rect 65942 40792 66154 40878
rect 69750 40892 69782 42646
rect 69930 40892 69962 42646
rect 69750 40806 69962 40892
rect 73592 40970 73646 42876
rect 73876 40970 73950 42876
rect 73592 40668 73950 40970
rect 73592 39664 73946 40668
rect 62064 39412 73946 39664
rect 76540 39654 87156 40040
rect 76524 39596 87156 39654
rect 62064 39342 73904 39412
rect 53414 34200 53622 34564
rect 59558 34446 59684 35834
rect 59892 34446 60238 35834
rect 76524 38980 77012 39596
rect 76524 35632 76712 38980
rect 76940 35632 77012 38980
rect 79960 38974 80304 39076
rect 76524 35080 77012 35632
rect 79960 35626 80038 38974
rect 80266 35626 80304 38974
rect 83270 38974 83614 39076
rect 79960 35524 80304 35626
rect 83270 35626 83348 38974
rect 83576 35626 83614 38974
rect 86622 39284 87110 39596
rect 83270 35524 83614 35626
rect 86622 35360 86742 39284
rect 86978 35360 87110 39284
rect 86622 35184 87110 35360
rect 76524 34976 76984 35080
rect 86578 35050 87110 35184
rect 86578 34976 87096 35050
rect 76524 34680 87096 34976
rect 76614 34664 87096 34680
rect 86578 34636 87096 34664
rect 48 28672 1326 29868
rect 1420 28672 1702 29868
rect 7794 29876 8002 30038
rect 48 24032 1702 28672
rect 7794 28680 7840 29876
rect 7934 28680 8002 29876
rect 14300 29884 14508 30046
rect 7794 28316 8002 28680
rect 14300 28688 14346 29884
rect 14440 28688 14508 29884
rect 20790 29868 20998 30030
rect 14300 28324 14508 28688
rect 20790 28672 20836 29868
rect 20930 28672 20998 29868
rect 27312 29884 27520 30046
rect 20790 28308 20998 28672
rect 27312 28688 27358 29884
rect 27452 28688 27520 29884
rect 33822 29890 34030 30052
rect 27312 28324 27520 28688
rect 33822 28694 33868 29890
rect 33962 28694 34030 29890
rect 40312 29890 40520 30052
rect 33822 28330 34030 28694
rect 40312 28694 40358 29890
rect 40452 28694 40520 29890
rect 46900 29912 47108 30074
rect 40312 28330 40520 28694
rect 46900 28716 46946 29912
rect 47040 28716 47108 29912
rect 53414 29926 53622 30088
rect 46900 28352 47108 28716
rect 53414 28730 53460 29926
rect 53554 28730 53622 29926
rect 59558 29896 60238 34446
rect 53414 28366 53622 28730
rect 59558 28426 59642 29896
rect 59974 28426 60238 29896
rect 48 22836 1326 24032
rect 1420 22836 1702 24032
rect 7794 24040 8002 24202
rect 48 18168 1702 22836
rect 7794 22844 7840 24040
rect 7934 22844 8002 24040
rect 14300 24048 14508 24210
rect 7794 22480 8002 22844
rect 14300 22852 14346 24048
rect 14440 22852 14508 24048
rect 20790 24032 20998 24194
rect 14300 22488 14508 22852
rect 20790 22836 20836 24032
rect 20930 22836 20998 24032
rect 27312 24048 27520 24210
rect 20790 22472 20998 22836
rect 27312 22852 27358 24048
rect 27452 22852 27520 24048
rect 33822 24054 34030 24216
rect 27312 22488 27520 22852
rect 33822 22858 33868 24054
rect 33962 22858 34030 24054
rect 40312 24054 40520 24216
rect 33822 22494 34030 22858
rect 40312 22858 40358 24054
rect 40452 22858 40520 24054
rect 46900 24076 47108 24238
rect 40312 22494 40520 22858
rect 46900 22880 46946 24076
rect 47040 22880 47108 24076
rect 53414 24090 53622 24252
rect 46900 22516 47108 22880
rect 53414 22894 53460 24090
rect 53554 22894 53622 24090
rect 59558 24250 60238 28426
rect 60858 27536 61940 27564
rect 60858 26870 101384 27536
rect 60858 26800 101452 26870
rect 60858 26440 61940 26800
rect 53414 22530 53622 22894
rect 59558 22696 59614 24250
rect 59864 22696 60238 24250
rect 48 16972 1326 18168
rect 1420 16972 1702 18168
rect 7794 18176 8002 18338
rect 48 12312 1702 16972
rect 7794 16980 7840 18176
rect 7934 16980 8002 18176
rect 14300 18184 14508 18346
rect 7794 16616 8002 16980
rect 14300 16988 14346 18184
rect 14440 16988 14508 18184
rect 20790 18168 20998 18330
rect 14300 16624 14508 16988
rect 20790 16972 20836 18168
rect 20930 16972 20998 18168
rect 27312 18184 27520 18346
rect 20790 16608 20998 16972
rect 27312 16988 27358 18184
rect 27452 16988 27520 18184
rect 33822 18190 34030 18352
rect 27312 16624 27520 16988
rect 33822 16994 33868 18190
rect 33962 16994 34030 18190
rect 40312 18190 40520 18352
rect 33822 16630 34030 16994
rect 40312 16994 40358 18190
rect 40452 16994 40520 18190
rect 46900 18212 47108 18374
rect 40312 16630 40520 16994
rect 46900 17016 46946 18212
rect 47040 17016 47108 18212
rect 53414 18226 53622 18388
rect 46900 16652 47108 17016
rect 53414 17030 53460 18226
rect 53554 17030 53622 18226
rect 59558 18464 60238 22696
rect 53414 16666 53622 17030
rect 59558 16980 59698 18464
rect 59892 16980 60238 18464
rect 48 11116 1336 12312
rect 1430 11116 1702 12312
rect 7804 12320 8012 12482
rect 48 6404 1702 11116
rect 7804 11124 7850 12320
rect 7944 11124 8012 12320
rect 14310 12328 14518 12490
rect 7804 10760 8012 11124
rect 14310 11132 14356 12328
rect 14450 11132 14518 12328
rect 20800 12312 21008 12474
rect 14310 10768 14518 11132
rect 20800 11116 20846 12312
rect 20940 11116 21008 12312
rect 27322 12328 27530 12490
rect 20800 10752 21008 11116
rect 27322 11132 27368 12328
rect 27462 11132 27530 12328
rect 33832 12334 34040 12496
rect 27322 10768 27530 11132
rect 33832 11138 33878 12334
rect 33972 11138 34040 12334
rect 40322 12334 40530 12496
rect 33832 10774 34040 11138
rect 40322 11138 40368 12334
rect 40462 11138 40530 12334
rect 46910 12356 47118 12518
rect 40322 10774 40530 11138
rect 46910 11160 46956 12356
rect 47050 11160 47118 12356
rect 53424 12370 53632 12532
rect 46910 10796 47118 11160
rect 53424 11174 53470 12370
rect 53564 11174 53632 12370
rect 59558 12542 60238 16980
rect 53424 10810 53632 11174
rect 59558 11168 59698 12542
rect 59934 11168 60238 12542
rect 48 5208 1354 6404
rect 1448 5208 1702 6404
rect 7822 6412 8030 6574
rect 48 1284 1702 5208
rect 7822 5216 7868 6412
rect 7962 5216 8030 6412
rect 14328 6420 14536 6582
rect 7822 4852 8030 5216
rect 14328 5224 14374 6420
rect 14468 5224 14536 6420
rect 20818 6404 21026 6566
rect 14328 4860 14536 5224
rect 20818 5208 20864 6404
rect 20958 5208 21026 6404
rect 27340 6420 27548 6582
rect 20818 4844 21026 5208
rect 27340 5224 27386 6420
rect 27480 5224 27548 6420
rect 33850 6426 34058 6588
rect 27340 4860 27548 5224
rect 33850 5230 33896 6426
rect 33990 5230 34058 6426
rect 40340 6426 40548 6588
rect 33850 4866 34058 5230
rect 40340 5230 40386 6426
rect 40480 5230 40548 6426
rect 46928 6448 47136 6610
rect 40340 4866 40548 5230
rect 46928 5252 46974 6448
rect 47068 5252 47136 6448
rect 53442 6462 53650 6624
rect 46928 4888 47136 5252
rect 53442 5266 53488 6462
rect 53582 5266 53650 6462
rect 59558 6714 60238 11168
rect 53442 4902 53650 5266
rect 59558 5340 59684 6714
rect 59850 5340 60238 6714
rect 59558 1284 60238 5340
rect 60922 24034 61936 26440
rect 60922 22838 61480 24034
rect 61574 22838 61936 24034
rect 67896 24032 68104 24194
rect 60922 18196 61936 22838
rect 67896 22836 67942 24032
rect 68036 22836 68104 24032
rect 100438 25188 101452 26800
rect 74590 24006 74798 24168
rect 67896 22472 68104 22836
rect 74590 22810 74636 24006
rect 74730 22810 74798 24006
rect 81052 24004 81260 24166
rect 74590 22446 74798 22810
rect 81052 22808 81098 24004
rect 81192 22808 81260 24004
rect 87824 23998 88032 24160
rect 81052 22444 81260 22808
rect 87824 22802 87870 23998
rect 87964 22802 88032 23998
rect 94286 23996 94494 24158
rect 87824 22438 88032 22802
rect 94286 22800 94332 23996
rect 94426 22800 94494 23996
rect 94286 22436 94494 22800
rect 100438 21336 100720 25188
rect 101232 21336 101452 25188
rect 100438 19110 101452 21336
rect 60922 17000 61486 18196
rect 61580 17000 61936 18196
rect 67904 18208 68112 18370
rect 60922 12338 61936 17000
rect 67904 17012 67950 18208
rect 68044 17012 68112 18208
rect 74596 18168 74804 18330
rect 67904 16648 68112 17012
rect 74596 16972 74642 18168
rect 74736 16972 74804 18168
rect 81060 18180 81268 18342
rect 74596 16608 74804 16972
rect 81060 16984 81106 18180
rect 81200 16984 81268 18180
rect 87830 18160 88038 18322
rect 81060 16620 81268 16984
rect 87830 16964 87876 18160
rect 87970 16964 88038 18160
rect 94294 18172 94502 18334
rect 87830 16600 88038 16964
rect 94294 16976 94340 18172
rect 94434 16976 94502 18172
rect 94294 16612 94502 16976
rect 100438 14992 100698 19110
rect 101188 14992 101452 19110
rect 60922 11142 61486 12338
rect 61580 11142 61936 12338
rect 67908 12336 68116 12498
rect 60922 6480 61936 11142
rect 67908 11140 67954 12336
rect 68048 11140 68116 12336
rect 100438 13700 101452 14992
rect 74596 12310 74804 12472
rect 67908 10776 68116 11140
rect 74596 11114 74642 12310
rect 74736 11114 74804 12310
rect 81064 12308 81272 12470
rect 74596 10750 74804 11114
rect 81064 11112 81110 12308
rect 81204 11112 81272 12308
rect 87830 12302 88038 12464
rect 81064 10748 81272 11112
rect 87830 11106 87876 12302
rect 87970 11106 88038 12302
rect 94298 12300 94506 12462
rect 87830 10742 88038 11106
rect 94298 11104 94344 12300
rect 94438 11104 94506 12300
rect 94298 10740 94506 11104
rect 100438 9516 100742 13700
rect 101232 9516 101452 13700
rect 60922 5284 61486 6480
rect 61580 5284 61936 6480
rect 67912 6478 68120 6640
rect 60922 2580 61936 5284
rect 67912 5282 67958 6478
rect 68052 5282 68120 6478
rect 100438 7468 101452 9516
rect 74596 6452 74804 6614
rect 67912 4918 68120 5282
rect 74596 5256 74642 6452
rect 74736 5256 74804 6452
rect 81068 6450 81276 6612
rect 74596 4892 74804 5256
rect 81068 5254 81114 6450
rect 81208 5254 81276 6450
rect 87830 6444 88038 6606
rect 81068 4890 81276 5254
rect 87830 5248 87876 6444
rect 87970 5248 88038 6444
rect 94302 6442 94510 6604
rect 87830 4884 88038 5248
rect 94302 5246 94348 6442
rect 94442 5246 94510 6442
rect 94302 4882 94510 5246
rect 100438 3350 100786 7468
rect 101166 3350 101452 7468
rect 100438 2580 101452 3350
rect 60908 2410 101452 2580
rect 60908 1844 101434 2410
rect 48 30 60292 1284
rect 59558 0 60238 30
<< mvnsubdiff >>
rect 70886 75030 82102 75164
rect 70886 74716 82118 75030
rect 70916 74012 71230 74716
rect 42232 73732 58078 73906
rect 70916 73864 71236 74012
rect 42232 73400 42904 73732
rect 45304 73730 58078 73732
rect 45304 73400 46912 73730
rect 42232 73398 46912 73400
rect 49312 73398 50924 73730
rect 53324 73398 54934 73730
rect 57334 73398 58078 73730
rect 42232 73350 58078 73398
rect 70944 73066 71236 73864
rect 81788 74014 82118 74716
rect 70944 72042 71042 73066
rect 42720 69534 45366 69560
rect 42720 69202 42896 69534
rect 45296 69202 45366 69534
rect 42720 69158 45366 69202
rect 46714 69534 49360 69560
rect 46714 69202 46890 69534
rect 49290 69202 49360 69534
rect 46714 69158 49360 69202
rect 50736 69534 53382 69560
rect 50736 69202 50912 69534
rect 53312 69202 53382 69534
rect 50736 69158 53382 69202
rect 54758 69534 57404 69560
rect 54758 69202 54934 69534
rect 57334 69202 57404 69534
rect 54758 69158 57404 69202
rect 70952 70320 71042 72042
rect 71182 72042 71236 73066
rect 74876 73046 75092 73106
rect 71182 70320 71228 72042
rect 70952 70266 71228 70320
rect 70952 69350 71220 70266
rect 74876 70300 74906 73046
rect 75046 70300 75092 73046
rect 78726 73060 78942 73120
rect 74876 70246 75092 70300
rect 78726 70314 78756 73060
rect 78896 70314 78942 73060
rect 78726 70260 78942 70314
rect 70952 69290 71224 69350
rect 20876 66106 21098 66112
rect 222 66090 594 66106
rect 20602 66090 21098 66106
rect 222 65970 21098 66090
rect 222 65934 19500 65970
rect 222 65930 16950 65934
rect 222 65928 6370 65930
rect 222 65786 1028 65928
rect 2542 65924 6370 65928
rect 2542 65786 3696 65924
rect 222 65782 3696 65786
rect 5210 65788 6370 65924
rect 7884 65788 9016 65930
rect 10530 65924 14324 65930
rect 10530 65788 11670 65924
rect 5210 65782 11670 65788
rect 13184 65788 14324 65924
rect 15838 65792 16950 65930
rect 18464 65792 19500 65934
rect 15838 65788 19500 65792
rect 13184 65782 19500 65788
rect 222 65776 19500 65782
rect 20566 65776 21098 65970
rect 222 65734 21098 65776
rect 70952 66544 71038 69290
rect 71178 66544 71224 69290
rect 74872 69270 75088 69330
rect 70952 66490 71224 66544
rect 222 57816 594 65734
rect 19392 65726 21098 65734
rect 19392 65724 20628 65726
rect 19364 59702 20600 59726
rect 944 59660 2556 59684
rect 944 59518 1000 59660
rect 2514 59518 2556 59660
rect 944 59490 2556 59518
rect 3612 59656 5224 59680
rect 3612 59514 3668 59656
rect 5182 59514 5224 59656
rect 3612 59486 5224 59514
rect 6286 59662 7898 59686
rect 6286 59520 6342 59662
rect 7856 59520 7898 59662
rect 6286 59492 7898 59520
rect 8932 59662 10544 59686
rect 8932 59520 8988 59662
rect 10502 59520 10544 59662
rect 8932 59492 10544 59520
rect 11586 59656 13198 59680
rect 11586 59514 11642 59656
rect 13156 59514 13198 59656
rect 11586 59486 13198 59514
rect 14240 59662 15852 59686
rect 14240 59520 14296 59662
rect 15810 59520 15852 59662
rect 14240 59492 15852 59520
rect 16866 59666 18478 59690
rect 16866 59524 16922 59666
rect 18436 59524 18478 59666
rect 16866 59496 18478 59524
rect 19364 59508 19472 59702
rect 20538 59508 20600 59702
rect 19364 59456 20600 59508
rect 222 56666 280 57816
rect 496 56666 594 57816
rect 222 47480 594 56666
rect 19364 53336 20600 53360
rect 944 53294 2556 53318
rect 944 53152 1000 53294
rect 2514 53152 2556 53294
rect 944 53124 2556 53152
rect 3612 53290 5224 53314
rect 3612 53148 3668 53290
rect 5182 53148 5224 53290
rect 3612 53120 5224 53148
rect 6286 53296 7898 53320
rect 6286 53154 6342 53296
rect 7856 53154 7898 53296
rect 6286 53126 7898 53154
rect 8932 53296 10544 53320
rect 8932 53154 8988 53296
rect 10502 53154 10544 53296
rect 8932 53126 10544 53154
rect 11586 53290 13198 53314
rect 11586 53148 11642 53290
rect 13156 53148 13198 53290
rect 11586 53120 13198 53148
rect 14240 53296 15852 53320
rect 14240 53154 14296 53296
rect 15810 53154 15852 53296
rect 14240 53126 15852 53154
rect 16866 53300 18478 53324
rect 16866 53158 16922 53300
rect 18436 53158 18478 53300
rect 16866 53130 18478 53158
rect 19364 53142 19472 53336
rect 20538 53142 20600 53336
rect 19364 53090 20600 53142
rect 20876 47480 21098 65726
rect 70952 65580 71220 66490
rect 74872 66524 74902 69270
rect 75042 66524 75088 69270
rect 78722 69284 78938 69344
rect 74872 66470 75088 66524
rect 78722 66538 78752 69284
rect 78892 66538 78938 69284
rect 78722 66484 78938 66538
rect 70952 65520 71224 65580
rect 42708 65060 45354 65086
rect 42708 64728 42884 65060
rect 45284 64728 45354 65060
rect 42708 64684 45354 64728
rect 46716 65058 49362 65084
rect 46716 64726 46892 65058
rect 49292 64726 49362 65058
rect 46716 64682 49362 64726
rect 50728 65058 53374 65084
rect 50728 64726 50904 65058
rect 53304 64726 53374 65058
rect 50728 64682 53374 64726
rect 54738 65058 57384 65084
rect 70952 65062 71038 65520
rect 54738 64726 54914 65058
rect 57314 64726 57384 65058
rect 54738 64682 57384 64726
rect 70960 62774 71038 65062
rect 71178 65070 71224 65520
rect 74872 65500 75088 65560
rect 71178 62774 71228 65070
rect 70960 61756 71228 62774
rect 74872 62754 74902 65500
rect 75042 62754 75088 65500
rect 78722 65514 78938 65574
rect 74872 62700 75088 62754
rect 78722 62768 78752 65514
rect 78892 62768 78938 65514
rect 78722 62714 78938 62768
rect 42700 60862 45346 60888
rect 42700 60530 42876 60862
rect 45276 60530 45346 60862
rect 42700 60486 45346 60530
rect 46694 60862 49340 60888
rect 46694 60530 46870 60862
rect 49270 60530 49340 60862
rect 46694 60486 49340 60530
rect 50716 60862 53362 60888
rect 50716 60530 50892 60862
rect 53292 60530 53362 60862
rect 50716 60486 53362 60530
rect 54738 60862 57384 60888
rect 54738 60530 54914 60862
rect 57314 60530 57384 60862
rect 54738 60486 57384 60530
rect 70960 59010 71038 61756
rect 71178 59010 71228 61756
rect 74872 61736 75088 61796
rect 70960 57980 71228 59010
rect 74872 58990 74902 61736
rect 75042 58990 75088 61736
rect 78722 61750 78938 61810
rect 74872 58936 75088 58990
rect 78722 59004 78752 61750
rect 78892 59004 78938 61750
rect 78722 58950 78938 59004
rect 42652 56472 45298 56498
rect 42652 56140 42828 56472
rect 45228 56140 45298 56472
rect 42652 56096 45298 56140
rect 46660 56470 49306 56496
rect 46660 56138 46836 56470
rect 49236 56138 49306 56470
rect 46660 56094 49306 56138
rect 50672 56470 53318 56496
rect 50672 56138 50848 56470
rect 53248 56138 53318 56470
rect 50672 56094 53318 56138
rect 54682 56470 57328 56496
rect 54682 56138 54858 56470
rect 57258 56138 57328 56470
rect 54682 56094 57328 56138
rect 70960 55234 71038 57980
rect 71178 55234 71228 57980
rect 74872 57960 75088 58020
rect 70960 54208 71228 55234
rect 74872 55214 74902 57960
rect 75042 55214 75088 57960
rect 78722 57974 78938 58034
rect 74872 55160 75088 55214
rect 78722 55228 78752 57974
rect 78892 55228 78938 57974
rect 78722 55174 78938 55228
rect 81818 54936 82118 74014
rect 42644 52274 45290 52300
rect 42644 51942 42820 52274
rect 45220 51942 45290 52274
rect 42644 51898 45290 51942
rect 46638 52274 49284 52300
rect 46638 51942 46814 52274
rect 49214 51942 49284 52274
rect 46638 51898 49284 51942
rect 50660 52274 53306 52300
rect 50660 51942 50836 52274
rect 53236 51942 53306 52274
rect 50660 51898 53306 51942
rect 54682 52274 57328 52300
rect 54682 51942 54858 52274
rect 57258 51942 57328 52274
rect 54682 51898 57328 51942
rect 70960 51462 71042 54208
rect 71182 51462 71228 54208
rect 74876 54188 75092 54248
rect 70960 51342 71228 51462
rect 70946 51064 71228 51342
rect 74876 51442 74906 54188
rect 75046 51442 75092 54188
rect 78726 54202 78942 54262
rect 74876 51388 75092 51442
rect 78726 51456 78756 54202
rect 78896 51456 78942 54202
rect 81818 54182 81910 54936
rect 82086 54182 82118 54936
rect 78726 51402 78942 51456
rect 81818 51268 82118 54182
rect 83272 54065 83303 54099
rect 83337 54065 83399 54099
rect 83433 54065 83495 54099
rect 83529 54065 83591 54099
rect 83625 54065 83687 54099
rect 83721 54065 83783 54099
rect 83817 54065 83879 54099
rect 83913 54065 83975 54099
rect 84009 54065 84071 54099
rect 84105 54065 84167 54099
rect 84201 54065 84263 54099
rect 84297 54065 84359 54099
rect 84393 54065 84455 54099
rect 84489 54065 84551 54099
rect 84585 54065 84647 54099
rect 84681 54065 84743 54099
rect 84777 54065 84839 54099
rect 84873 54065 84935 54099
rect 84969 54065 85031 54099
rect 85065 54065 85127 54099
rect 85161 54065 85223 54099
rect 85257 54065 85319 54099
rect 85353 54065 85415 54099
rect 85449 54065 85511 54099
rect 85545 54065 85607 54099
rect 85641 54065 85703 54099
rect 85737 54065 85799 54099
rect 85833 54065 85895 54099
rect 85929 54065 85991 54099
rect 86025 54065 86087 54099
rect 86121 54065 86183 54099
rect 86217 54065 86279 54099
rect 86313 54065 86344 54099
rect 70946 50626 71214 51064
rect 81818 50626 82148 51268
rect 70916 50192 82148 50626
rect 70916 50162 82088 50192
rect 42092 48178 57938 48310
rect 42092 48166 46660 48178
rect 42092 47902 42766 48166
rect 44904 47914 46660 48166
rect 49352 48152 57938 48178
rect 49352 48140 54448 48152
rect 49352 47914 50790 48140
rect 53312 47928 54448 48140
rect 57206 47928 57938 48152
rect 53312 47914 57938 47928
rect 44904 47902 57938 47914
rect 42092 47754 57938 47902
rect 222 47408 21098 47480
rect 222 47404 17048 47408
rect 222 47370 9118 47404
rect 222 47240 2592 47370
rect 4384 47244 9118 47370
rect 10578 47386 17048 47404
rect 10578 47244 14218 47386
rect 4384 47240 14218 47244
rect 222 47226 14218 47240
rect 15628 47262 17048 47386
rect 18368 47378 21098 47408
rect 18368 47262 19456 47378
rect 15628 47226 19456 47262
rect 222 47222 19456 47226
rect 20474 47222 21098 47378
rect 222 47116 21098 47222
rect 222 47114 594 47116
<< mvpsubdiffcont >>
rect 24368 55766 25098 55868
rect 28714 55872 29532 55970
rect 22980 54924 23102 55346
rect 24374 53876 25104 53978
rect 28720 53982 29538 54080
rect 28736 52040 29554 52138
rect 24390 51934 25120 52036
rect 83303 53251 83337 53285
rect 83399 53251 83433 53285
rect 83495 53251 83529 53285
rect 83591 53251 83625 53285
rect 83687 53251 83721 53285
rect 83783 53251 83817 53285
rect 83879 53251 83913 53285
rect 83975 53251 84009 53285
rect 84071 53251 84105 53285
rect 84167 53251 84201 53285
rect 84263 53251 84297 53285
rect 84359 53251 84393 53285
rect 84455 53251 84489 53285
rect 84551 53251 84585 53285
rect 84647 53251 84681 53285
rect 84743 53251 84777 53285
rect 84839 53251 84873 53285
rect 84935 53251 84969 53285
rect 85031 53251 85065 53285
rect 85127 53251 85161 53285
rect 85223 53251 85257 53285
rect 85319 53251 85353 53285
rect 85415 53251 85449 53285
rect 85511 53251 85545 53285
rect 85607 53251 85641 53285
rect 85703 53251 85737 53285
rect 85799 53251 85833 53285
rect 85895 53251 85929 53285
rect 85991 53251 86025 53285
rect 86087 53251 86121 53285
rect 86183 53251 86217 53285
rect 86279 53251 86313 53285
rect 24240 44696 25328 44998
rect 38946 44424 42360 45148
rect 1326 40322 1420 41518
rect 7840 40330 7934 41526
rect 14346 40338 14440 41534
rect 20836 40322 20930 41518
rect 27358 40338 27452 41534
rect 33868 40344 33962 41540
rect 40358 40344 40452 41540
rect 46946 40366 47040 41562
rect 53460 40380 53554 41576
rect 68330 43808 68980 43950
rect 59572 40204 59836 41772
rect 1326 34506 1420 35702
rect 7840 34514 7934 35710
rect 14346 34522 14440 35718
rect 20836 34506 20930 35702
rect 27358 34522 27452 35718
rect 33868 34528 33962 35724
rect 40358 34528 40452 35724
rect 46946 34550 47040 35746
rect 53460 34564 53554 35760
rect 62180 40876 62328 42630
rect 65974 40878 66122 42632
rect 69782 40892 69930 42646
rect 73646 40970 73876 42876
rect 59684 34446 59892 35834
rect 76712 35632 76940 38980
rect 80038 35626 80266 38974
rect 83348 35626 83576 38974
rect 86742 35360 86978 39284
rect 1326 28672 1420 29868
rect 7840 28680 7934 29876
rect 14346 28688 14440 29884
rect 20836 28672 20930 29868
rect 27358 28688 27452 29884
rect 33868 28694 33962 29890
rect 40358 28694 40452 29890
rect 46946 28716 47040 29912
rect 53460 28730 53554 29926
rect 59642 28426 59974 29896
rect 1326 22836 1420 24032
rect 7840 22844 7934 24040
rect 14346 22852 14440 24048
rect 20836 22836 20930 24032
rect 27358 22852 27452 24048
rect 33868 22858 33962 24054
rect 40358 22858 40452 24054
rect 46946 22880 47040 24076
rect 53460 22894 53554 24090
rect 59614 22696 59864 24250
rect 1326 16972 1420 18168
rect 7840 16980 7934 18176
rect 14346 16988 14440 18184
rect 20836 16972 20930 18168
rect 27358 16988 27452 18184
rect 33868 16994 33962 18190
rect 40358 16994 40452 18190
rect 46946 17016 47040 18212
rect 53460 17030 53554 18226
rect 59698 16980 59892 18464
rect 1336 11116 1430 12312
rect 7850 11124 7944 12320
rect 14356 11132 14450 12328
rect 20846 11116 20940 12312
rect 27368 11132 27462 12328
rect 33878 11138 33972 12334
rect 40368 11138 40462 12334
rect 46956 11160 47050 12356
rect 53470 11174 53564 12370
rect 59698 11168 59934 12542
rect 1354 5208 1448 6404
rect 7868 5216 7962 6412
rect 14374 5224 14468 6420
rect 20864 5208 20958 6404
rect 27386 5224 27480 6420
rect 33896 5230 33990 6426
rect 40386 5230 40480 6426
rect 46974 5252 47068 6448
rect 53488 5266 53582 6462
rect 59684 5340 59850 6714
rect 61480 22838 61574 24034
rect 67942 22836 68036 24032
rect 74636 22810 74730 24006
rect 81098 22808 81192 24004
rect 87870 22802 87964 23998
rect 94332 22800 94426 23996
rect 100720 21336 101232 25188
rect 61486 17000 61580 18196
rect 67950 17012 68044 18208
rect 74642 16972 74736 18168
rect 81106 16984 81200 18180
rect 87876 16964 87970 18160
rect 94340 16976 94434 18172
rect 100698 14992 101188 19110
rect 61486 11142 61580 12338
rect 67954 11140 68048 12336
rect 74642 11114 74736 12310
rect 81110 11112 81204 12308
rect 87876 11106 87970 12302
rect 94344 11104 94438 12300
rect 100742 9516 101232 13700
rect 61486 5284 61580 6480
rect 67958 5282 68052 6478
rect 74642 5256 74736 6452
rect 81114 5254 81208 6450
rect 87876 5248 87970 6444
rect 94348 5246 94442 6442
rect 100786 3350 101166 7468
<< mvnsubdiffcont >>
rect 42904 73400 45304 73732
rect 46912 73398 49312 73730
rect 50924 73398 53324 73730
rect 54934 73398 57334 73730
rect 42896 69202 45296 69534
rect 46890 69202 49290 69534
rect 50912 69202 53312 69534
rect 54934 69202 57334 69534
rect 71042 70320 71182 73066
rect 74906 70300 75046 73046
rect 78756 70314 78896 73060
rect 1028 65786 2542 65928
rect 3696 65782 5210 65924
rect 6370 65788 7884 65930
rect 9016 65788 10530 65930
rect 11670 65782 13184 65924
rect 14324 65788 15838 65930
rect 16950 65792 18464 65934
rect 19500 65776 20566 65970
rect 71038 66544 71178 69290
rect 1000 59518 2514 59660
rect 3668 59514 5182 59656
rect 6342 59520 7856 59662
rect 8988 59520 10502 59662
rect 11642 59514 13156 59656
rect 14296 59520 15810 59662
rect 16922 59524 18436 59666
rect 19472 59508 20538 59702
rect 280 56666 496 57816
rect 1000 53152 2514 53294
rect 3668 53148 5182 53290
rect 6342 53154 7856 53296
rect 8988 53154 10502 53296
rect 11642 53148 13156 53290
rect 14296 53154 15810 53296
rect 16922 53158 18436 53300
rect 19472 53142 20538 53336
rect 74902 66524 75042 69270
rect 78752 66538 78892 69284
rect 42884 64728 45284 65060
rect 46892 64726 49292 65058
rect 50904 64726 53304 65058
rect 54914 64726 57314 65058
rect 71038 62774 71178 65520
rect 74902 62754 75042 65500
rect 78752 62768 78892 65514
rect 42876 60530 45276 60862
rect 46870 60530 49270 60862
rect 50892 60530 53292 60862
rect 54914 60530 57314 60862
rect 71038 59010 71178 61756
rect 74902 58990 75042 61736
rect 78752 59004 78892 61750
rect 42828 56140 45228 56472
rect 46836 56138 49236 56470
rect 50848 56138 53248 56470
rect 54858 56138 57258 56470
rect 71038 55234 71178 57980
rect 74902 55214 75042 57960
rect 78752 55228 78892 57974
rect 42820 51942 45220 52274
rect 46814 51942 49214 52274
rect 50836 51942 53236 52274
rect 54858 51942 57258 52274
rect 71042 51462 71182 54208
rect 74906 51442 75046 54188
rect 78756 51456 78896 54202
rect 81910 54182 82086 54936
rect 83303 54065 83337 54099
rect 83399 54065 83433 54099
rect 83495 54065 83529 54099
rect 83591 54065 83625 54099
rect 83687 54065 83721 54099
rect 83783 54065 83817 54099
rect 83879 54065 83913 54099
rect 83975 54065 84009 54099
rect 84071 54065 84105 54099
rect 84167 54065 84201 54099
rect 84263 54065 84297 54099
rect 84359 54065 84393 54099
rect 84455 54065 84489 54099
rect 84551 54065 84585 54099
rect 84647 54065 84681 54099
rect 84743 54065 84777 54099
rect 84839 54065 84873 54099
rect 84935 54065 84969 54099
rect 85031 54065 85065 54099
rect 85127 54065 85161 54099
rect 85223 54065 85257 54099
rect 85319 54065 85353 54099
rect 85415 54065 85449 54099
rect 85511 54065 85545 54099
rect 85607 54065 85641 54099
rect 85703 54065 85737 54099
rect 85799 54065 85833 54099
rect 85895 54065 85929 54099
rect 85991 54065 86025 54099
rect 86087 54065 86121 54099
rect 86183 54065 86217 54099
rect 86279 54065 86313 54099
rect 42766 47902 44904 48166
rect 46660 47914 49352 48178
rect 50790 47914 53312 48140
rect 54448 47928 57206 48152
rect 2592 47240 4384 47370
rect 9118 47244 10578 47404
rect 14218 47226 15628 47386
rect 17048 47262 18368 47408
rect 19456 47222 20474 47378
<< poly >>
rect 79978 74590 81316 74624
rect 72226 74496 73396 74538
rect 72226 74372 72590 74496
rect 71844 74370 72590 74372
rect 72878 74372 73396 74496
rect 79978 74406 80390 74590
rect 80836 74406 81316 74590
rect 72878 74370 73774 74372
rect 71844 74280 73774 74370
rect 79978 74366 81316 74406
rect 71384 74274 73958 74280
rect 71384 74254 71984 74274
rect 72042 74254 72642 74274
rect 72700 74254 73300 74274
rect 73358 74254 73958 74274
rect 75708 74260 77638 74352
rect 79558 74274 81488 74366
rect 79098 74268 81672 74274
rect 75248 74254 77822 74260
rect 42170 72582 42196 73182
rect 42796 73104 42822 73182
rect 42864 73104 42890 73182
rect 42796 72664 42890 73104
rect 42796 72582 42822 72664
rect 42864 72582 42890 72664
rect 43490 73102 43516 73182
rect 43558 73102 43584 73182
rect 43490 72662 43584 73102
rect 43490 72582 43516 72662
rect 43558 72582 43584 72662
rect 44184 73116 44210 73182
rect 44252 73116 44278 73182
rect 44184 72676 44278 73116
rect 44184 72582 44210 72676
rect 44252 72582 44278 72676
rect 44878 73096 44904 73182
rect 44946 73096 44972 73182
rect 44878 72650 44972 73096
rect 44878 72582 44904 72650
rect 44946 72582 44972 72650
rect 45572 72936 45598 73182
rect 45572 72912 45660 72936
rect 46178 72912 46204 73180
rect 45572 72678 46204 72912
rect 45572 72582 45660 72678
rect 45590 72524 45660 72582
rect 46178 72580 46204 72678
rect 46804 73102 46830 73180
rect 46872 73102 46898 73180
rect 46804 72662 46898 73102
rect 46804 72580 46830 72662
rect 46872 72580 46898 72662
rect 47498 73100 47524 73180
rect 47566 73100 47592 73180
rect 47498 72660 47592 73100
rect 47498 72580 47524 72660
rect 47566 72580 47592 72660
rect 48192 73114 48218 73180
rect 48260 73114 48286 73180
rect 48192 72674 48286 73114
rect 48192 72580 48218 72674
rect 48260 72580 48286 72674
rect 48886 73094 48912 73180
rect 48954 73094 48980 73180
rect 48886 72648 48980 73094
rect 48886 72580 48912 72648
rect 48954 72580 48980 72648
rect 49580 72934 49606 73180
rect 49580 72916 49668 72934
rect 50190 72916 50216 73180
rect 49580 72682 50216 72916
rect 49580 72580 49668 72682
rect 50190 72580 50216 72682
rect 50816 73102 50842 73180
rect 50884 73102 50910 73180
rect 50816 72662 50910 73102
rect 50816 72580 50842 72662
rect 50884 72580 50910 72662
rect 51510 73100 51536 73180
rect 51578 73100 51604 73180
rect 51510 72660 51604 73100
rect 51510 72580 51536 72660
rect 51578 72580 51604 72660
rect 52204 73114 52230 73180
rect 52272 73114 52298 73180
rect 52204 72674 52298 73114
rect 52204 72580 52230 72674
rect 52272 72580 52298 72674
rect 52898 73094 52924 73180
rect 52966 73094 52992 73180
rect 52898 72648 52992 73094
rect 52898 72580 52924 72648
rect 52966 72580 52992 72648
rect 53592 72934 53618 73180
rect 53592 72906 53680 72934
rect 54200 72906 54226 73180
rect 53592 72672 54226 72906
rect 53592 72580 53680 72672
rect 54200 72580 54226 72672
rect 54826 73102 54852 73180
rect 54894 73102 54920 73180
rect 54826 72662 54920 73102
rect 54826 72580 54852 72662
rect 54894 72580 54920 72662
rect 55520 73100 55546 73180
rect 55588 73100 55614 73180
rect 55520 72660 55614 73100
rect 55520 72580 55546 72660
rect 55588 72580 55614 72660
rect 56214 73114 56240 73180
rect 56282 73114 56308 73180
rect 56214 72674 56308 73114
rect 56214 72580 56240 72674
rect 56282 72580 56308 72674
rect 56908 73094 56934 73180
rect 56976 73094 57002 73180
rect 56908 72648 57002 73094
rect 56908 72580 56934 72648
rect 56976 72580 57002 72648
rect 57602 72934 57628 73180
rect 75248 74234 75848 74254
rect 75906 74234 76506 74254
rect 76564 74234 77164 74254
rect 77222 74234 77822 74254
rect 79098 74248 79698 74268
rect 79756 74248 80356 74268
rect 80414 74248 81014 74268
rect 81072 74248 81672 74268
rect 71384 73628 71984 73654
rect 72042 73628 72642 73654
rect 72700 73628 73300 73654
rect 73358 73628 73958 73654
rect 71714 73432 71792 73628
rect 72162 73432 72240 73628
rect 72910 73432 72982 73628
rect 73462 73432 73534 73628
rect 75248 73608 75848 73634
rect 75906 73608 76506 73634
rect 76564 73608 77164 73634
rect 77222 73608 77822 73634
rect 79098 73622 79698 73648
rect 79756 73622 80356 73648
rect 80414 73622 81014 73648
rect 81072 73622 81672 73648
rect 71702 73366 73792 73432
rect 75578 73412 75656 73608
rect 76026 73412 76104 73608
rect 76774 73412 76846 73608
rect 77326 73412 77398 73608
rect 79428 73426 79506 73622
rect 79876 73426 79954 73622
rect 80624 73426 80696 73622
rect 81176 73426 81248 73622
rect 71356 73362 73930 73366
rect 71356 73340 71956 73362
rect 72014 73340 72614 73362
rect 72672 73340 73272 73362
rect 73330 73340 73930 73362
rect 75566 73346 77656 73412
rect 79416 73360 81506 73426
rect 79070 73356 81644 73360
rect 75220 73342 77794 73346
rect 57602 72580 57690 72934
rect 42170 71924 42196 72524
rect 42796 72434 42822 72524
rect 42864 72434 42890 72524
rect 42796 71994 42890 72434
rect 42796 71924 42822 71994
rect 42864 71924 42890 71994
rect 43490 72458 43516 72524
rect 43558 72458 43584 72524
rect 43490 72018 43584 72458
rect 43490 71924 43516 72018
rect 43558 71924 43584 72018
rect 44184 72442 44210 72524
rect 44252 72442 44278 72524
rect 44184 72002 44278 72442
rect 44184 71924 44210 72002
rect 44252 71924 44278 72002
rect 44878 72454 44904 72524
rect 44946 72454 44972 72524
rect 44878 72014 44972 72454
rect 44878 71924 44904 72014
rect 44946 71924 44972 72014
rect 45572 72406 45660 72524
rect 49598 72522 49668 72580
rect 53610 72522 53680 72580
rect 57620 72522 57690 72580
rect 46178 72406 46204 72522
rect 45572 72172 46204 72406
rect 45572 71924 45660 72172
rect 45590 71866 45660 71924
rect 46178 71922 46204 72172
rect 46804 72432 46830 72522
rect 46872 72432 46898 72522
rect 46804 71992 46898 72432
rect 46804 71922 46830 71992
rect 46872 71922 46898 71992
rect 47498 72456 47524 72522
rect 47566 72456 47592 72522
rect 47498 72016 47592 72456
rect 47498 71922 47524 72016
rect 47566 71922 47592 72016
rect 48192 72440 48218 72522
rect 48260 72440 48286 72522
rect 48192 72000 48286 72440
rect 48192 71922 48218 72000
rect 48260 71922 48286 72000
rect 48886 72452 48912 72522
rect 48954 72452 48980 72522
rect 48886 72012 48980 72452
rect 48886 71922 48912 72012
rect 48954 71922 48980 72012
rect 49580 72406 49668 72522
rect 50190 72406 50216 72522
rect 49580 72172 50216 72406
rect 49580 71922 49668 72172
rect 50190 71922 50216 72172
rect 50816 72432 50842 72522
rect 50884 72432 50910 72522
rect 50816 71992 50910 72432
rect 50816 71922 50842 71992
rect 50884 71922 50910 71992
rect 51510 72456 51536 72522
rect 51578 72456 51604 72522
rect 51510 72016 51604 72456
rect 51510 71922 51536 72016
rect 51578 71922 51604 72016
rect 52204 72440 52230 72522
rect 52272 72440 52298 72522
rect 52204 72000 52298 72440
rect 52204 71922 52230 72000
rect 52272 71922 52298 72000
rect 52898 72452 52924 72522
rect 52966 72452 52992 72522
rect 52898 72012 52992 72452
rect 52898 71922 52924 72012
rect 52966 71922 52992 72012
rect 53592 72448 53680 72522
rect 54200 72448 54226 72522
rect 53592 72214 54226 72448
rect 53592 71922 53680 72214
rect 54200 71922 54226 72214
rect 54826 72432 54852 72522
rect 54894 72432 54920 72522
rect 54826 71992 54920 72432
rect 54826 71922 54852 71992
rect 54894 71922 54920 71992
rect 55520 72456 55546 72522
rect 55588 72456 55614 72522
rect 55520 72016 55614 72456
rect 55520 71922 55546 72016
rect 55588 71922 55614 72016
rect 56214 72440 56240 72522
rect 56282 72440 56308 72522
rect 56214 72000 56308 72440
rect 56214 71922 56240 72000
rect 56282 71922 56308 72000
rect 56908 72452 56934 72522
rect 56976 72452 57002 72522
rect 56908 72012 57002 72452
rect 56908 71922 56934 72012
rect 56976 71922 57002 72012
rect 57602 71922 57690 72522
rect 42170 71266 42196 71866
rect 42796 71758 42822 71866
rect 42864 71758 42890 71866
rect 42796 71318 42890 71758
rect 42796 71266 42822 71318
rect 42864 71266 42890 71318
rect 43490 71770 43516 71866
rect 43558 71770 43584 71866
rect 43490 71330 43584 71770
rect 43490 71266 43516 71330
rect 43558 71266 43584 71330
rect 44184 71748 44210 71866
rect 44252 71748 44278 71866
rect 44184 71308 44278 71748
rect 44184 71266 44210 71308
rect 44252 71266 44278 71308
rect 44878 71720 44904 71866
rect 44946 71720 44972 71866
rect 44878 71280 44972 71720
rect 44878 71266 44904 71280
rect 44946 71266 44972 71280
rect 45572 71728 45660 71866
rect 49598 71864 49668 71922
rect 53610 71864 53680 71922
rect 57620 71864 57690 71922
rect 46178 71728 46204 71864
rect 45572 71494 46204 71728
rect 45572 71266 45660 71494
rect 45590 71208 45660 71266
rect 46178 71264 46204 71494
rect 46804 71756 46830 71864
rect 46872 71756 46898 71864
rect 46804 71316 46898 71756
rect 46804 71264 46830 71316
rect 46872 71264 46898 71316
rect 47498 71768 47524 71864
rect 47566 71768 47592 71864
rect 47498 71328 47592 71768
rect 47498 71264 47524 71328
rect 47566 71264 47592 71328
rect 48192 71746 48218 71864
rect 48260 71746 48286 71864
rect 48192 71306 48286 71746
rect 48192 71264 48218 71306
rect 48260 71264 48286 71306
rect 48886 71718 48912 71864
rect 48954 71718 48980 71864
rect 48886 71278 48980 71718
rect 48886 71264 48912 71278
rect 48954 71264 48980 71278
rect 49580 71734 49668 71864
rect 50190 71734 50216 71864
rect 49580 71500 50216 71734
rect 49580 71264 49668 71500
rect 50190 71264 50216 71500
rect 50816 71756 50842 71864
rect 50884 71756 50910 71864
rect 50816 71316 50910 71756
rect 50816 71264 50842 71316
rect 50884 71264 50910 71316
rect 51510 71768 51536 71864
rect 51578 71768 51604 71864
rect 51510 71328 51604 71768
rect 51510 71264 51536 71328
rect 51578 71264 51604 71328
rect 52204 71746 52230 71864
rect 52272 71746 52298 71864
rect 52204 71306 52298 71746
rect 52204 71264 52230 71306
rect 52272 71264 52298 71306
rect 52898 71718 52924 71864
rect 52966 71718 52992 71864
rect 52898 71278 52992 71718
rect 52898 71264 52924 71278
rect 52966 71264 52992 71278
rect 53592 71718 53680 71864
rect 54200 71718 54226 71864
rect 53592 71484 54226 71718
rect 53592 71264 53680 71484
rect 54200 71264 54226 71484
rect 54826 71756 54852 71864
rect 54894 71756 54920 71864
rect 54826 71316 54920 71756
rect 54826 71264 54852 71316
rect 54894 71264 54920 71316
rect 55520 71768 55546 71864
rect 55588 71768 55614 71864
rect 55520 71328 55614 71768
rect 55520 71264 55546 71328
rect 55588 71264 55614 71328
rect 56214 71746 56240 71864
rect 56282 71746 56308 71864
rect 56214 71306 56308 71746
rect 56214 71264 56240 71306
rect 56282 71264 56308 71306
rect 56908 71718 56934 71864
rect 56976 71718 57002 71864
rect 56908 71278 57002 71718
rect 56908 71264 56934 71278
rect 56976 71264 57002 71278
rect 57602 71264 57690 71864
rect 42170 70608 42196 71208
rect 42796 71126 42822 71208
rect 42864 71126 42890 71208
rect 42796 70686 42890 71126
rect 42796 70608 42822 70686
rect 42864 70608 42890 70686
rect 43490 71148 43516 71208
rect 43558 71148 43584 71208
rect 43490 70708 43584 71148
rect 43490 70608 43516 70708
rect 43558 70608 43584 70708
rect 44184 71148 44210 71208
rect 44252 71148 44278 71208
rect 44184 70708 44278 71148
rect 44184 70608 44210 70708
rect 44252 70608 44278 70708
rect 44878 71136 44904 71208
rect 44946 71136 44972 71208
rect 44878 70696 44972 71136
rect 44878 70608 44904 70696
rect 44946 70608 44972 70696
rect 45572 71126 45660 71208
rect 49598 71206 49668 71264
rect 53610 71206 53680 71264
rect 57620 71206 57690 71264
rect 46178 71126 46204 71206
rect 45572 70892 46204 71126
rect 45572 70608 45660 70892
rect 45590 70550 45660 70608
rect 46178 70606 46204 70892
rect 46804 71124 46830 71206
rect 46872 71124 46898 71206
rect 46804 70684 46898 71124
rect 46804 70606 46830 70684
rect 46872 70606 46898 70684
rect 47498 71146 47524 71206
rect 47566 71146 47592 71206
rect 47498 70706 47592 71146
rect 47498 70606 47524 70706
rect 47566 70606 47592 70706
rect 48192 71146 48218 71206
rect 48260 71146 48286 71206
rect 48192 70706 48286 71146
rect 48192 70606 48218 70706
rect 48260 70606 48286 70706
rect 48886 71134 48912 71206
rect 48954 71134 48980 71206
rect 48886 70694 48980 71134
rect 48886 70606 48912 70694
rect 48954 70606 48980 70694
rect 49580 71092 49668 71206
rect 50190 71092 50216 71206
rect 49580 70858 50216 71092
rect 49580 70606 49668 70858
rect 50190 70606 50216 70858
rect 50816 71124 50842 71206
rect 50884 71124 50910 71206
rect 50816 70684 50910 71124
rect 50816 70606 50842 70684
rect 50884 70606 50910 70684
rect 51510 71146 51536 71206
rect 51578 71146 51604 71206
rect 51510 70706 51604 71146
rect 51510 70606 51536 70706
rect 51578 70606 51604 70706
rect 52204 71146 52230 71206
rect 52272 71146 52298 71206
rect 52204 70706 52298 71146
rect 52204 70606 52230 70706
rect 52272 70606 52298 70706
rect 52898 71134 52924 71206
rect 52966 71134 52992 71206
rect 52898 70694 52992 71134
rect 52898 70606 52924 70694
rect 52966 70606 52992 70694
rect 53592 71116 53680 71206
rect 54200 71116 54226 71206
rect 53592 70882 54226 71116
rect 53592 70606 53680 70882
rect 54200 70606 54226 70882
rect 54826 71124 54852 71206
rect 54894 71124 54920 71206
rect 54826 70684 54920 71124
rect 54826 70606 54852 70684
rect 54894 70606 54920 70684
rect 55520 71146 55546 71206
rect 55588 71146 55614 71206
rect 55520 70706 55614 71146
rect 55520 70606 55546 70706
rect 55588 70606 55614 70706
rect 56214 71146 56240 71206
rect 56282 71146 56308 71206
rect 56214 70706 56308 71146
rect 56214 70606 56240 70706
rect 56282 70606 56308 70706
rect 56908 71134 56934 71206
rect 56976 71134 57002 71206
rect 56908 70694 57002 71134
rect 56908 70606 56934 70694
rect 56976 70606 57002 70694
rect 57602 70624 57690 71206
rect 57602 70606 57880 70624
rect 42170 69950 42196 70550
rect 42796 70418 42822 70550
rect 42864 70418 42890 70550
rect 42796 69978 42890 70418
rect 42796 69950 42822 69978
rect 42864 69950 42890 69978
rect 43490 70460 43516 70550
rect 43558 70460 43584 70550
rect 43490 70020 43584 70460
rect 43490 69950 43516 70020
rect 43558 69950 43584 70020
rect 44184 70472 44210 70550
rect 44252 70472 44278 70550
rect 44184 70032 44278 70472
rect 44184 69950 44210 70032
rect 44252 69950 44278 70032
rect 44878 70498 44904 70550
rect 44946 70498 44972 70550
rect 44878 70058 44972 70498
rect 44878 69950 44904 70058
rect 44946 69950 44972 70058
rect 45572 70524 45660 70550
rect 49598 70548 49668 70606
rect 53610 70548 53680 70606
rect 57620 70548 57880 70606
rect 46178 70524 46204 70548
rect 45572 70290 46204 70524
rect 45572 70270 45660 70290
rect 45572 69950 45598 70270
rect 46178 69948 46204 70290
rect 46804 70416 46830 70548
rect 46872 70416 46898 70548
rect 46804 69976 46898 70416
rect 46804 69948 46830 69976
rect 46872 69948 46898 69976
rect 47498 70458 47524 70548
rect 47566 70458 47592 70548
rect 47498 70018 47592 70458
rect 47498 69948 47524 70018
rect 47566 69948 47592 70018
rect 48192 70470 48218 70548
rect 48260 70470 48286 70548
rect 48192 70030 48286 70470
rect 48192 69948 48218 70030
rect 48260 69948 48286 70030
rect 48886 70496 48912 70548
rect 48954 70496 48980 70548
rect 48886 70056 48980 70496
rect 48886 69948 48912 70056
rect 48954 69948 48980 70056
rect 49580 70500 49668 70548
rect 50190 70500 50216 70548
rect 49580 70266 50216 70500
rect 49580 69948 49606 70266
rect 50190 69948 50216 70266
rect 50816 70416 50842 70548
rect 50884 70416 50910 70548
rect 50816 69976 50910 70416
rect 50816 69948 50842 69976
rect 50884 69948 50910 69976
rect 51510 70458 51536 70548
rect 51578 70458 51604 70548
rect 51510 70018 51604 70458
rect 51510 69948 51536 70018
rect 51578 69948 51604 70018
rect 52204 70470 52230 70548
rect 52272 70470 52298 70548
rect 52204 70030 52298 70470
rect 52204 69948 52230 70030
rect 52272 69948 52298 70030
rect 52898 70496 52924 70548
rect 52966 70496 52992 70548
rect 52898 70056 52992 70496
rect 52898 69948 52924 70056
rect 52966 69948 52992 70056
rect 53592 70544 53680 70548
rect 54200 70544 54226 70548
rect 53592 70310 54226 70544
rect 53592 70268 53680 70310
rect 53592 69948 53618 70268
rect 54200 69948 54226 70310
rect 54826 70416 54852 70548
rect 54894 70416 54920 70548
rect 54826 69976 54920 70416
rect 54826 69948 54852 69976
rect 54894 69948 54920 69976
rect 55520 70458 55546 70548
rect 55588 70458 55614 70548
rect 55520 70018 55614 70458
rect 55520 69948 55546 70018
rect 55588 69948 55614 70018
rect 56214 70470 56240 70548
rect 56282 70470 56308 70548
rect 56214 70030 56308 70470
rect 56214 69948 56240 70030
rect 56282 69948 56308 70030
rect 56908 70496 56934 70548
rect 56976 70496 57002 70548
rect 56908 70056 57002 70496
rect 56908 69948 56934 70056
rect 56976 69948 57002 70056
rect 57602 70268 57880 70548
rect 57602 69948 57628 70268
rect 57678 69722 57880 70268
rect 57678 69438 57710 69722
rect 57854 69438 57880 69722
rect 42162 68384 42188 68984
rect 42788 68906 42814 68984
rect 42856 68906 42882 68984
rect 42788 68466 42882 68906
rect 42788 68384 42814 68466
rect 42856 68384 42882 68466
rect 43482 68904 43508 68984
rect 43550 68904 43576 68984
rect 43482 68464 43576 68904
rect 43482 68384 43508 68464
rect 43550 68384 43576 68464
rect 44176 68918 44202 68984
rect 44244 68918 44270 68984
rect 44176 68478 44270 68918
rect 44176 68384 44202 68478
rect 44244 68384 44270 68478
rect 44870 68898 44896 68984
rect 44938 68898 44964 68984
rect 44870 68452 44964 68898
rect 44870 68384 44896 68452
rect 44938 68384 44964 68452
rect 45564 68738 45590 68984
rect 45564 68702 45652 68738
rect 46156 68702 46182 68984
rect 45564 68466 46182 68702
rect 45564 68384 45652 68466
rect 46156 68384 46182 68466
rect 46782 68906 46808 68984
rect 46850 68906 46876 68984
rect 46782 68466 46876 68906
rect 46782 68384 46808 68466
rect 46850 68384 46876 68466
rect 47476 68904 47502 68984
rect 47544 68904 47570 68984
rect 47476 68464 47570 68904
rect 47476 68384 47502 68464
rect 47544 68384 47570 68464
rect 48170 68918 48196 68984
rect 48238 68918 48264 68984
rect 48170 68478 48264 68918
rect 48170 68384 48196 68478
rect 48238 68384 48264 68478
rect 48864 68898 48890 68984
rect 48932 68898 48958 68984
rect 48864 68452 48958 68898
rect 48864 68384 48890 68452
rect 48932 68384 48958 68452
rect 49558 68738 49584 68984
rect 49558 68698 49646 68738
rect 50178 68698 50204 68984
rect 49558 68462 50204 68698
rect 49558 68384 49646 68462
rect 50178 68384 50204 68462
rect 50804 68906 50830 68984
rect 50872 68906 50898 68984
rect 50804 68466 50898 68906
rect 50804 68384 50830 68466
rect 50872 68384 50898 68466
rect 51498 68904 51524 68984
rect 51566 68904 51592 68984
rect 51498 68464 51592 68904
rect 51498 68384 51524 68464
rect 51566 68384 51592 68464
rect 52192 68918 52218 68984
rect 52260 68918 52286 68984
rect 52192 68478 52286 68918
rect 52192 68384 52218 68478
rect 52260 68384 52286 68478
rect 52886 68898 52912 68984
rect 52954 68898 52980 68984
rect 52886 68452 52980 68898
rect 52886 68384 52912 68452
rect 52954 68384 52980 68452
rect 53580 68738 53606 68984
rect 53580 68698 53668 68738
rect 54200 68698 54226 68984
rect 53580 68462 54226 68698
rect 53580 68384 53668 68462
rect 54200 68384 54226 68462
rect 54826 68906 54852 68984
rect 54894 68906 54920 68984
rect 54826 68466 54920 68906
rect 54826 68384 54852 68466
rect 54894 68384 54920 68466
rect 55520 68904 55546 68984
rect 55588 68904 55614 68984
rect 55520 68464 55614 68904
rect 55520 68384 55546 68464
rect 55588 68384 55614 68464
rect 56214 68918 56240 68984
rect 56282 68918 56308 68984
rect 56214 68478 56308 68918
rect 56214 68384 56240 68478
rect 56282 68384 56308 68478
rect 56908 68898 56934 68984
rect 56976 68898 57002 68984
rect 56908 68452 57002 68898
rect 56908 68384 56934 68452
rect 56976 68384 57002 68452
rect 57602 68738 57628 68984
rect 57678 68738 57880 69438
rect 57602 68506 57880 68738
rect 75220 73320 75820 73342
rect 75878 73320 76478 73342
rect 76536 73320 77136 73342
rect 77194 73320 77794 73342
rect 79070 73334 79670 73356
rect 79728 73334 80328 73356
rect 80386 73334 80986 73356
rect 81044 73334 81644 73356
rect 71356 72714 71956 72740
rect 72014 72714 72614 72740
rect 72672 72714 73272 72740
rect 73330 72714 73930 72740
rect 71416 72672 71840 72714
rect 72154 72672 72578 72714
rect 72736 72672 73160 72714
rect 73408 72672 73832 72714
rect 71356 72646 71956 72672
rect 72014 72646 72614 72672
rect 72672 72646 73272 72672
rect 73330 72646 73930 72672
rect 71356 72020 71956 72046
rect 72014 72020 72614 72046
rect 72672 72020 73272 72046
rect 73330 72020 73930 72046
rect 71410 71978 71834 72020
rect 72122 71978 72546 72020
rect 72732 71978 73156 72020
rect 73448 71978 73872 72020
rect 71356 71952 71956 71978
rect 72014 71952 72614 71978
rect 72672 71952 73272 71978
rect 73330 71952 73930 71978
rect 71356 71326 71956 71352
rect 72014 71326 72614 71352
rect 72672 71326 73272 71352
rect 73330 71326 73930 71352
rect 71396 71284 71820 71326
rect 72142 71284 72566 71326
rect 72770 71284 73194 71326
rect 73406 71284 73830 71326
rect 71356 71258 71956 71284
rect 72014 71258 72614 71284
rect 72672 71258 73272 71284
rect 73330 71258 73930 71284
rect 71356 70632 71956 70658
rect 72014 70632 72614 70658
rect 72672 70632 73272 70658
rect 73330 70632 73930 70658
rect 71392 70590 71816 70632
rect 72172 70590 72596 70632
rect 72722 70590 73146 70632
rect 73440 70590 73864 70632
rect 71356 70564 71956 70590
rect 72014 70564 72614 70590
rect 72672 70564 73272 70590
rect 73330 70564 73930 70590
rect 75220 72694 75820 72720
rect 75878 72694 76478 72720
rect 76536 72694 77136 72720
rect 77194 72694 77794 72720
rect 75280 72652 75704 72694
rect 76018 72652 76442 72694
rect 76600 72652 77024 72694
rect 77272 72652 77696 72694
rect 75220 72626 75820 72652
rect 75878 72626 76478 72652
rect 76536 72626 77136 72652
rect 77194 72626 77794 72652
rect 75220 72000 75820 72026
rect 75878 72000 76478 72026
rect 76536 72000 77136 72026
rect 77194 72000 77794 72026
rect 75274 71958 75698 72000
rect 75986 71958 76410 72000
rect 76596 71958 77020 72000
rect 77312 71958 77736 72000
rect 75220 71932 75820 71958
rect 75878 71932 76478 71958
rect 76536 71932 77136 71958
rect 77194 71932 77794 71958
rect 75220 71306 75820 71332
rect 75878 71306 76478 71332
rect 76536 71306 77136 71332
rect 77194 71306 77794 71332
rect 75260 71264 75684 71306
rect 76006 71264 76430 71306
rect 76634 71264 77058 71306
rect 77270 71264 77694 71306
rect 75220 71238 75820 71264
rect 75878 71238 76478 71264
rect 76536 71238 77136 71264
rect 77194 71238 77794 71264
rect 75220 70612 75820 70638
rect 75878 70612 76478 70638
rect 76536 70612 77136 70638
rect 77194 70612 77794 70638
rect 75256 70570 75680 70612
rect 76036 70570 76460 70612
rect 76586 70570 77010 70612
rect 77304 70570 77728 70612
rect 75220 70544 75820 70570
rect 75878 70544 76478 70570
rect 76536 70544 77136 70570
rect 77194 70544 77794 70570
rect 71356 69938 71956 69964
rect 72014 69938 72614 69964
rect 72672 69938 73272 69964
rect 73330 69938 73930 69964
rect 79070 72708 79670 72734
rect 79728 72708 80328 72734
rect 80386 72708 80986 72734
rect 81044 72708 81644 72734
rect 79130 72666 79554 72708
rect 79868 72666 80292 72708
rect 80450 72666 80874 72708
rect 81122 72666 81546 72708
rect 79070 72640 79670 72666
rect 79728 72640 80328 72666
rect 80386 72640 80986 72666
rect 81044 72640 81644 72666
rect 79070 72014 79670 72040
rect 79728 72014 80328 72040
rect 80386 72014 80986 72040
rect 81044 72014 81644 72040
rect 79124 71972 79548 72014
rect 79836 71972 80260 72014
rect 80446 71972 80870 72014
rect 81162 71972 81586 72014
rect 79070 71946 79670 71972
rect 79728 71946 80328 71972
rect 80386 71946 80986 71972
rect 81044 71946 81644 71972
rect 79070 71320 79670 71346
rect 79728 71320 80328 71346
rect 80386 71320 80986 71346
rect 81044 71320 81644 71346
rect 79110 71278 79534 71320
rect 79856 71278 80280 71320
rect 80484 71278 80908 71320
rect 81120 71278 81544 71320
rect 79070 71252 79670 71278
rect 79728 71252 80328 71278
rect 80386 71252 80986 71278
rect 81044 71252 81644 71278
rect 79070 70626 79670 70652
rect 79728 70626 80328 70652
rect 80386 70626 80986 70652
rect 81044 70626 81644 70652
rect 79106 70584 79530 70626
rect 79886 70584 80310 70626
rect 80436 70584 80860 70626
rect 81154 70584 81578 70626
rect 79070 70558 79670 70584
rect 79728 70558 80328 70584
rect 80386 70558 80986 70584
rect 81044 70558 81644 70584
rect 71718 69656 71824 69938
rect 72126 69656 72232 69938
rect 72834 69656 72940 69938
rect 73436 69656 73542 69938
rect 75220 69918 75820 69944
rect 75878 69918 76478 69944
rect 76536 69918 77136 69944
rect 77194 69918 77794 69944
rect 79070 69932 79670 69958
rect 79728 69932 80328 69958
rect 80386 69932 80986 69958
rect 81044 69932 81644 69958
rect 71698 69590 73788 69656
rect 75582 69636 75688 69918
rect 75990 69636 76096 69918
rect 76698 69636 76804 69918
rect 77300 69636 77406 69918
rect 79432 69650 79538 69932
rect 79840 69650 79946 69932
rect 80548 69650 80654 69932
rect 81150 69650 81256 69932
rect 71352 69586 73926 69590
rect 71352 69564 71952 69586
rect 72010 69564 72610 69586
rect 72668 69564 73268 69586
rect 73326 69564 73926 69586
rect 75562 69570 77652 69636
rect 79412 69584 81502 69650
rect 79066 69580 81640 69584
rect 75216 69566 77790 69570
rect 57602 68384 57690 68506
rect 45582 68326 45652 68384
rect 49576 68326 49646 68384
rect 53598 68326 53668 68384
rect 57620 68326 57690 68384
rect 42162 67726 42188 68326
rect 42788 68236 42814 68326
rect 42856 68236 42882 68326
rect 42788 67796 42882 68236
rect 42788 67726 42814 67796
rect 42856 67726 42882 67796
rect 43482 68260 43508 68326
rect 43550 68260 43576 68326
rect 43482 67820 43576 68260
rect 43482 67726 43508 67820
rect 43550 67726 43576 67820
rect 44176 68244 44202 68326
rect 44244 68244 44270 68326
rect 44176 67804 44270 68244
rect 44176 67726 44202 67804
rect 44244 67726 44270 67804
rect 44870 68256 44896 68326
rect 44938 68256 44964 68326
rect 44870 67816 44964 68256
rect 44870 67726 44896 67816
rect 44938 67726 44964 67816
rect 45564 68206 45652 68326
rect 46156 68206 46182 68326
rect 45564 67970 46182 68206
rect 45564 67726 45652 67970
rect 46156 67726 46182 67970
rect 46782 68236 46808 68326
rect 46850 68236 46876 68326
rect 46782 67796 46876 68236
rect 46782 67726 46808 67796
rect 46850 67726 46876 67796
rect 47476 68260 47502 68326
rect 47544 68260 47570 68326
rect 47476 67820 47570 68260
rect 47476 67726 47502 67820
rect 47544 67726 47570 67820
rect 48170 68244 48196 68326
rect 48238 68244 48264 68326
rect 48170 67804 48264 68244
rect 48170 67726 48196 67804
rect 48238 67726 48264 67804
rect 48864 68256 48890 68326
rect 48932 68256 48958 68326
rect 48864 67816 48958 68256
rect 48864 67726 48890 67816
rect 48932 67726 48958 67816
rect 49558 68166 49646 68326
rect 50178 68166 50204 68326
rect 49558 67930 50204 68166
rect 49558 67726 49646 67930
rect 50178 67726 50204 67930
rect 50804 68236 50830 68326
rect 50872 68236 50898 68326
rect 50804 67796 50898 68236
rect 50804 67726 50830 67796
rect 50872 67726 50898 67796
rect 51498 68260 51524 68326
rect 51566 68260 51592 68326
rect 51498 67820 51592 68260
rect 51498 67726 51524 67820
rect 51566 67726 51592 67820
rect 52192 68244 52218 68326
rect 52260 68244 52286 68326
rect 52192 67804 52286 68244
rect 52192 67726 52218 67804
rect 52260 67726 52286 67804
rect 52886 68256 52912 68326
rect 52954 68256 52980 68326
rect 52886 67816 52980 68256
rect 52886 67726 52912 67816
rect 52954 67726 52980 67816
rect 53580 68176 53668 68326
rect 54200 68176 54226 68326
rect 53580 67940 54226 68176
rect 53580 67726 53668 67940
rect 54200 67726 54226 67940
rect 54826 68236 54852 68326
rect 54894 68236 54920 68326
rect 54826 67796 54920 68236
rect 54826 67726 54852 67796
rect 54894 67726 54920 67796
rect 55520 68260 55546 68326
rect 55588 68260 55614 68326
rect 55520 67820 55614 68260
rect 55520 67726 55546 67820
rect 55588 67726 55614 67820
rect 56214 68244 56240 68326
rect 56282 68244 56308 68326
rect 56214 67804 56308 68244
rect 56214 67726 56240 67804
rect 56282 67726 56308 67804
rect 56908 68256 56934 68326
rect 56976 68256 57002 68326
rect 56908 67816 57002 68256
rect 56908 67726 56934 67816
rect 56976 67726 57002 67816
rect 57602 67726 57690 68326
rect 45582 67668 45652 67726
rect 49576 67668 49646 67726
rect 53598 67668 53668 67726
rect 57620 67668 57690 67726
rect 42162 67068 42188 67668
rect 42788 67560 42814 67668
rect 42856 67560 42882 67668
rect 42788 67120 42882 67560
rect 42788 67068 42814 67120
rect 42856 67068 42882 67120
rect 43482 67572 43508 67668
rect 43550 67572 43576 67668
rect 43482 67132 43576 67572
rect 43482 67068 43508 67132
rect 43550 67068 43576 67132
rect 44176 67550 44202 67668
rect 44244 67550 44270 67668
rect 44176 67110 44270 67550
rect 44176 67068 44202 67110
rect 44244 67068 44270 67110
rect 44870 67522 44896 67668
rect 44938 67522 44964 67668
rect 44870 67082 44964 67522
rect 44870 67068 44896 67082
rect 44938 67068 44964 67082
rect 45564 67526 45652 67668
rect 46156 67526 46182 67668
rect 45564 67290 46182 67526
rect 45564 67068 45652 67290
rect 46156 67068 46182 67290
rect 46782 67560 46808 67668
rect 46850 67560 46876 67668
rect 46782 67120 46876 67560
rect 46782 67068 46808 67120
rect 46850 67068 46876 67120
rect 47476 67572 47502 67668
rect 47544 67572 47570 67668
rect 47476 67132 47570 67572
rect 47476 67068 47502 67132
rect 47544 67068 47570 67132
rect 48170 67550 48196 67668
rect 48238 67550 48264 67668
rect 48170 67110 48264 67550
rect 48170 67068 48196 67110
rect 48238 67068 48264 67110
rect 48864 67522 48890 67668
rect 48932 67522 48958 67668
rect 48864 67082 48958 67522
rect 48864 67068 48890 67082
rect 48932 67068 48958 67082
rect 49558 67474 49646 67668
rect 50178 67474 50204 67668
rect 49558 67238 50204 67474
rect 49558 67068 49646 67238
rect 50178 67068 50204 67238
rect 50804 67560 50830 67668
rect 50872 67560 50898 67668
rect 50804 67120 50898 67560
rect 50804 67068 50830 67120
rect 50872 67068 50898 67120
rect 51498 67572 51524 67668
rect 51566 67572 51592 67668
rect 51498 67132 51592 67572
rect 51498 67068 51524 67132
rect 51566 67068 51592 67132
rect 52192 67550 52218 67668
rect 52260 67550 52286 67668
rect 52192 67110 52286 67550
rect 52192 67068 52218 67110
rect 52260 67068 52286 67110
rect 52886 67522 52912 67668
rect 52954 67522 52980 67668
rect 52886 67082 52980 67522
rect 52886 67068 52912 67082
rect 52954 67068 52980 67082
rect 53580 67526 53668 67668
rect 54200 67526 54226 67668
rect 53580 67290 54226 67526
rect 53580 67068 53668 67290
rect 54200 67068 54226 67290
rect 54826 67560 54852 67668
rect 54894 67560 54920 67668
rect 54826 67120 54920 67560
rect 54826 67068 54852 67120
rect 54894 67068 54920 67120
rect 55520 67572 55546 67668
rect 55588 67572 55614 67668
rect 55520 67132 55614 67572
rect 55520 67068 55546 67132
rect 55588 67068 55614 67132
rect 56214 67550 56240 67668
rect 56282 67550 56308 67668
rect 56214 67110 56308 67550
rect 56214 67068 56240 67110
rect 56282 67068 56308 67110
rect 56908 67522 56934 67668
rect 56976 67522 57002 67668
rect 56908 67082 57002 67522
rect 56908 67068 56934 67082
rect 56976 67068 57002 67082
rect 57602 67068 57690 67668
rect 45582 67010 45652 67068
rect 49576 67010 49646 67068
rect 53598 67010 53668 67068
rect 57620 67010 57690 67068
rect 42162 66410 42188 67010
rect 42788 66928 42814 67010
rect 42856 66928 42882 67010
rect 42788 66488 42882 66928
rect 42788 66410 42814 66488
rect 42856 66410 42882 66488
rect 43482 66950 43508 67010
rect 43550 66950 43576 67010
rect 43482 66510 43576 66950
rect 43482 66410 43508 66510
rect 43550 66410 43576 66510
rect 44176 66950 44202 67010
rect 44244 66950 44270 67010
rect 44176 66510 44270 66950
rect 44176 66410 44202 66510
rect 44244 66410 44270 66510
rect 44870 66938 44896 67010
rect 44938 66938 44964 67010
rect 44870 66498 44964 66938
rect 44870 66410 44896 66498
rect 44938 66410 44964 66498
rect 45564 66832 45652 67010
rect 46156 66832 46182 67010
rect 45564 66596 46182 66832
rect 45564 66410 45652 66596
rect 46156 66410 46182 66596
rect 46782 66928 46808 67010
rect 46850 66928 46876 67010
rect 46782 66488 46876 66928
rect 46782 66410 46808 66488
rect 46850 66410 46876 66488
rect 47476 66950 47502 67010
rect 47544 66950 47570 67010
rect 47476 66510 47570 66950
rect 47476 66410 47502 66510
rect 47544 66410 47570 66510
rect 48170 66950 48196 67010
rect 48238 66950 48264 67010
rect 48170 66510 48264 66950
rect 48170 66410 48196 66510
rect 48238 66410 48264 66510
rect 48864 66938 48890 67010
rect 48932 66938 48958 67010
rect 48864 66498 48958 66938
rect 48864 66410 48890 66498
rect 48932 66410 48958 66498
rect 49558 66832 49646 67010
rect 50178 66832 50204 67010
rect 49558 66596 50204 66832
rect 49558 66410 49646 66596
rect 50178 66410 50204 66596
rect 50804 66928 50830 67010
rect 50872 66928 50898 67010
rect 50804 66488 50898 66928
rect 50804 66410 50830 66488
rect 50872 66410 50898 66488
rect 51498 66950 51524 67010
rect 51566 66950 51592 67010
rect 51498 66510 51592 66950
rect 51498 66410 51524 66510
rect 51566 66410 51592 66510
rect 52192 66950 52218 67010
rect 52260 66950 52286 67010
rect 52192 66510 52286 66950
rect 52192 66410 52218 66510
rect 52260 66410 52286 66510
rect 52886 66938 52912 67010
rect 52954 66938 52980 67010
rect 52886 66498 52980 66938
rect 52886 66410 52912 66498
rect 52954 66410 52980 66498
rect 53580 66938 53668 67010
rect 54200 66938 54226 67010
rect 53580 66702 54226 66938
rect 53580 66410 53668 66702
rect 54200 66410 54226 66702
rect 54826 66928 54852 67010
rect 54894 66928 54920 67010
rect 54826 66488 54920 66928
rect 54826 66410 54852 66488
rect 54894 66410 54920 66488
rect 55520 66950 55546 67010
rect 55588 66950 55614 67010
rect 55520 66510 55614 66950
rect 55520 66410 55546 66510
rect 55588 66410 55614 66510
rect 56214 66950 56240 67010
rect 56282 66950 56308 67010
rect 56214 66510 56308 66950
rect 56214 66410 56240 66510
rect 56282 66410 56308 66510
rect 56908 66938 56934 67010
rect 56976 66938 57002 67010
rect 56908 66498 57002 66938
rect 56908 66410 56934 66498
rect 56976 66410 57002 66498
rect 57602 66410 57690 67010
rect 45582 66352 45652 66410
rect 49576 66352 49646 66410
rect 53598 66352 53668 66410
rect 57620 66352 57690 66410
rect 42162 65752 42188 66352
rect 42788 66220 42814 66352
rect 42856 66220 42882 66352
rect 42788 65780 42882 66220
rect 42788 65752 42814 65780
rect 42856 65752 42882 65780
rect 43482 66262 43508 66352
rect 43550 66262 43576 66352
rect 43482 65822 43576 66262
rect 43482 65752 43508 65822
rect 43550 65752 43576 65822
rect 44176 66274 44202 66352
rect 44244 66274 44270 66352
rect 44176 65834 44270 66274
rect 44176 65752 44202 65834
rect 44244 65752 44270 65834
rect 44870 66300 44896 66352
rect 44938 66300 44964 66352
rect 44870 65860 44964 66300
rect 44870 65752 44896 65860
rect 44938 65752 44964 65860
rect 45564 66322 45652 66352
rect 46156 66322 46182 66352
rect 45564 66086 46182 66322
rect 45564 66072 45652 66086
rect 45564 65752 45590 66072
rect 46156 65752 46182 66086
rect 46782 66220 46808 66352
rect 46850 66220 46876 66352
rect 46782 65780 46876 66220
rect 46782 65752 46808 65780
rect 46850 65752 46876 65780
rect 47476 66262 47502 66352
rect 47544 66262 47570 66352
rect 47476 65822 47570 66262
rect 47476 65752 47502 65822
rect 47544 65752 47570 65822
rect 48170 66274 48196 66352
rect 48238 66274 48264 66352
rect 48170 65834 48264 66274
rect 48170 65752 48196 65834
rect 48238 65752 48264 65834
rect 48864 66300 48890 66352
rect 48932 66300 48958 66352
rect 48864 65860 48958 66300
rect 48864 65752 48890 65860
rect 48932 65752 48958 65860
rect 49558 66306 49646 66352
rect 50178 66306 50204 66352
rect 49558 66070 50204 66306
rect 49558 65752 49584 66070
rect 50178 65752 50204 66070
rect 50804 66220 50830 66352
rect 50872 66220 50898 66352
rect 50804 65780 50898 66220
rect 50804 65752 50830 65780
rect 50872 65752 50898 65780
rect 51498 66262 51524 66352
rect 51566 66262 51592 66352
rect 51498 65822 51592 66262
rect 51498 65752 51524 65822
rect 51566 65752 51592 65822
rect 52192 66274 52218 66352
rect 52260 66274 52286 66352
rect 52192 65834 52286 66274
rect 52192 65752 52218 65834
rect 52260 65752 52286 65834
rect 52886 66300 52912 66352
rect 52954 66300 52980 66352
rect 52886 65860 52980 66300
rect 52886 65752 52912 65860
rect 52954 65752 52980 65860
rect 53580 66336 53668 66352
rect 54200 66336 54226 66352
rect 53580 66100 54226 66336
rect 53580 66072 53668 66100
rect 53580 65752 53606 66072
rect 54200 65752 54226 66100
rect 54826 66220 54852 66352
rect 54894 66220 54920 66352
rect 54826 65780 54920 66220
rect 54826 65752 54852 65780
rect 54894 65752 54920 65780
rect 55520 66262 55546 66352
rect 55588 66262 55614 66352
rect 55520 65822 55614 66262
rect 55520 65752 55546 65822
rect 55588 65752 55614 65822
rect 56214 66274 56240 66352
rect 56282 66274 56308 66352
rect 56214 65834 56308 66274
rect 56214 65752 56240 65834
rect 56282 65752 56308 65834
rect 56908 66300 56934 66352
rect 56976 66300 57002 66352
rect 56908 65860 57002 66300
rect 56908 65752 56934 65860
rect 56976 65752 57002 65860
rect 57602 66072 57690 66352
rect 75216 69544 75816 69566
rect 75874 69544 76474 69566
rect 76532 69544 77132 69566
rect 77190 69544 77790 69566
rect 79066 69558 79666 69580
rect 79724 69558 80324 69580
rect 80382 69558 80982 69580
rect 81040 69558 81640 69580
rect 71352 68938 71952 68964
rect 72010 68938 72610 68964
rect 72668 68938 73268 68964
rect 73326 68938 73926 68964
rect 71412 68896 71836 68938
rect 72150 68896 72574 68938
rect 72732 68896 73156 68938
rect 73404 68896 73828 68938
rect 71352 68870 71952 68896
rect 72010 68870 72610 68896
rect 72668 68870 73268 68896
rect 73326 68870 73926 68896
rect 71352 68244 71952 68270
rect 72010 68244 72610 68270
rect 72668 68244 73268 68270
rect 73326 68244 73926 68270
rect 71406 68202 71830 68244
rect 72118 68202 72542 68244
rect 72728 68202 73152 68244
rect 73444 68202 73868 68244
rect 71352 68176 71952 68202
rect 72010 68176 72610 68202
rect 72668 68176 73268 68202
rect 73326 68176 73926 68202
rect 71352 67550 71952 67576
rect 72010 67550 72610 67576
rect 72668 67550 73268 67576
rect 73326 67550 73926 67576
rect 71392 67508 71816 67550
rect 72138 67508 72562 67550
rect 72766 67508 73190 67550
rect 73402 67508 73826 67550
rect 71352 67482 71952 67508
rect 72010 67482 72610 67508
rect 72668 67482 73268 67508
rect 73326 67482 73926 67508
rect 71352 66856 71952 66882
rect 72010 66856 72610 66882
rect 72668 66856 73268 66882
rect 73326 66856 73926 66882
rect 71388 66814 71812 66856
rect 72168 66814 72592 66856
rect 72718 66814 73142 66856
rect 73436 66814 73860 66856
rect 71352 66788 71952 66814
rect 72010 66788 72610 66814
rect 72668 66788 73268 66814
rect 73326 66788 73926 66814
rect 57602 65752 57628 66072
rect 726 64924 752 65524
rect 1352 65428 1378 65524
rect 1420 65428 1446 65524
rect 1352 65060 1446 65428
rect 1352 64924 1378 65060
rect 1420 64924 1446 65060
rect 2046 65434 2072 65524
rect 2114 65434 2140 65524
rect 2046 65066 2140 65434
rect 2046 64924 2072 65066
rect 2114 64924 2140 65066
rect 2740 65150 2766 65524
rect 2740 65128 2792 65150
rect 3394 65128 3420 65520
rect 2740 64984 3420 65128
rect 2740 64924 2792 64984
rect 2762 64866 2792 64924
rect 3394 64920 3420 64984
rect 4020 65424 4046 65520
rect 4088 65424 4114 65520
rect 4020 65056 4114 65424
rect 4020 64920 4046 65056
rect 4088 64920 4114 65056
rect 4714 65430 4740 65520
rect 4782 65430 4808 65520
rect 4714 65062 4808 65430
rect 4714 64920 4740 65062
rect 4782 64920 4808 65062
rect 5408 65146 5434 65520
rect 5408 65126 5460 65146
rect 6068 65126 6094 65526
rect 5408 64982 6094 65126
rect 5408 64920 5460 64982
rect 6068 64926 6094 64982
rect 6694 65430 6720 65526
rect 6762 65430 6788 65526
rect 6694 65062 6788 65430
rect 6694 64926 6720 65062
rect 6762 64926 6788 65062
rect 7388 65436 7414 65526
rect 7456 65436 7482 65526
rect 7388 65068 7482 65436
rect 7388 64926 7414 65068
rect 7456 64926 7482 65068
rect 8082 65430 8108 65526
rect 8082 65166 8142 65430
rect 8714 65166 8740 65526
rect 8082 64996 8740 65166
rect 8082 64926 8134 64996
rect 8714 64926 8740 64996
rect 9340 65430 9366 65526
rect 9408 65430 9434 65526
rect 9340 65062 9434 65430
rect 9340 64926 9366 65062
rect 9408 64926 9434 65062
rect 10034 65436 10060 65526
rect 10102 65436 10128 65526
rect 10034 65068 10128 65436
rect 10034 64926 10060 65068
rect 10102 64926 10128 65068
rect 10728 65518 10754 65526
rect 10728 65368 10792 65518
rect 11368 65368 11394 65520
rect 10728 65190 11394 65368
rect 10728 65120 10792 65190
rect 10728 64926 10780 65120
rect 726 64266 752 64866
rect 1352 64752 1378 64866
rect 1420 64752 1446 64866
rect 1352 64384 1446 64752
rect 1352 64266 1378 64384
rect 1420 64266 1446 64384
rect 2046 64748 2072 64866
rect 2114 64748 2140 64866
rect 2046 64380 2140 64748
rect 2046 64266 2072 64380
rect 2114 64266 2140 64380
rect 2740 64728 2792 64866
rect 5430 64862 5460 64920
rect 8104 64868 8134 64926
rect 10750 64868 10780 64926
rect 11368 64920 11394 65190
rect 11994 65424 12020 65520
rect 12062 65424 12088 65520
rect 11994 65056 12088 65424
rect 11994 64920 12020 65056
rect 12062 64920 12088 65056
rect 12688 65430 12714 65520
rect 12756 65430 12782 65520
rect 12688 65062 12782 65430
rect 12688 64920 12714 65062
rect 12756 64920 12782 65062
rect 13382 65148 13408 65520
rect 14022 65148 14048 65526
rect 13382 64970 14048 65148
rect 13382 64920 13434 64970
rect 14022 64926 14048 64970
rect 14648 65430 14674 65526
rect 14716 65430 14742 65526
rect 14648 65062 14742 65430
rect 14648 64926 14674 65062
rect 14716 64926 14742 65062
rect 15342 65436 15368 65526
rect 15410 65436 15436 65526
rect 15342 65068 15436 65436
rect 15342 64926 15368 65068
rect 15410 64926 15436 65068
rect 16036 65152 16062 65526
rect 16036 65148 16088 65152
rect 16648 65148 16674 65530
rect 16036 64990 16674 65148
rect 16036 64926 16088 64990
rect 16648 64930 16674 64990
rect 17274 65434 17300 65530
rect 17342 65434 17368 65530
rect 17274 65066 17368 65434
rect 17274 64930 17300 65066
rect 17342 64930 17368 65066
rect 17968 65440 17994 65530
rect 18036 65440 18062 65530
rect 17968 65072 18062 65440
rect 17968 64930 17994 65072
rect 18036 64930 18062 65072
rect 18662 65160 18688 65530
rect 19332 65160 19358 65574
rect 18662 65024 19358 65160
rect 18662 64930 18714 65024
rect 19332 64974 19358 65024
rect 19958 65462 19984 65574
rect 20026 65462 20052 65574
rect 19958 65090 20052 65462
rect 19958 64974 19984 65090
rect 20026 64974 20052 65090
rect 20652 65192 20678 65574
rect 20652 64974 20758 65192
rect 3394 64728 3420 64862
rect 2740 64584 3420 64728
rect 2740 64266 2792 64584
rect 2762 64208 2792 64266
rect 3394 64262 3420 64584
rect 4020 64748 4046 64862
rect 4088 64748 4114 64862
rect 4020 64380 4114 64748
rect 4020 64262 4046 64380
rect 4088 64262 4114 64380
rect 4714 64744 4740 64862
rect 4782 64744 4808 64862
rect 4714 64376 4808 64744
rect 4714 64262 4740 64376
rect 4782 64262 4808 64376
rect 5408 64632 5460 64862
rect 6068 64632 6094 64868
rect 5408 64488 6094 64632
rect 5408 64262 5460 64488
rect 6068 64268 6094 64488
rect 6694 64754 6720 64868
rect 6762 64754 6788 64868
rect 6694 64386 6788 64754
rect 6694 64268 6720 64386
rect 6762 64268 6788 64386
rect 7388 64750 7414 64868
rect 7456 64750 7482 64868
rect 7388 64382 7482 64750
rect 7388 64268 7414 64382
rect 7456 64268 7482 64382
rect 8082 64666 8134 64868
rect 8714 64666 8740 64868
rect 8082 64496 8740 64666
rect 8082 64268 8134 64496
rect 8714 64268 8740 64496
rect 9340 64754 9366 64868
rect 9408 64754 9434 64868
rect 9340 64386 9434 64754
rect 9340 64268 9366 64386
rect 9408 64268 9434 64386
rect 10034 64750 10060 64868
rect 10102 64750 10128 64868
rect 10034 64382 10128 64750
rect 10034 64268 10060 64382
rect 10102 64268 10128 64382
rect 10728 64712 10780 64868
rect 13404 64862 13434 64920
rect 16058 64868 16088 64926
rect 18684 64872 18714 64930
rect 20672 64916 20758 64974
rect 11368 64712 11394 64862
rect 10728 64534 11394 64712
rect 10728 64268 10780 64534
rect 726 63608 752 64208
rect 1352 64090 1378 64208
rect 1420 64090 1446 64208
rect 1352 63722 1446 64090
rect 1352 63608 1378 63722
rect 1420 63608 1446 63722
rect 2046 64136 2072 64208
rect 2114 64136 2140 64208
rect 2046 63768 2140 64136
rect 2046 63608 2072 63768
rect 2114 63608 2140 63768
rect 2740 63982 2792 64208
rect 5430 64204 5460 64262
rect 8104 64210 8134 64268
rect 10750 64210 10780 64268
rect 11368 64262 11394 64534
rect 11994 64748 12020 64862
rect 12062 64748 12088 64862
rect 11994 64380 12088 64748
rect 11994 64262 12020 64380
rect 12062 64262 12088 64380
rect 12688 64744 12714 64862
rect 12756 64744 12782 64862
rect 12688 64376 12782 64744
rect 12688 64262 12714 64376
rect 12756 64262 12782 64376
rect 13382 64742 13434 64862
rect 14022 64742 14048 64868
rect 13382 64564 14048 64742
rect 13382 64262 13434 64564
rect 14022 64268 14048 64564
rect 14648 64754 14674 64868
rect 14716 64754 14742 64868
rect 14648 64386 14742 64754
rect 14648 64268 14674 64386
rect 14716 64268 14742 64386
rect 15342 64750 15368 64868
rect 15410 64750 15436 64868
rect 15342 64382 15436 64750
rect 15342 64268 15368 64382
rect 15410 64268 15436 64382
rect 16036 64722 16088 64868
rect 16648 64722 16674 64872
rect 16036 64564 16674 64722
rect 16036 64268 16088 64564
rect 16648 64272 16674 64564
rect 17274 64758 17300 64872
rect 17342 64758 17368 64872
rect 17274 64390 17368 64758
rect 17274 64272 17300 64390
rect 17342 64272 17368 64390
rect 17968 64754 17994 64872
rect 18036 64754 18062 64872
rect 17968 64386 18062 64754
rect 17968 64272 17994 64386
rect 18036 64272 18062 64386
rect 18662 64734 18714 64872
rect 19332 64734 19358 64916
rect 18662 64598 19358 64734
rect 18662 64272 18714 64598
rect 19332 64316 19358 64598
rect 19958 64780 19984 64916
rect 20026 64780 20052 64916
rect 19958 64408 20052 64780
rect 19958 64316 19984 64408
rect 20026 64316 20052 64408
rect 20652 64316 20758 64916
rect 3394 63982 3420 64204
rect 2740 63838 3420 63982
rect 2740 63608 2792 63838
rect 2762 63550 2792 63608
rect 3394 63604 3420 63838
rect 4020 64086 4046 64204
rect 4088 64086 4114 64204
rect 4020 63718 4114 64086
rect 4020 63604 4046 63718
rect 4088 63604 4114 63718
rect 4714 64132 4740 64204
rect 4782 64132 4808 64204
rect 4714 63764 4808 64132
rect 4714 63604 4740 63764
rect 4782 63604 4808 63764
rect 5408 64014 5460 64204
rect 6068 64014 6094 64210
rect 5408 63870 6094 64014
rect 5408 63604 5460 63870
rect 6068 63610 6094 63870
rect 6694 64092 6720 64210
rect 6762 64092 6788 64210
rect 6694 63724 6788 64092
rect 6694 63610 6720 63724
rect 6762 63610 6788 63724
rect 7388 64138 7414 64210
rect 7456 64138 7482 64210
rect 7388 63770 7482 64138
rect 7388 63610 7414 63770
rect 7456 63610 7482 63770
rect 8082 63998 8134 64210
rect 8714 63998 8740 64210
rect 8082 63820 8740 63998
rect 8082 63610 8134 63820
rect 8714 63610 8740 63820
rect 9340 64092 9366 64210
rect 9408 64092 9434 64210
rect 9340 63724 9434 64092
rect 9340 63610 9366 63724
rect 9408 63610 9434 63724
rect 10034 64138 10060 64210
rect 10102 64138 10128 64210
rect 10034 63770 10128 64138
rect 10034 63610 10060 63770
rect 10102 63610 10128 63770
rect 10728 64054 10780 64210
rect 13404 64204 13434 64262
rect 16058 64210 16088 64268
rect 18684 64214 18714 64272
rect 20672 64258 20758 64316
rect 11368 64054 11394 64204
rect 10728 63876 11394 64054
rect 10728 63610 10780 63876
rect 726 62950 752 63550
rect 1352 63444 1378 63550
rect 1420 63444 1446 63550
rect 1352 63076 1446 63444
rect 1352 62950 1378 63076
rect 1420 62950 1446 63076
rect 2046 63442 2072 63550
rect 2114 63442 2140 63550
rect 2046 63074 2140 63442
rect 2046 62950 2072 63074
rect 2114 62950 2140 63074
rect 2740 63276 2792 63550
rect 5430 63546 5460 63604
rect 8104 63552 8134 63610
rect 10750 63552 10780 63610
rect 11368 63604 11394 63876
rect 11994 64086 12020 64204
rect 12062 64086 12088 64204
rect 11994 63718 12088 64086
rect 11994 63604 12020 63718
rect 12062 63604 12088 63718
rect 12688 64132 12714 64204
rect 12756 64132 12782 64204
rect 12688 63764 12782 64132
rect 12688 63604 12714 63764
rect 12756 63604 12782 63764
rect 13382 64070 13434 64204
rect 14022 64070 14048 64210
rect 13382 63892 14048 64070
rect 13382 63604 13434 63892
rect 14022 63610 14048 63892
rect 14648 64092 14674 64210
rect 14716 64092 14742 64210
rect 14648 63724 14742 64092
rect 14648 63610 14674 63724
rect 14716 63610 14742 63724
rect 15342 64138 15368 64210
rect 15410 64138 15436 64210
rect 15342 63770 15436 64138
rect 15342 63610 15368 63770
rect 15410 63610 15436 63770
rect 16036 64014 16088 64210
rect 16648 64014 16674 64214
rect 16036 63856 16674 64014
rect 16036 63610 16088 63856
rect 16648 63614 16674 63856
rect 17274 64096 17300 64214
rect 17342 64096 17368 64214
rect 17274 63728 17368 64096
rect 17274 63614 17300 63728
rect 17342 63614 17368 63728
rect 17968 64142 17994 64214
rect 18036 64142 18062 64214
rect 17968 63774 18062 64142
rect 17968 63614 17994 63774
rect 18036 63614 18062 63774
rect 18662 64062 18714 64214
rect 19332 64062 19358 64258
rect 18662 63926 19358 64062
rect 18662 63614 18714 63926
rect 19332 63658 19358 63926
rect 19958 64154 19984 64258
rect 20026 64154 20052 64258
rect 19958 63782 20052 64154
rect 19958 63658 19984 63782
rect 20026 63658 20052 63782
rect 20652 64192 20758 64258
rect 20652 64128 20826 64192
rect 20652 64054 20714 64128
rect 20798 64054 20826 64128
rect 20652 63964 20826 64054
rect 20652 63658 20758 63964
rect 3394 63276 3420 63546
rect 2740 63132 3420 63276
rect 2740 62950 2792 63132
rect 2762 62892 2792 62950
rect 3394 62946 3420 63132
rect 4020 63440 4046 63546
rect 4088 63440 4114 63546
rect 4020 63072 4114 63440
rect 4020 62946 4046 63072
rect 4088 62946 4114 63072
rect 4714 63438 4740 63546
rect 4782 63438 4808 63546
rect 4714 63070 4808 63438
rect 4714 62946 4740 63070
rect 4782 62946 4808 63070
rect 5408 63366 5460 63546
rect 6068 63366 6094 63552
rect 5408 63222 6094 63366
rect 5408 62946 5460 63222
rect 6068 62952 6094 63222
rect 6694 63446 6720 63552
rect 6762 63446 6788 63552
rect 6694 63078 6788 63446
rect 6694 62952 6720 63078
rect 6762 62952 6788 63078
rect 7388 63444 7414 63552
rect 7456 63444 7482 63552
rect 7388 63076 7482 63444
rect 7388 62952 7414 63076
rect 7456 62952 7482 63076
rect 8082 63376 8134 63552
rect 8714 63376 8740 63552
rect 8082 63198 8740 63376
rect 8082 62952 8134 63198
rect 8714 62952 8740 63198
rect 9340 63446 9366 63552
rect 9408 63446 9434 63552
rect 9340 63078 9434 63446
rect 9340 62952 9366 63078
rect 9408 62952 9434 63078
rect 10034 63444 10060 63552
rect 10102 63444 10128 63552
rect 10034 63076 10128 63444
rect 10034 62952 10060 63076
rect 10102 62952 10128 63076
rect 10728 63436 10780 63552
rect 13404 63546 13434 63604
rect 16058 63552 16088 63610
rect 18684 63556 18714 63614
rect 20672 63600 20758 63658
rect 11368 63436 11394 63546
rect 10728 63258 11394 63436
rect 10728 62952 10780 63258
rect 726 62292 752 62892
rect 1352 62752 1378 62892
rect 1420 62752 1446 62892
rect 1352 62384 1446 62752
rect 1352 62292 1378 62384
rect 1420 62292 1446 62384
rect 2046 62774 2072 62892
rect 2114 62774 2140 62892
rect 2046 62406 2140 62774
rect 2046 62292 2072 62406
rect 2114 62292 2140 62406
rect 2740 62698 2792 62892
rect 5430 62888 5460 62946
rect 8104 62894 8134 62952
rect 10750 62894 10780 62952
rect 11368 62946 11394 63258
rect 11994 63440 12020 63546
rect 12062 63440 12088 63546
rect 11994 63072 12088 63440
rect 11994 62946 12020 63072
rect 12062 62946 12088 63072
rect 12688 63438 12714 63546
rect 12756 63438 12782 63546
rect 12688 63070 12782 63438
rect 12688 62946 12714 63070
rect 12756 62946 12782 63070
rect 13382 63444 13434 63546
rect 14022 63444 14048 63552
rect 13382 63266 14048 63444
rect 13382 62946 13434 63266
rect 14022 62952 14048 63266
rect 14648 63446 14674 63552
rect 14716 63446 14742 63552
rect 14648 63078 14742 63446
rect 14648 62952 14674 63078
rect 14716 62952 14742 63078
rect 15342 63444 15368 63552
rect 15410 63444 15436 63552
rect 15342 63076 15436 63444
rect 15342 62952 15368 63076
rect 15410 62952 15436 63076
rect 16036 63346 16088 63552
rect 16648 63346 16674 63556
rect 16036 63188 16674 63346
rect 16036 62952 16088 63188
rect 16648 62956 16674 63188
rect 17274 63450 17300 63556
rect 17342 63450 17368 63556
rect 17274 63082 17368 63450
rect 17274 62956 17300 63082
rect 17342 62956 17368 63082
rect 17968 63448 17994 63556
rect 18036 63448 18062 63556
rect 17968 63080 18062 63448
rect 17968 62956 17994 63080
rect 18036 62956 18062 63080
rect 18662 63380 18714 63556
rect 19332 63380 19358 63600
rect 18662 63244 19358 63380
rect 18662 62956 18714 63244
rect 19332 63000 19358 63244
rect 19958 63456 19984 63600
rect 20026 63456 20052 63600
rect 19958 63084 20052 63456
rect 19958 63000 19984 63084
rect 20026 63000 20052 63084
rect 20652 63000 20758 63600
rect 3394 62698 3420 62888
rect 2740 62554 3420 62698
rect 2740 62292 2792 62554
rect 2762 62234 2792 62292
rect 3394 62288 3420 62554
rect 4020 62748 4046 62888
rect 4088 62748 4114 62888
rect 4020 62380 4114 62748
rect 4020 62288 4046 62380
rect 4088 62288 4114 62380
rect 4714 62770 4740 62888
rect 4782 62770 4808 62888
rect 4714 62402 4808 62770
rect 4714 62288 4740 62402
rect 4782 62288 4808 62402
rect 5408 62740 5460 62888
rect 6068 62740 6094 62894
rect 5408 62596 6094 62740
rect 5408 62288 5460 62596
rect 6068 62294 6094 62596
rect 6694 62754 6720 62894
rect 6762 62754 6788 62894
rect 6694 62386 6788 62754
rect 6694 62294 6720 62386
rect 6762 62294 6788 62386
rect 7388 62776 7414 62894
rect 7456 62776 7482 62894
rect 7388 62408 7482 62776
rect 7388 62294 7414 62408
rect 7456 62294 7482 62408
rect 8082 62844 8134 62894
rect 8714 62844 8740 62894
rect 8082 62666 8740 62844
rect 8082 62294 8134 62666
rect 8714 62294 8740 62666
rect 9340 62754 9366 62894
rect 9408 62754 9434 62894
rect 9340 62386 9434 62754
rect 9340 62294 9366 62386
rect 9408 62294 9434 62386
rect 10034 62776 10060 62894
rect 10102 62776 10128 62894
rect 10034 62408 10128 62776
rect 10034 62294 10060 62408
rect 10102 62294 10128 62408
rect 10728 62738 10780 62894
rect 13404 62888 13434 62946
rect 16058 62894 16088 62952
rect 18684 62898 18714 62956
rect 20672 62942 20758 63000
rect 11368 62738 11394 62888
rect 10728 62560 11394 62738
rect 10728 62294 10780 62560
rect 726 61634 752 62234
rect 1352 62086 1378 62234
rect 1420 62086 1446 62234
rect 1352 61718 1446 62086
rect 1352 61634 1378 61718
rect 1420 61634 1446 61718
rect 2046 62072 2072 62234
rect 2114 62072 2140 62234
rect 2046 61704 2140 62072
rect 2046 61634 2072 61704
rect 2114 61634 2140 61704
rect 2740 62124 2792 62234
rect 5430 62230 5460 62288
rect 8104 62236 8134 62294
rect 10750 62236 10780 62294
rect 11368 62288 11394 62560
rect 11994 62748 12020 62888
rect 12062 62748 12088 62888
rect 11994 62380 12088 62748
rect 11994 62288 12020 62380
rect 12062 62288 12088 62380
rect 12688 62770 12714 62888
rect 12756 62770 12782 62888
rect 12688 62402 12782 62770
rect 12688 62288 12714 62402
rect 12756 62288 12782 62402
rect 13382 62708 13434 62888
rect 14022 62708 14048 62894
rect 13382 62530 14048 62708
rect 13382 62288 13434 62530
rect 14022 62294 14048 62530
rect 14648 62754 14674 62894
rect 14716 62754 14742 62894
rect 14648 62386 14742 62754
rect 14648 62294 14674 62386
rect 14716 62294 14742 62386
rect 15342 62776 15368 62894
rect 15410 62776 15436 62894
rect 15342 62408 15436 62776
rect 15342 62294 15368 62408
rect 15410 62294 15436 62408
rect 16036 62686 16088 62894
rect 16648 62686 16674 62898
rect 16036 62528 16674 62686
rect 16036 62294 16088 62528
rect 16648 62298 16674 62528
rect 17274 62758 17300 62898
rect 17342 62758 17368 62898
rect 17274 62390 17368 62758
rect 17274 62298 17300 62390
rect 17342 62298 17368 62390
rect 17968 62780 17994 62898
rect 18036 62780 18062 62898
rect 17968 62412 18062 62780
rect 17968 62298 17994 62412
rect 18036 62298 18062 62412
rect 18662 62758 18714 62898
rect 19332 62758 19358 62942
rect 18662 62622 19358 62758
rect 18662 62298 18714 62622
rect 19332 62342 19358 62622
rect 19958 62826 19984 62942
rect 20026 62826 20052 62942
rect 19958 62454 20052 62826
rect 19958 62342 19984 62454
rect 20026 62342 20052 62454
rect 20652 62342 20758 62942
rect 3394 62124 3420 62230
rect 2740 61980 3420 62124
rect 2740 61634 2792 61980
rect 2762 61576 2792 61634
rect 3394 61630 3420 61980
rect 4020 62082 4046 62230
rect 4088 62082 4114 62230
rect 4020 61714 4114 62082
rect 4020 61630 4046 61714
rect 4088 61630 4114 61714
rect 4714 62068 4740 62230
rect 4782 62068 4808 62230
rect 4714 61700 4808 62068
rect 4714 61630 4740 61700
rect 4782 61630 4808 61700
rect 5408 62036 5460 62230
rect 6068 62036 6094 62236
rect 5408 61892 6094 62036
rect 5408 61630 5460 61892
rect 6068 61636 6094 61892
rect 6694 62088 6720 62236
rect 6762 62088 6788 62236
rect 6694 61720 6788 62088
rect 6694 61636 6720 61720
rect 6762 61636 6788 61720
rect 7388 62074 7414 62236
rect 7456 62074 7482 62236
rect 7388 61706 7482 62074
rect 7388 61636 7414 61706
rect 7456 61636 7482 61706
rect 8082 62102 8134 62236
rect 8714 62102 8740 62236
rect 8082 61924 8740 62102
rect 8082 61636 8134 61924
rect 8714 61636 8740 61924
rect 9340 62088 9366 62236
rect 9408 62088 9434 62236
rect 9340 61720 9434 62088
rect 9340 61636 9366 61720
rect 9408 61636 9434 61720
rect 10034 62074 10060 62236
rect 10102 62074 10128 62236
rect 10034 61706 10128 62074
rect 10034 61636 10060 61706
rect 10102 61636 10128 61706
rect 10728 62108 10780 62236
rect 13404 62230 13434 62288
rect 16058 62236 16088 62294
rect 18684 62240 18714 62298
rect 20672 62284 20758 62342
rect 11368 62108 11394 62230
rect 10728 61930 11394 62108
rect 10728 61636 10780 61930
rect 726 60976 752 61576
rect 1352 61414 1378 61576
rect 1420 61414 1446 61576
rect 1352 61046 1446 61414
rect 1352 60976 1378 61046
rect 1420 60976 1446 61046
rect 2046 61418 2072 61576
rect 2114 61418 2140 61576
rect 2046 61050 2140 61418
rect 2046 60976 2072 61050
rect 2114 60976 2140 61050
rect 2740 61500 2792 61576
rect 5430 61572 5460 61630
rect 8104 61578 8134 61636
rect 10750 61578 10780 61636
rect 11368 61630 11394 61930
rect 11994 62082 12020 62230
rect 12062 62082 12088 62230
rect 11994 61714 12088 62082
rect 11994 61630 12020 61714
rect 12062 61630 12088 61714
rect 12688 62068 12714 62230
rect 12756 62068 12782 62230
rect 12688 61700 12782 62068
rect 12688 61630 12714 61700
rect 12756 61630 12782 61700
rect 13382 62098 13434 62230
rect 14022 62098 14048 62236
rect 13382 61920 14048 62098
rect 13382 61630 13434 61920
rect 14022 61636 14048 61920
rect 14648 62088 14674 62236
rect 14716 62088 14742 62236
rect 14648 61720 14742 62088
rect 14648 61636 14674 61720
rect 14716 61636 14742 61720
rect 15342 62074 15368 62236
rect 15410 62074 15436 62236
rect 15342 61706 15436 62074
rect 15342 61636 15368 61706
rect 15410 61636 15436 61706
rect 16036 62022 16088 62236
rect 16648 62022 16674 62240
rect 16036 61864 16674 62022
rect 16036 61636 16088 61864
rect 16648 61640 16674 61864
rect 17274 62092 17300 62240
rect 17342 62092 17368 62240
rect 17274 61724 17368 62092
rect 17274 61640 17300 61724
rect 17342 61640 17368 61724
rect 17968 62078 17994 62240
rect 18036 62078 18062 62240
rect 17968 61710 18062 62078
rect 17968 61640 17994 61710
rect 18036 61640 18062 61710
rect 18662 62052 18714 62240
rect 19332 62052 19358 62284
rect 18662 61916 19358 62052
rect 18662 61640 18714 61916
rect 19332 61684 19358 61916
rect 19958 62162 19984 62284
rect 20026 62162 20052 62284
rect 19958 61790 20052 62162
rect 19958 61684 19984 61790
rect 20026 61684 20052 61790
rect 20652 61684 20758 62284
rect 3394 61500 3420 61572
rect 2740 61356 3420 61500
rect 2740 60976 2792 61356
rect 2762 60918 2792 60976
rect 3394 60972 3420 61356
rect 4020 61410 4046 61572
rect 4088 61410 4114 61572
rect 4020 61042 4114 61410
rect 4020 60972 4046 61042
rect 4088 60972 4114 61042
rect 4714 61414 4740 61572
rect 4782 61414 4808 61572
rect 4714 61046 4808 61414
rect 4714 60972 4740 61046
rect 4782 60972 4808 61046
rect 5408 61472 5460 61572
rect 6068 61472 6094 61578
rect 5408 61328 6094 61472
rect 5408 60972 5460 61328
rect 6068 60978 6094 61328
rect 6694 61416 6720 61578
rect 6762 61416 6788 61578
rect 6694 61048 6788 61416
rect 6694 60978 6720 61048
rect 6762 60978 6788 61048
rect 7388 61420 7414 61578
rect 7456 61420 7482 61578
rect 7388 61052 7482 61420
rect 7388 60978 7414 61052
rect 7456 60978 7482 61052
rect 8082 61472 8134 61578
rect 8714 61472 8740 61578
rect 8082 61294 8740 61472
rect 8082 60978 8134 61294
rect 8714 60978 8740 61294
rect 9340 61416 9366 61578
rect 9408 61416 9434 61578
rect 9340 61048 9434 61416
rect 9340 60978 9366 61048
rect 9408 60978 9434 61048
rect 10034 61420 10060 61578
rect 10102 61420 10128 61578
rect 10034 61052 10128 61420
rect 10034 60978 10060 61052
rect 10102 60978 10128 61052
rect 10728 61460 10780 61578
rect 13404 61572 13434 61630
rect 16058 61578 16088 61636
rect 18684 61582 18714 61640
rect 20672 61626 20758 61684
rect 11368 61460 11394 61572
rect 10728 61282 11394 61460
rect 10728 60978 10780 61282
rect 726 60318 752 60918
rect 1352 60790 1378 60918
rect 1420 60790 1446 60918
rect 1352 60436 1446 60790
rect 1352 60318 1378 60436
rect 1420 60318 1446 60436
rect 2046 60778 2072 60918
rect 2114 60778 2140 60918
rect 2046 60424 2140 60778
rect 2046 60318 2072 60424
rect 2114 60318 2140 60424
rect 2740 60614 2792 60918
rect 5430 60914 5460 60972
rect 8104 60920 8134 60978
rect 10750 60920 10780 60978
rect 11368 60972 11394 61282
rect 11994 61410 12020 61572
rect 12062 61410 12088 61572
rect 11994 61042 12088 61410
rect 11994 60972 12020 61042
rect 12062 60972 12088 61042
rect 12688 61414 12714 61572
rect 12756 61414 12782 61572
rect 12688 61046 12782 61414
rect 12688 60972 12714 61046
rect 12756 60972 12782 61046
rect 13382 61430 13434 61572
rect 14022 61430 14048 61578
rect 13382 61252 14048 61430
rect 13382 60972 13434 61252
rect 14022 60978 14048 61252
rect 14648 61416 14674 61578
rect 14716 61416 14742 61578
rect 14648 61048 14742 61416
rect 14648 60978 14674 61048
rect 14716 60978 14742 61048
rect 15342 61420 15368 61578
rect 15410 61420 15436 61578
rect 15342 61052 15436 61420
rect 15342 60978 15368 61052
rect 15410 60978 15436 61052
rect 16036 61418 16088 61578
rect 16648 61418 16674 61582
rect 16036 61260 16674 61418
rect 16036 60978 16088 61260
rect 16648 60982 16674 61260
rect 17274 61420 17300 61582
rect 17342 61420 17368 61582
rect 17274 61052 17368 61420
rect 17274 60982 17300 61052
rect 17342 60982 17368 61052
rect 17968 61424 17994 61582
rect 18036 61424 18062 61582
rect 17968 61056 18062 61424
rect 17968 60982 17994 61056
rect 18036 60982 18062 61056
rect 18662 61438 18714 61582
rect 19332 61438 19358 61626
rect 18662 61302 19358 61438
rect 18662 60982 18714 61302
rect 19332 61026 19358 61302
rect 19958 61496 19984 61626
rect 20026 61496 20052 61626
rect 19958 61124 20052 61496
rect 19958 61026 19984 61124
rect 20026 61026 20052 61124
rect 20652 61026 20758 61626
rect 3394 60614 3420 60914
rect 2740 60470 3420 60614
rect 2740 60354 2792 60470
rect 2740 60318 2766 60354
rect 3394 60314 3420 60470
rect 4020 60786 4046 60914
rect 4088 60786 4114 60914
rect 4020 60432 4114 60786
rect 4020 60314 4046 60432
rect 4088 60314 4114 60432
rect 4714 60774 4740 60914
rect 4782 60774 4808 60914
rect 4714 60420 4808 60774
rect 4714 60314 4740 60420
rect 4782 60314 4808 60420
rect 5408 60588 5460 60914
rect 6068 60588 6094 60920
rect 5408 60444 6094 60588
rect 5408 60350 5460 60444
rect 5408 60314 5434 60350
rect 6068 60320 6094 60444
rect 6694 60792 6720 60920
rect 6762 60792 6788 60920
rect 6694 60438 6788 60792
rect 6694 60320 6720 60438
rect 6762 60320 6788 60438
rect 7388 60780 7414 60920
rect 7456 60780 7482 60920
rect 7388 60426 7482 60780
rect 7388 60320 7414 60426
rect 7456 60320 7482 60426
rect 8082 60622 8134 60920
rect 8714 60622 8740 60920
rect 8082 60444 8740 60622
rect 8082 60356 8134 60444
rect 8082 60320 8108 60356
rect 8714 60320 8740 60444
rect 9340 60792 9366 60920
rect 9408 60792 9434 60920
rect 9340 60438 9434 60792
rect 9340 60320 9366 60438
rect 9408 60320 9434 60438
rect 10034 60780 10060 60920
rect 10102 60780 10128 60920
rect 10034 60426 10128 60780
rect 10034 60320 10060 60426
rect 10102 60320 10128 60426
rect 10728 60622 10780 60920
rect 13404 60914 13434 60972
rect 16058 60920 16088 60978
rect 18684 60924 18714 60982
rect 20672 60968 20758 61026
rect 11368 60622 11394 60914
rect 10728 60444 11394 60622
rect 10728 60356 10780 60444
rect 10728 60320 10754 60356
rect 11368 60314 11394 60444
rect 11994 60786 12020 60914
rect 12062 60786 12088 60914
rect 11994 60432 12088 60786
rect 11994 60314 12020 60432
rect 12062 60314 12088 60432
rect 12688 60774 12714 60914
rect 12756 60774 12782 60914
rect 12688 60420 12782 60774
rect 12688 60314 12714 60420
rect 12756 60314 12782 60420
rect 13382 60600 13434 60914
rect 14022 60600 14048 60920
rect 13382 60422 14048 60600
rect 13382 60350 13434 60422
rect 13382 60314 13408 60350
rect 14022 60320 14048 60422
rect 14648 60792 14674 60920
rect 14716 60792 14742 60920
rect 14648 60438 14742 60792
rect 14648 60320 14674 60438
rect 14716 60320 14742 60438
rect 15342 60780 15368 60920
rect 15410 60780 15436 60920
rect 15342 60426 15436 60780
rect 15342 60320 15368 60426
rect 15410 60320 15436 60426
rect 16036 60612 16088 60920
rect 16648 60612 16674 60924
rect 16036 60468 16674 60612
rect 16036 60356 16088 60468
rect 16036 60320 16062 60356
rect 16648 60324 16674 60468
rect 17274 60796 17300 60924
rect 17342 60796 17368 60924
rect 17274 60442 17368 60796
rect 17274 60324 17300 60442
rect 17342 60324 17368 60442
rect 17968 60784 17994 60924
rect 18036 60784 18062 60924
rect 17968 60430 18062 60784
rect 17968 60324 17994 60430
rect 18036 60324 18062 60430
rect 18662 60694 18714 60924
rect 19332 60694 19358 60968
rect 18662 60558 19358 60694
rect 18662 60360 18714 60558
rect 19332 60368 19358 60558
rect 19958 60884 19984 60968
rect 20026 60884 20052 60968
rect 19958 60512 20052 60884
rect 19958 60368 19984 60512
rect 20026 60368 20052 60512
rect 20652 60474 20758 60968
rect 20652 60368 20678 60474
rect 18662 60324 18688 60360
rect 698 58656 724 59256
rect 1324 59160 1350 59256
rect 1392 59160 1418 59256
rect 1324 58792 1418 59160
rect 1324 58656 1350 58792
rect 1392 58656 1418 58792
rect 2018 59166 2044 59256
rect 2086 59166 2112 59256
rect 2018 58798 2112 59166
rect 2018 58656 2044 58798
rect 2086 58656 2112 58798
rect 2712 58882 2738 59256
rect 2712 58860 2764 58882
rect 3366 58860 3392 59252
rect 2712 58716 3392 58860
rect 2712 58656 2764 58716
rect 2734 58598 2764 58656
rect 3366 58652 3392 58716
rect 3992 59156 4018 59252
rect 4060 59156 4086 59252
rect 3992 58788 4086 59156
rect 3992 58652 4018 58788
rect 4060 58652 4086 58788
rect 4686 59162 4712 59252
rect 4754 59162 4780 59252
rect 4686 58794 4780 59162
rect 4686 58652 4712 58794
rect 4754 58652 4780 58794
rect 5380 58878 5406 59252
rect 5380 58858 5432 58878
rect 6040 58858 6066 59258
rect 5380 58714 6066 58858
rect 5380 58652 5432 58714
rect 6040 58658 6066 58714
rect 6666 59162 6692 59258
rect 6734 59162 6760 59258
rect 6666 58794 6760 59162
rect 6666 58658 6692 58794
rect 6734 58658 6760 58794
rect 7360 59168 7386 59258
rect 7428 59168 7454 59258
rect 7360 58800 7454 59168
rect 7360 58658 7386 58800
rect 7428 58658 7454 58800
rect 8054 59162 8080 59258
rect 8054 58898 8114 59162
rect 8686 58898 8712 59258
rect 8054 58728 8712 58898
rect 8054 58658 8106 58728
rect 8686 58658 8712 58728
rect 9312 59162 9338 59258
rect 9380 59162 9406 59258
rect 9312 58794 9406 59162
rect 9312 58658 9338 58794
rect 9380 58658 9406 58794
rect 10006 59168 10032 59258
rect 10074 59168 10100 59258
rect 10006 58800 10100 59168
rect 10006 58658 10032 58800
rect 10074 58658 10100 58800
rect 10700 59250 10726 59258
rect 10700 59100 10764 59250
rect 11340 59100 11366 59252
rect 10700 58922 11366 59100
rect 10700 58852 10764 58922
rect 10700 58658 10752 58852
rect 698 57998 724 58598
rect 1324 58484 1350 58598
rect 1392 58484 1418 58598
rect 1324 58116 1418 58484
rect 1324 57998 1350 58116
rect 1392 57998 1418 58116
rect 2018 58480 2044 58598
rect 2086 58480 2112 58598
rect 2018 58112 2112 58480
rect 2018 57998 2044 58112
rect 2086 57998 2112 58112
rect 2712 58460 2764 58598
rect 5402 58594 5432 58652
rect 8076 58600 8106 58658
rect 10722 58600 10752 58658
rect 11340 58652 11366 58922
rect 11966 59156 11992 59252
rect 12034 59156 12060 59252
rect 11966 58788 12060 59156
rect 11966 58652 11992 58788
rect 12034 58652 12060 58788
rect 12660 59162 12686 59252
rect 12728 59162 12754 59252
rect 12660 58794 12754 59162
rect 12660 58652 12686 58794
rect 12728 58652 12754 58794
rect 13354 58880 13380 59252
rect 13994 58880 14020 59258
rect 13354 58702 14020 58880
rect 13354 58652 13406 58702
rect 13994 58658 14020 58702
rect 14620 59162 14646 59258
rect 14688 59162 14714 59258
rect 14620 58794 14714 59162
rect 14620 58658 14646 58794
rect 14688 58658 14714 58794
rect 15314 59168 15340 59258
rect 15382 59168 15408 59258
rect 15314 58800 15408 59168
rect 15314 58658 15340 58800
rect 15382 58658 15408 58800
rect 16008 58884 16034 59258
rect 16008 58880 16060 58884
rect 16620 58880 16646 59262
rect 16008 58722 16646 58880
rect 16008 58658 16060 58722
rect 16620 58662 16646 58722
rect 17246 59166 17272 59262
rect 17314 59166 17340 59262
rect 17246 58798 17340 59166
rect 17246 58662 17272 58798
rect 17314 58662 17340 58798
rect 17940 59172 17966 59262
rect 18008 59172 18034 59262
rect 17940 58804 18034 59172
rect 17940 58662 17966 58804
rect 18008 58662 18034 58804
rect 18634 58892 18660 59262
rect 19304 58892 19330 59306
rect 18634 58756 19330 58892
rect 18634 58662 18686 58756
rect 19304 58706 19330 58756
rect 19930 59194 19956 59306
rect 19998 59194 20024 59306
rect 19930 58822 20024 59194
rect 19930 58706 19956 58822
rect 19998 58706 20024 58822
rect 20624 59080 20650 59306
rect 20624 58706 20726 59080
rect 3366 58460 3392 58594
rect 2712 58316 3392 58460
rect 2712 57998 2764 58316
rect 2734 57940 2764 57998
rect 3366 57994 3392 58316
rect 3992 58480 4018 58594
rect 4060 58480 4086 58594
rect 3992 58112 4086 58480
rect 3992 57994 4018 58112
rect 4060 57994 4086 58112
rect 4686 58476 4712 58594
rect 4754 58476 4780 58594
rect 4686 58108 4780 58476
rect 4686 57994 4712 58108
rect 4754 57994 4780 58108
rect 5380 58364 5432 58594
rect 6040 58364 6066 58600
rect 5380 58220 6066 58364
rect 5380 57994 5432 58220
rect 6040 58000 6066 58220
rect 6666 58486 6692 58600
rect 6734 58486 6760 58600
rect 6666 58118 6760 58486
rect 6666 58000 6692 58118
rect 6734 58000 6760 58118
rect 7360 58482 7386 58600
rect 7428 58482 7454 58600
rect 7360 58114 7454 58482
rect 7360 58000 7386 58114
rect 7428 58000 7454 58114
rect 8054 58398 8106 58600
rect 8686 58398 8712 58600
rect 8054 58228 8712 58398
rect 8054 58000 8106 58228
rect 8686 58000 8712 58228
rect 9312 58486 9338 58600
rect 9380 58486 9406 58600
rect 9312 58118 9406 58486
rect 9312 58000 9338 58118
rect 9380 58000 9406 58118
rect 10006 58482 10032 58600
rect 10074 58482 10100 58600
rect 10006 58114 10100 58482
rect 10006 58000 10032 58114
rect 10074 58000 10100 58114
rect 10700 58444 10752 58600
rect 13376 58594 13406 58652
rect 16030 58600 16060 58658
rect 18656 58604 18686 58662
rect 20640 58648 20726 58706
rect 11340 58444 11366 58594
rect 10700 58266 11366 58444
rect 10700 58000 10752 58266
rect 698 57340 724 57940
rect 1324 57822 1350 57940
rect 1392 57822 1418 57940
rect 1324 57454 1418 57822
rect 1324 57340 1350 57454
rect 1392 57340 1418 57454
rect 2018 57868 2044 57940
rect 2086 57868 2112 57940
rect 2018 57500 2112 57868
rect 2018 57340 2044 57500
rect 2086 57340 2112 57500
rect 2712 57714 2764 57940
rect 5402 57936 5432 57994
rect 8076 57942 8106 58000
rect 10722 57942 10752 58000
rect 11340 57994 11366 58266
rect 11966 58480 11992 58594
rect 12034 58480 12060 58594
rect 11966 58112 12060 58480
rect 11966 57994 11992 58112
rect 12034 57994 12060 58112
rect 12660 58476 12686 58594
rect 12728 58476 12754 58594
rect 12660 58108 12754 58476
rect 12660 57994 12686 58108
rect 12728 57994 12754 58108
rect 13354 58474 13406 58594
rect 13994 58474 14020 58600
rect 13354 58296 14020 58474
rect 13354 57994 13406 58296
rect 13994 58000 14020 58296
rect 14620 58486 14646 58600
rect 14688 58486 14714 58600
rect 14620 58118 14714 58486
rect 14620 58000 14646 58118
rect 14688 58000 14714 58118
rect 15314 58482 15340 58600
rect 15382 58482 15408 58600
rect 15314 58114 15408 58482
rect 15314 58000 15340 58114
rect 15382 58000 15408 58114
rect 16008 58454 16060 58600
rect 16620 58454 16646 58604
rect 16008 58296 16646 58454
rect 16008 58000 16060 58296
rect 16620 58004 16646 58296
rect 17246 58490 17272 58604
rect 17314 58490 17340 58604
rect 17246 58122 17340 58490
rect 17246 58004 17272 58122
rect 17314 58004 17340 58122
rect 17940 58486 17966 58604
rect 18008 58486 18034 58604
rect 17940 58118 18034 58486
rect 17940 58004 17966 58118
rect 18008 58004 18034 58118
rect 18634 58466 18686 58604
rect 19304 58466 19330 58648
rect 18634 58330 19330 58466
rect 18634 58004 18686 58330
rect 19304 58048 19330 58330
rect 19930 58512 19956 58648
rect 19998 58512 20024 58648
rect 19930 58140 20024 58512
rect 19930 58048 19956 58140
rect 19998 58048 20024 58140
rect 20624 58048 20726 58648
rect 3366 57714 3392 57936
rect 2712 57570 3392 57714
rect 2712 57340 2764 57570
rect 2734 57282 2764 57340
rect 3366 57336 3392 57570
rect 3992 57818 4018 57936
rect 4060 57818 4086 57936
rect 3992 57450 4086 57818
rect 3992 57336 4018 57450
rect 4060 57336 4086 57450
rect 4686 57864 4712 57936
rect 4754 57864 4780 57936
rect 4686 57496 4780 57864
rect 4686 57336 4712 57496
rect 4754 57336 4780 57496
rect 5380 57746 5432 57936
rect 6040 57746 6066 57942
rect 5380 57602 6066 57746
rect 5380 57336 5432 57602
rect 6040 57342 6066 57602
rect 6666 57824 6692 57942
rect 6734 57824 6760 57942
rect 6666 57456 6760 57824
rect 6666 57342 6692 57456
rect 6734 57342 6760 57456
rect 7360 57870 7386 57942
rect 7428 57870 7454 57942
rect 7360 57502 7454 57870
rect 7360 57342 7386 57502
rect 7428 57342 7454 57502
rect 8054 57730 8106 57942
rect 8686 57730 8712 57942
rect 8054 57552 8712 57730
rect 8054 57342 8106 57552
rect 8686 57342 8712 57552
rect 9312 57824 9338 57942
rect 9380 57824 9406 57942
rect 9312 57456 9406 57824
rect 9312 57342 9338 57456
rect 9380 57342 9406 57456
rect 10006 57870 10032 57942
rect 10074 57870 10100 57942
rect 10006 57502 10100 57870
rect 10006 57342 10032 57502
rect 10074 57342 10100 57502
rect 10700 57786 10752 57942
rect 13376 57936 13406 57994
rect 16030 57942 16060 58000
rect 18656 57946 18686 58004
rect 20640 57990 20726 58048
rect 11340 57786 11366 57936
rect 10700 57608 11366 57786
rect 10700 57342 10752 57608
rect 698 56682 724 57282
rect 1324 57176 1350 57282
rect 1392 57176 1418 57282
rect 1324 56808 1418 57176
rect 1324 56682 1350 56808
rect 1392 56682 1418 56808
rect 2018 57174 2044 57282
rect 2086 57174 2112 57282
rect 2018 56806 2112 57174
rect 2018 56682 2044 56806
rect 2086 56682 2112 56806
rect 2712 57008 2764 57282
rect 5402 57278 5432 57336
rect 8076 57284 8106 57342
rect 10722 57284 10752 57342
rect 11340 57336 11366 57608
rect 11966 57818 11992 57936
rect 12034 57818 12060 57936
rect 11966 57450 12060 57818
rect 11966 57336 11992 57450
rect 12034 57336 12060 57450
rect 12660 57864 12686 57936
rect 12728 57864 12754 57936
rect 12660 57496 12754 57864
rect 12660 57336 12686 57496
rect 12728 57336 12754 57496
rect 13354 57802 13406 57936
rect 13994 57802 14020 57942
rect 13354 57624 14020 57802
rect 13354 57336 13406 57624
rect 13994 57342 14020 57624
rect 14620 57824 14646 57942
rect 14688 57824 14714 57942
rect 14620 57456 14714 57824
rect 14620 57342 14646 57456
rect 14688 57342 14714 57456
rect 15314 57870 15340 57942
rect 15382 57870 15408 57942
rect 15314 57502 15408 57870
rect 15314 57342 15340 57502
rect 15382 57342 15408 57502
rect 16008 57746 16060 57942
rect 16620 57746 16646 57946
rect 16008 57588 16646 57746
rect 16008 57342 16060 57588
rect 16620 57346 16646 57588
rect 17246 57828 17272 57946
rect 17314 57828 17340 57946
rect 17246 57460 17340 57828
rect 17246 57346 17272 57460
rect 17314 57346 17340 57460
rect 17940 57874 17966 57946
rect 18008 57874 18034 57946
rect 17940 57506 18034 57874
rect 17940 57346 17966 57506
rect 18008 57346 18034 57506
rect 18634 57794 18686 57946
rect 19304 57794 19330 57990
rect 18634 57658 19330 57794
rect 18634 57346 18686 57658
rect 19304 57390 19330 57658
rect 19930 57886 19956 57990
rect 19998 57886 20024 57990
rect 19930 57514 20024 57886
rect 19930 57390 19956 57514
rect 19998 57390 20024 57514
rect 20624 57390 20726 57990
rect 3366 57008 3392 57278
rect 2712 56864 3392 57008
rect 2712 56682 2764 56864
rect 2734 56624 2764 56682
rect 3366 56678 3392 56864
rect 3992 57172 4018 57278
rect 4060 57172 4086 57278
rect 3992 56804 4086 57172
rect 3992 56678 4018 56804
rect 4060 56678 4086 56804
rect 4686 57170 4712 57278
rect 4754 57170 4780 57278
rect 4686 56802 4780 57170
rect 4686 56678 4712 56802
rect 4754 56678 4780 56802
rect 5380 57098 5432 57278
rect 6040 57098 6066 57284
rect 5380 56954 6066 57098
rect 5380 56678 5432 56954
rect 6040 56684 6066 56954
rect 6666 57178 6692 57284
rect 6734 57178 6760 57284
rect 6666 56810 6760 57178
rect 6666 56684 6692 56810
rect 6734 56684 6760 56810
rect 7360 57176 7386 57284
rect 7428 57176 7454 57284
rect 7360 56808 7454 57176
rect 7360 56684 7386 56808
rect 7428 56684 7454 56808
rect 8054 57108 8106 57284
rect 8686 57108 8712 57284
rect 8054 56930 8712 57108
rect 8054 56684 8106 56930
rect 8686 56684 8712 56930
rect 9312 57178 9338 57284
rect 9380 57178 9406 57284
rect 9312 56810 9406 57178
rect 9312 56684 9338 56810
rect 9380 56684 9406 56810
rect 10006 57176 10032 57284
rect 10074 57176 10100 57284
rect 10006 56808 10100 57176
rect 10006 56684 10032 56808
rect 10074 56684 10100 56808
rect 10700 57168 10752 57284
rect 13376 57278 13406 57336
rect 16030 57284 16060 57342
rect 18656 57288 18686 57346
rect 20640 57332 20726 57390
rect 11340 57168 11366 57278
rect 10700 56990 11366 57168
rect 10700 56684 10752 56990
rect 698 56024 724 56624
rect 1324 56484 1350 56624
rect 1392 56484 1418 56624
rect 1324 56116 1418 56484
rect 1324 56024 1350 56116
rect 1392 56024 1418 56116
rect 2018 56506 2044 56624
rect 2086 56506 2112 56624
rect 2018 56138 2112 56506
rect 2018 56024 2044 56138
rect 2086 56024 2112 56138
rect 2712 56430 2764 56624
rect 5402 56620 5432 56678
rect 8076 56626 8106 56684
rect 10722 56626 10752 56684
rect 11340 56678 11366 56990
rect 11966 57172 11992 57278
rect 12034 57172 12060 57278
rect 11966 56804 12060 57172
rect 11966 56678 11992 56804
rect 12034 56678 12060 56804
rect 12660 57170 12686 57278
rect 12728 57170 12754 57278
rect 12660 56802 12754 57170
rect 12660 56678 12686 56802
rect 12728 56678 12754 56802
rect 13354 57176 13406 57278
rect 13994 57176 14020 57284
rect 13354 56998 14020 57176
rect 13354 56678 13406 56998
rect 13994 56684 14020 56998
rect 14620 57178 14646 57284
rect 14688 57178 14714 57284
rect 14620 56810 14714 57178
rect 14620 56684 14646 56810
rect 14688 56684 14714 56810
rect 15314 57176 15340 57284
rect 15382 57176 15408 57284
rect 15314 56808 15408 57176
rect 15314 56684 15340 56808
rect 15382 56684 15408 56808
rect 16008 57078 16060 57284
rect 16620 57078 16646 57288
rect 16008 56920 16646 57078
rect 16008 56684 16060 56920
rect 16620 56688 16646 56920
rect 17246 57182 17272 57288
rect 17314 57182 17340 57288
rect 17246 56814 17340 57182
rect 17246 56688 17272 56814
rect 17314 56688 17340 56814
rect 17940 57180 17966 57288
rect 18008 57180 18034 57288
rect 17940 56812 18034 57180
rect 17940 56688 17966 56812
rect 18008 56688 18034 56812
rect 18634 57112 18686 57288
rect 19304 57112 19330 57332
rect 18634 56976 19330 57112
rect 18634 56688 18686 56976
rect 19304 56732 19330 56976
rect 19930 57188 19956 57332
rect 19998 57188 20024 57332
rect 19930 56816 20024 57188
rect 19930 56732 19956 56816
rect 19998 56732 20024 56816
rect 20624 56732 20726 57332
rect 3366 56430 3392 56620
rect 2712 56286 3392 56430
rect 2712 56024 2764 56286
rect 2734 55966 2764 56024
rect 3366 56020 3392 56286
rect 3992 56480 4018 56620
rect 4060 56480 4086 56620
rect 3992 56112 4086 56480
rect 3992 56020 4018 56112
rect 4060 56020 4086 56112
rect 4686 56502 4712 56620
rect 4754 56502 4780 56620
rect 4686 56134 4780 56502
rect 4686 56020 4712 56134
rect 4754 56020 4780 56134
rect 5380 56472 5432 56620
rect 6040 56472 6066 56626
rect 5380 56328 6066 56472
rect 5380 56020 5432 56328
rect 6040 56026 6066 56328
rect 6666 56486 6692 56626
rect 6734 56486 6760 56626
rect 6666 56118 6760 56486
rect 6666 56026 6692 56118
rect 6734 56026 6760 56118
rect 7360 56508 7386 56626
rect 7428 56508 7454 56626
rect 7360 56140 7454 56508
rect 7360 56026 7386 56140
rect 7428 56026 7454 56140
rect 8054 56576 8106 56626
rect 8686 56576 8712 56626
rect 8054 56398 8712 56576
rect 8054 56026 8106 56398
rect 8686 56026 8712 56398
rect 9312 56486 9338 56626
rect 9380 56486 9406 56626
rect 9312 56118 9406 56486
rect 9312 56026 9338 56118
rect 9380 56026 9406 56118
rect 10006 56508 10032 56626
rect 10074 56508 10100 56626
rect 10006 56140 10100 56508
rect 10006 56026 10032 56140
rect 10074 56026 10100 56140
rect 10700 56470 10752 56626
rect 13376 56620 13406 56678
rect 16030 56626 16060 56684
rect 18656 56630 18686 56688
rect 20640 56674 20726 56732
rect 11340 56470 11366 56620
rect 10700 56292 11366 56470
rect 10700 56026 10752 56292
rect 698 55366 724 55966
rect 1324 55818 1350 55966
rect 1392 55818 1418 55966
rect 1324 55450 1418 55818
rect 1324 55366 1350 55450
rect 1392 55366 1418 55450
rect 2018 55804 2044 55966
rect 2086 55804 2112 55966
rect 2018 55436 2112 55804
rect 2018 55366 2044 55436
rect 2086 55366 2112 55436
rect 2712 55856 2764 55966
rect 5402 55962 5432 56020
rect 8076 55968 8106 56026
rect 10722 55968 10752 56026
rect 11340 56020 11366 56292
rect 11966 56480 11992 56620
rect 12034 56480 12060 56620
rect 11966 56112 12060 56480
rect 11966 56020 11992 56112
rect 12034 56020 12060 56112
rect 12660 56502 12686 56620
rect 12728 56502 12754 56620
rect 12660 56134 12754 56502
rect 12660 56020 12686 56134
rect 12728 56020 12754 56134
rect 13354 56440 13406 56620
rect 13994 56440 14020 56626
rect 13354 56262 14020 56440
rect 13354 56020 13406 56262
rect 13994 56026 14020 56262
rect 14620 56486 14646 56626
rect 14688 56486 14714 56626
rect 14620 56118 14714 56486
rect 14620 56026 14646 56118
rect 14688 56026 14714 56118
rect 15314 56508 15340 56626
rect 15382 56508 15408 56626
rect 15314 56140 15408 56508
rect 15314 56026 15340 56140
rect 15382 56026 15408 56140
rect 16008 56418 16060 56626
rect 16620 56418 16646 56630
rect 16008 56260 16646 56418
rect 16008 56026 16060 56260
rect 16620 56030 16646 56260
rect 17246 56490 17272 56630
rect 17314 56490 17340 56630
rect 17246 56122 17340 56490
rect 17246 56030 17272 56122
rect 17314 56030 17340 56122
rect 17940 56512 17966 56630
rect 18008 56512 18034 56630
rect 17940 56144 18034 56512
rect 17940 56030 17966 56144
rect 18008 56030 18034 56144
rect 18634 56490 18686 56630
rect 19304 56490 19330 56674
rect 18634 56354 19330 56490
rect 18634 56030 18686 56354
rect 19304 56074 19330 56354
rect 19930 56558 19956 56674
rect 19998 56558 20024 56674
rect 19930 56186 20024 56558
rect 19930 56074 19956 56186
rect 19998 56074 20024 56186
rect 20624 56074 20726 56674
rect 3366 55856 3392 55962
rect 2712 55712 3392 55856
rect 2712 55366 2764 55712
rect 2734 55308 2764 55366
rect 3366 55362 3392 55712
rect 3992 55814 4018 55962
rect 4060 55814 4086 55962
rect 3992 55446 4086 55814
rect 3992 55362 4018 55446
rect 4060 55362 4086 55446
rect 4686 55800 4712 55962
rect 4754 55800 4780 55962
rect 4686 55432 4780 55800
rect 4686 55362 4712 55432
rect 4754 55362 4780 55432
rect 5380 55768 5432 55962
rect 6040 55768 6066 55968
rect 5380 55624 6066 55768
rect 5380 55362 5432 55624
rect 6040 55368 6066 55624
rect 6666 55820 6692 55968
rect 6734 55820 6760 55968
rect 6666 55452 6760 55820
rect 6666 55368 6692 55452
rect 6734 55368 6760 55452
rect 7360 55806 7386 55968
rect 7428 55806 7454 55968
rect 7360 55438 7454 55806
rect 7360 55368 7386 55438
rect 7428 55368 7454 55438
rect 8054 55834 8106 55968
rect 8686 55834 8712 55968
rect 8054 55656 8712 55834
rect 8054 55368 8106 55656
rect 8686 55368 8712 55656
rect 9312 55820 9338 55968
rect 9380 55820 9406 55968
rect 9312 55452 9406 55820
rect 9312 55368 9338 55452
rect 9380 55368 9406 55452
rect 10006 55806 10032 55968
rect 10074 55806 10100 55968
rect 10006 55438 10100 55806
rect 10006 55368 10032 55438
rect 10074 55368 10100 55438
rect 10700 55840 10752 55968
rect 13376 55962 13406 56020
rect 16030 55968 16060 56026
rect 18656 55972 18686 56030
rect 20640 56016 20726 56074
rect 11340 55840 11366 55962
rect 10700 55662 11366 55840
rect 10700 55368 10752 55662
rect 698 54708 724 55308
rect 1324 55146 1350 55308
rect 1392 55146 1418 55308
rect 1324 54778 1418 55146
rect 1324 54708 1350 54778
rect 1392 54708 1418 54778
rect 2018 55150 2044 55308
rect 2086 55150 2112 55308
rect 2018 54782 2112 55150
rect 2018 54708 2044 54782
rect 2086 54708 2112 54782
rect 2712 55232 2764 55308
rect 5402 55304 5432 55362
rect 8076 55310 8106 55368
rect 10722 55310 10752 55368
rect 11340 55362 11366 55662
rect 11966 55814 11992 55962
rect 12034 55814 12060 55962
rect 11966 55446 12060 55814
rect 11966 55362 11992 55446
rect 12034 55362 12060 55446
rect 12660 55800 12686 55962
rect 12728 55800 12754 55962
rect 12660 55432 12754 55800
rect 12660 55362 12686 55432
rect 12728 55362 12754 55432
rect 13354 55830 13406 55962
rect 13994 55830 14020 55968
rect 13354 55652 14020 55830
rect 13354 55362 13406 55652
rect 13994 55368 14020 55652
rect 14620 55820 14646 55968
rect 14688 55820 14714 55968
rect 14620 55452 14714 55820
rect 14620 55368 14646 55452
rect 14688 55368 14714 55452
rect 15314 55806 15340 55968
rect 15382 55806 15408 55968
rect 15314 55438 15408 55806
rect 15314 55368 15340 55438
rect 15382 55368 15408 55438
rect 16008 55754 16060 55968
rect 16620 55754 16646 55972
rect 16008 55596 16646 55754
rect 16008 55368 16060 55596
rect 16620 55372 16646 55596
rect 17246 55824 17272 55972
rect 17314 55824 17340 55972
rect 17246 55456 17340 55824
rect 17246 55372 17272 55456
rect 17314 55372 17340 55456
rect 17940 55810 17966 55972
rect 18008 55810 18034 55972
rect 17940 55442 18034 55810
rect 17940 55372 17966 55442
rect 18008 55372 18034 55442
rect 18634 55784 18686 55972
rect 19304 55784 19330 56016
rect 18634 55648 19330 55784
rect 18634 55372 18686 55648
rect 19304 55416 19330 55648
rect 19930 55894 19956 56016
rect 19998 55894 20024 56016
rect 19930 55522 20024 55894
rect 19930 55416 19956 55522
rect 19998 55416 20024 55522
rect 20624 55416 20726 56016
rect 3366 55232 3392 55304
rect 2712 55088 3392 55232
rect 2712 54708 2764 55088
rect 2734 54650 2764 54708
rect 3366 54704 3392 55088
rect 3992 55142 4018 55304
rect 4060 55142 4086 55304
rect 3992 54774 4086 55142
rect 3992 54704 4018 54774
rect 4060 54704 4086 54774
rect 4686 55146 4712 55304
rect 4754 55146 4780 55304
rect 4686 54778 4780 55146
rect 4686 54704 4712 54778
rect 4754 54704 4780 54778
rect 5380 55204 5432 55304
rect 6040 55204 6066 55310
rect 5380 55060 6066 55204
rect 5380 54704 5432 55060
rect 6040 54710 6066 55060
rect 6666 55148 6692 55310
rect 6734 55148 6760 55310
rect 6666 54780 6760 55148
rect 6666 54710 6692 54780
rect 6734 54710 6760 54780
rect 7360 55152 7386 55310
rect 7428 55152 7454 55310
rect 7360 54784 7454 55152
rect 7360 54710 7386 54784
rect 7428 54710 7454 54784
rect 8054 55204 8106 55310
rect 8686 55204 8712 55310
rect 8054 55026 8712 55204
rect 8054 54710 8106 55026
rect 8686 54710 8712 55026
rect 9312 55148 9338 55310
rect 9380 55148 9406 55310
rect 9312 54780 9406 55148
rect 9312 54710 9338 54780
rect 9380 54710 9406 54780
rect 10006 55152 10032 55310
rect 10074 55152 10100 55310
rect 10006 54784 10100 55152
rect 10006 54710 10032 54784
rect 10074 54710 10100 54784
rect 10700 55192 10752 55310
rect 13376 55304 13406 55362
rect 16030 55310 16060 55368
rect 18656 55314 18686 55372
rect 20640 55358 20726 55416
rect 11340 55192 11366 55304
rect 10700 55014 11366 55192
rect 10700 54710 10752 55014
rect 698 54050 724 54650
rect 1324 54522 1350 54650
rect 1392 54522 1418 54650
rect 1324 54168 1418 54522
rect 1324 54050 1350 54168
rect 1392 54050 1418 54168
rect 2018 54510 2044 54650
rect 2086 54510 2112 54650
rect 2018 54156 2112 54510
rect 2018 54050 2044 54156
rect 2086 54050 2112 54156
rect 2712 54346 2764 54650
rect 5402 54646 5432 54704
rect 8076 54652 8106 54710
rect 10722 54652 10752 54710
rect 11340 54704 11366 55014
rect 11966 55142 11992 55304
rect 12034 55142 12060 55304
rect 11966 54774 12060 55142
rect 11966 54704 11992 54774
rect 12034 54704 12060 54774
rect 12660 55146 12686 55304
rect 12728 55146 12754 55304
rect 12660 54778 12754 55146
rect 12660 54704 12686 54778
rect 12728 54704 12754 54778
rect 13354 55162 13406 55304
rect 13994 55162 14020 55310
rect 13354 54984 14020 55162
rect 13354 54704 13406 54984
rect 13994 54710 14020 54984
rect 14620 55148 14646 55310
rect 14688 55148 14714 55310
rect 14620 54780 14714 55148
rect 14620 54710 14646 54780
rect 14688 54710 14714 54780
rect 15314 55152 15340 55310
rect 15382 55152 15408 55310
rect 15314 54784 15408 55152
rect 15314 54710 15340 54784
rect 15382 54710 15408 54784
rect 16008 55150 16060 55310
rect 16620 55150 16646 55314
rect 16008 54992 16646 55150
rect 16008 54710 16060 54992
rect 16620 54714 16646 54992
rect 17246 55152 17272 55314
rect 17314 55152 17340 55314
rect 17246 54784 17340 55152
rect 17246 54714 17272 54784
rect 17314 54714 17340 54784
rect 17940 55156 17966 55314
rect 18008 55156 18034 55314
rect 17940 54788 18034 55156
rect 17940 54714 17966 54788
rect 18008 54714 18034 54788
rect 18634 55170 18686 55314
rect 19304 55170 19330 55358
rect 18634 55034 19330 55170
rect 18634 54714 18686 55034
rect 19304 54758 19330 55034
rect 19930 55228 19956 55358
rect 19998 55228 20024 55358
rect 19930 54856 20024 55228
rect 19930 54758 19956 54856
rect 19998 54758 20024 54856
rect 20624 54758 20726 55358
rect 3366 54346 3392 54646
rect 2712 54202 3392 54346
rect 2712 54086 2764 54202
rect 2712 54050 2738 54086
rect 3366 54046 3392 54202
rect 3992 54518 4018 54646
rect 4060 54518 4086 54646
rect 3992 54164 4086 54518
rect 3992 54046 4018 54164
rect 4060 54046 4086 54164
rect 4686 54506 4712 54646
rect 4754 54506 4780 54646
rect 4686 54152 4780 54506
rect 4686 54046 4712 54152
rect 4754 54046 4780 54152
rect 5380 54320 5432 54646
rect 6040 54320 6066 54652
rect 5380 54176 6066 54320
rect 5380 54082 5432 54176
rect 5380 54046 5406 54082
rect 6040 54052 6066 54176
rect 6666 54524 6692 54652
rect 6734 54524 6760 54652
rect 6666 54170 6760 54524
rect 6666 54052 6692 54170
rect 6734 54052 6760 54170
rect 7360 54512 7386 54652
rect 7428 54512 7454 54652
rect 7360 54158 7454 54512
rect 7360 54052 7386 54158
rect 7428 54052 7454 54158
rect 8054 54354 8106 54652
rect 8686 54354 8712 54652
rect 8054 54176 8712 54354
rect 8054 54088 8106 54176
rect 8054 54052 8080 54088
rect 8686 54052 8712 54176
rect 9312 54524 9338 54652
rect 9380 54524 9406 54652
rect 9312 54170 9406 54524
rect 9312 54052 9338 54170
rect 9380 54052 9406 54170
rect 10006 54512 10032 54652
rect 10074 54512 10100 54652
rect 10006 54158 10100 54512
rect 10006 54052 10032 54158
rect 10074 54052 10100 54158
rect 10700 54354 10752 54652
rect 13376 54646 13406 54704
rect 16030 54652 16060 54710
rect 18656 54656 18686 54714
rect 20640 54740 20726 54758
rect 20640 54700 20840 54740
rect 11340 54354 11366 54646
rect 10700 54176 11366 54354
rect 10700 54088 10752 54176
rect 10700 54052 10726 54088
rect 11340 54046 11366 54176
rect 11966 54518 11992 54646
rect 12034 54518 12060 54646
rect 11966 54164 12060 54518
rect 11966 54046 11992 54164
rect 12034 54046 12060 54164
rect 12660 54506 12686 54646
rect 12728 54506 12754 54646
rect 12660 54152 12754 54506
rect 12660 54046 12686 54152
rect 12728 54046 12754 54152
rect 13354 54332 13406 54646
rect 13994 54332 14020 54652
rect 13354 54154 14020 54332
rect 13354 54082 13406 54154
rect 13354 54046 13380 54082
rect 13994 54052 14020 54154
rect 14620 54524 14646 54652
rect 14688 54524 14714 54652
rect 14620 54170 14714 54524
rect 14620 54052 14646 54170
rect 14688 54052 14714 54170
rect 15314 54512 15340 54652
rect 15382 54512 15408 54652
rect 15314 54158 15408 54512
rect 15314 54052 15340 54158
rect 15382 54052 15408 54158
rect 16008 54344 16060 54652
rect 16620 54344 16646 54656
rect 16008 54200 16646 54344
rect 16008 54088 16060 54200
rect 16008 54052 16034 54088
rect 16620 54056 16646 54200
rect 17246 54528 17272 54656
rect 17314 54528 17340 54656
rect 17246 54174 17340 54528
rect 17246 54056 17272 54174
rect 17314 54056 17340 54174
rect 17940 54516 17966 54656
rect 18008 54516 18034 54656
rect 17940 54162 18034 54516
rect 17940 54056 17966 54162
rect 18008 54056 18034 54162
rect 18634 54426 18686 54656
rect 19304 54426 19330 54700
rect 18634 54290 19330 54426
rect 18634 54092 18686 54290
rect 19304 54100 19330 54290
rect 19930 54616 19956 54700
rect 19998 54616 20024 54700
rect 19930 54244 20024 54616
rect 19930 54100 19956 54244
rect 19998 54100 20024 54244
rect 20624 54660 20840 54700
rect 20624 54424 20678 54660
rect 20792 54424 20840 54660
rect 20624 54364 20840 54424
rect 20624 54362 20726 54364
rect 20624 54100 20650 54362
rect 18634 54056 18660 54092
rect 698 52290 724 52890
rect 1324 52794 1350 52890
rect 1392 52794 1418 52890
rect 1324 52426 1418 52794
rect 1324 52290 1350 52426
rect 1392 52290 1418 52426
rect 2018 52800 2044 52890
rect 2086 52800 2112 52890
rect 2018 52432 2112 52800
rect 2018 52290 2044 52432
rect 2086 52290 2112 52432
rect 2712 52516 2738 52890
rect 2712 52494 2764 52516
rect 3366 52494 3392 52886
rect 2712 52350 3392 52494
rect 2712 52290 2764 52350
rect 2734 52232 2764 52290
rect 3366 52286 3392 52350
rect 3992 52790 4018 52886
rect 4060 52790 4086 52886
rect 3992 52422 4086 52790
rect 3992 52286 4018 52422
rect 4060 52286 4086 52422
rect 4686 52796 4712 52886
rect 4754 52796 4780 52886
rect 4686 52428 4780 52796
rect 4686 52286 4712 52428
rect 4754 52286 4780 52428
rect 5380 52512 5406 52886
rect 5380 52492 5432 52512
rect 6040 52492 6066 52892
rect 5380 52348 6066 52492
rect 5380 52286 5432 52348
rect 6040 52292 6066 52348
rect 6666 52796 6692 52892
rect 6734 52796 6760 52892
rect 6666 52428 6760 52796
rect 6666 52292 6692 52428
rect 6734 52292 6760 52428
rect 7360 52802 7386 52892
rect 7428 52802 7454 52892
rect 7360 52434 7454 52802
rect 7360 52292 7386 52434
rect 7428 52292 7454 52434
rect 8054 52796 8080 52892
rect 8054 52532 8114 52796
rect 8686 52532 8712 52892
rect 8054 52362 8712 52532
rect 8054 52292 8106 52362
rect 8686 52292 8712 52362
rect 9312 52796 9338 52892
rect 9380 52796 9406 52892
rect 9312 52428 9406 52796
rect 9312 52292 9338 52428
rect 9380 52292 9406 52428
rect 10006 52802 10032 52892
rect 10074 52802 10100 52892
rect 10006 52434 10100 52802
rect 10006 52292 10032 52434
rect 10074 52292 10100 52434
rect 10700 52884 10726 52892
rect 10700 52734 10764 52884
rect 11340 52734 11366 52886
rect 10700 52556 11366 52734
rect 10700 52486 10764 52556
rect 10700 52292 10752 52486
rect 698 51632 724 52232
rect 1324 52118 1350 52232
rect 1392 52118 1418 52232
rect 1324 51750 1418 52118
rect 1324 51632 1350 51750
rect 1392 51632 1418 51750
rect 2018 52114 2044 52232
rect 2086 52114 2112 52232
rect 2018 51746 2112 52114
rect 2018 51632 2044 51746
rect 2086 51632 2112 51746
rect 2712 52094 2764 52232
rect 5402 52228 5432 52286
rect 8076 52234 8106 52292
rect 10722 52234 10752 52292
rect 11340 52286 11366 52556
rect 11966 52790 11992 52886
rect 12034 52790 12060 52886
rect 11966 52422 12060 52790
rect 11966 52286 11992 52422
rect 12034 52286 12060 52422
rect 12660 52796 12686 52886
rect 12728 52796 12754 52886
rect 12660 52428 12754 52796
rect 12660 52286 12686 52428
rect 12728 52286 12754 52428
rect 13354 52514 13380 52886
rect 13994 52514 14020 52892
rect 13354 52336 14020 52514
rect 13354 52286 13406 52336
rect 13994 52292 14020 52336
rect 14620 52796 14646 52892
rect 14688 52796 14714 52892
rect 14620 52428 14714 52796
rect 14620 52292 14646 52428
rect 14688 52292 14714 52428
rect 15314 52802 15340 52892
rect 15382 52802 15408 52892
rect 15314 52434 15408 52802
rect 15314 52292 15340 52434
rect 15382 52292 15408 52434
rect 16008 52518 16034 52892
rect 16008 52514 16060 52518
rect 16620 52514 16646 52896
rect 16008 52356 16646 52514
rect 16008 52292 16060 52356
rect 16620 52296 16646 52356
rect 17246 52800 17272 52896
rect 17314 52800 17340 52896
rect 17246 52432 17340 52800
rect 17246 52296 17272 52432
rect 17314 52296 17340 52432
rect 17940 52806 17966 52896
rect 18008 52806 18034 52896
rect 17940 52438 18034 52806
rect 17940 52296 17966 52438
rect 18008 52296 18034 52438
rect 18634 52526 18660 52896
rect 19304 52526 19330 52940
rect 18634 52390 19330 52526
rect 18634 52296 18686 52390
rect 19304 52340 19330 52390
rect 19930 52828 19956 52940
rect 19998 52828 20024 52940
rect 19930 52456 20024 52828
rect 19930 52340 19956 52456
rect 19998 52340 20024 52456
rect 20624 52696 20650 52940
rect 20624 52340 20712 52696
rect 3366 52094 3392 52228
rect 2712 51950 3392 52094
rect 2712 51632 2764 51950
rect 2734 51574 2764 51632
rect 3366 51628 3392 51950
rect 3992 52114 4018 52228
rect 4060 52114 4086 52228
rect 3992 51746 4086 52114
rect 3992 51628 4018 51746
rect 4060 51628 4086 51746
rect 4686 52110 4712 52228
rect 4754 52110 4780 52228
rect 4686 51742 4780 52110
rect 4686 51628 4712 51742
rect 4754 51628 4780 51742
rect 5380 51998 5432 52228
rect 6040 51998 6066 52234
rect 5380 51854 6066 51998
rect 5380 51628 5432 51854
rect 6040 51634 6066 51854
rect 6666 52120 6692 52234
rect 6734 52120 6760 52234
rect 6666 51752 6760 52120
rect 6666 51634 6692 51752
rect 6734 51634 6760 51752
rect 7360 52116 7386 52234
rect 7428 52116 7454 52234
rect 7360 51748 7454 52116
rect 7360 51634 7386 51748
rect 7428 51634 7454 51748
rect 8054 52032 8106 52234
rect 8686 52032 8712 52234
rect 8054 51862 8712 52032
rect 8054 51634 8106 51862
rect 8686 51634 8712 51862
rect 9312 52120 9338 52234
rect 9380 52120 9406 52234
rect 9312 51752 9406 52120
rect 9312 51634 9338 51752
rect 9380 51634 9406 51752
rect 10006 52116 10032 52234
rect 10074 52116 10100 52234
rect 10006 51748 10100 52116
rect 10006 51634 10032 51748
rect 10074 51634 10100 51748
rect 10700 52078 10752 52234
rect 13376 52228 13406 52286
rect 16030 52234 16060 52292
rect 18656 52238 18686 52296
rect 20644 52282 20712 52340
rect 11340 52078 11366 52228
rect 10700 51900 11366 52078
rect 10700 51634 10752 51900
rect 698 50974 724 51574
rect 1324 51456 1350 51574
rect 1392 51456 1418 51574
rect 1324 51088 1418 51456
rect 1324 50974 1350 51088
rect 1392 50974 1418 51088
rect 2018 51502 2044 51574
rect 2086 51502 2112 51574
rect 2018 51134 2112 51502
rect 2018 50974 2044 51134
rect 2086 50974 2112 51134
rect 2712 51348 2764 51574
rect 5402 51570 5432 51628
rect 8076 51576 8106 51634
rect 10722 51576 10752 51634
rect 11340 51628 11366 51900
rect 11966 52114 11992 52228
rect 12034 52114 12060 52228
rect 11966 51746 12060 52114
rect 11966 51628 11992 51746
rect 12034 51628 12060 51746
rect 12660 52110 12686 52228
rect 12728 52110 12754 52228
rect 12660 51742 12754 52110
rect 12660 51628 12686 51742
rect 12728 51628 12754 51742
rect 13354 52108 13406 52228
rect 13994 52108 14020 52234
rect 13354 51930 14020 52108
rect 13354 51628 13406 51930
rect 13994 51634 14020 51930
rect 14620 52120 14646 52234
rect 14688 52120 14714 52234
rect 14620 51752 14714 52120
rect 14620 51634 14646 51752
rect 14688 51634 14714 51752
rect 15314 52116 15340 52234
rect 15382 52116 15408 52234
rect 15314 51748 15408 52116
rect 15314 51634 15340 51748
rect 15382 51634 15408 51748
rect 16008 52088 16060 52234
rect 16620 52088 16646 52238
rect 16008 51930 16646 52088
rect 16008 51634 16060 51930
rect 16620 51638 16646 51930
rect 17246 52124 17272 52238
rect 17314 52124 17340 52238
rect 17246 51756 17340 52124
rect 17246 51638 17272 51756
rect 17314 51638 17340 51756
rect 17940 52120 17966 52238
rect 18008 52120 18034 52238
rect 17940 51752 18034 52120
rect 17940 51638 17966 51752
rect 18008 51638 18034 51752
rect 18634 52100 18686 52238
rect 19304 52100 19330 52282
rect 18634 51964 19330 52100
rect 18634 51638 18686 51964
rect 19304 51682 19330 51964
rect 19930 52146 19956 52282
rect 19998 52146 20024 52282
rect 19930 51774 20024 52146
rect 19930 51682 19956 51774
rect 19998 51682 20024 51774
rect 20624 51682 20712 52282
rect 3366 51348 3392 51570
rect 2712 51204 3392 51348
rect 2712 50974 2764 51204
rect 2734 50916 2764 50974
rect 3366 50970 3392 51204
rect 3992 51452 4018 51570
rect 4060 51452 4086 51570
rect 3992 51084 4086 51452
rect 3992 50970 4018 51084
rect 4060 50970 4086 51084
rect 4686 51498 4712 51570
rect 4754 51498 4780 51570
rect 4686 51130 4780 51498
rect 4686 50970 4712 51130
rect 4754 50970 4780 51130
rect 5380 51380 5432 51570
rect 6040 51380 6066 51576
rect 5380 51236 6066 51380
rect 5380 50970 5432 51236
rect 6040 50976 6066 51236
rect 6666 51458 6692 51576
rect 6734 51458 6760 51576
rect 6666 51090 6760 51458
rect 6666 50976 6692 51090
rect 6734 50976 6760 51090
rect 7360 51504 7386 51576
rect 7428 51504 7454 51576
rect 7360 51136 7454 51504
rect 7360 50976 7386 51136
rect 7428 50976 7454 51136
rect 8054 51364 8106 51576
rect 8686 51364 8712 51576
rect 8054 51186 8712 51364
rect 8054 50976 8106 51186
rect 8686 50976 8712 51186
rect 9312 51458 9338 51576
rect 9380 51458 9406 51576
rect 9312 51090 9406 51458
rect 9312 50976 9338 51090
rect 9380 50976 9406 51090
rect 10006 51504 10032 51576
rect 10074 51504 10100 51576
rect 10006 51136 10100 51504
rect 10006 50976 10032 51136
rect 10074 50976 10100 51136
rect 10700 51420 10752 51576
rect 13376 51570 13406 51628
rect 16030 51576 16060 51634
rect 18656 51580 18686 51638
rect 20644 51624 20712 51682
rect 11340 51420 11366 51570
rect 10700 51242 11366 51420
rect 10700 50976 10752 51242
rect 698 50316 724 50916
rect 1324 50810 1350 50916
rect 1392 50810 1418 50916
rect 1324 50442 1418 50810
rect 1324 50316 1350 50442
rect 1392 50316 1418 50442
rect 2018 50808 2044 50916
rect 2086 50808 2112 50916
rect 2018 50440 2112 50808
rect 2018 50316 2044 50440
rect 2086 50316 2112 50440
rect 2712 50642 2764 50916
rect 5402 50912 5432 50970
rect 8076 50918 8106 50976
rect 10722 50918 10752 50976
rect 11340 50970 11366 51242
rect 11966 51452 11992 51570
rect 12034 51452 12060 51570
rect 11966 51084 12060 51452
rect 11966 50970 11992 51084
rect 12034 50970 12060 51084
rect 12660 51498 12686 51570
rect 12728 51498 12754 51570
rect 12660 51130 12754 51498
rect 12660 50970 12686 51130
rect 12728 50970 12754 51130
rect 13354 51436 13406 51570
rect 13994 51436 14020 51576
rect 13354 51258 14020 51436
rect 13354 50970 13406 51258
rect 13994 50976 14020 51258
rect 14620 51458 14646 51576
rect 14688 51458 14714 51576
rect 14620 51090 14714 51458
rect 14620 50976 14646 51090
rect 14688 50976 14714 51090
rect 15314 51504 15340 51576
rect 15382 51504 15408 51576
rect 15314 51136 15408 51504
rect 15314 50976 15340 51136
rect 15382 50976 15408 51136
rect 16008 51380 16060 51576
rect 16620 51380 16646 51580
rect 16008 51222 16646 51380
rect 16008 50976 16060 51222
rect 16620 50980 16646 51222
rect 17246 51462 17272 51580
rect 17314 51462 17340 51580
rect 17246 51094 17340 51462
rect 17246 50980 17272 51094
rect 17314 50980 17340 51094
rect 17940 51508 17966 51580
rect 18008 51508 18034 51580
rect 17940 51140 18034 51508
rect 17940 50980 17966 51140
rect 18008 50980 18034 51140
rect 18634 51428 18686 51580
rect 19304 51428 19330 51624
rect 18634 51292 19330 51428
rect 18634 50980 18686 51292
rect 19304 51024 19330 51292
rect 19930 51520 19956 51624
rect 19998 51520 20024 51624
rect 19930 51148 20024 51520
rect 19930 51024 19956 51148
rect 19998 51024 20024 51148
rect 20624 51024 20712 51624
rect 3366 50642 3392 50912
rect 2712 50498 3392 50642
rect 2712 50316 2764 50498
rect 2734 50258 2764 50316
rect 3366 50312 3392 50498
rect 3992 50806 4018 50912
rect 4060 50806 4086 50912
rect 3992 50438 4086 50806
rect 3992 50312 4018 50438
rect 4060 50312 4086 50438
rect 4686 50804 4712 50912
rect 4754 50804 4780 50912
rect 4686 50436 4780 50804
rect 4686 50312 4712 50436
rect 4754 50312 4780 50436
rect 5380 50732 5432 50912
rect 6040 50732 6066 50918
rect 5380 50588 6066 50732
rect 5380 50312 5432 50588
rect 6040 50318 6066 50588
rect 6666 50812 6692 50918
rect 6734 50812 6760 50918
rect 6666 50444 6760 50812
rect 6666 50318 6692 50444
rect 6734 50318 6760 50444
rect 7360 50810 7386 50918
rect 7428 50810 7454 50918
rect 7360 50442 7454 50810
rect 7360 50318 7386 50442
rect 7428 50318 7454 50442
rect 8054 50742 8106 50918
rect 8686 50742 8712 50918
rect 8054 50564 8712 50742
rect 8054 50318 8106 50564
rect 8686 50318 8712 50564
rect 9312 50812 9338 50918
rect 9380 50812 9406 50918
rect 9312 50444 9406 50812
rect 9312 50318 9338 50444
rect 9380 50318 9406 50444
rect 10006 50810 10032 50918
rect 10074 50810 10100 50918
rect 10006 50442 10100 50810
rect 10006 50318 10032 50442
rect 10074 50318 10100 50442
rect 10700 50802 10752 50918
rect 13376 50912 13406 50970
rect 16030 50918 16060 50976
rect 18656 50922 18686 50980
rect 20644 50966 20712 51024
rect 11340 50802 11366 50912
rect 10700 50624 11366 50802
rect 10700 50318 10752 50624
rect 698 49658 724 50258
rect 1324 50118 1350 50258
rect 1392 50118 1418 50258
rect 1324 49750 1418 50118
rect 1324 49658 1350 49750
rect 1392 49658 1418 49750
rect 2018 50140 2044 50258
rect 2086 50140 2112 50258
rect 2018 49772 2112 50140
rect 2018 49658 2044 49772
rect 2086 49658 2112 49772
rect 2712 50064 2764 50258
rect 5402 50254 5432 50312
rect 8076 50260 8106 50318
rect 10722 50260 10752 50318
rect 11340 50312 11366 50624
rect 11966 50806 11992 50912
rect 12034 50806 12060 50912
rect 11966 50438 12060 50806
rect 11966 50312 11992 50438
rect 12034 50312 12060 50438
rect 12660 50804 12686 50912
rect 12728 50804 12754 50912
rect 12660 50436 12754 50804
rect 12660 50312 12686 50436
rect 12728 50312 12754 50436
rect 13354 50810 13406 50912
rect 13994 50810 14020 50918
rect 13354 50632 14020 50810
rect 13354 50312 13406 50632
rect 13994 50318 14020 50632
rect 14620 50812 14646 50918
rect 14688 50812 14714 50918
rect 14620 50444 14714 50812
rect 14620 50318 14646 50444
rect 14688 50318 14714 50444
rect 15314 50810 15340 50918
rect 15382 50810 15408 50918
rect 15314 50442 15408 50810
rect 15314 50318 15340 50442
rect 15382 50318 15408 50442
rect 16008 50712 16060 50918
rect 16620 50712 16646 50922
rect 16008 50554 16646 50712
rect 16008 50318 16060 50554
rect 16620 50322 16646 50554
rect 17246 50816 17272 50922
rect 17314 50816 17340 50922
rect 17246 50448 17340 50816
rect 17246 50322 17272 50448
rect 17314 50322 17340 50448
rect 17940 50814 17966 50922
rect 18008 50814 18034 50922
rect 17940 50446 18034 50814
rect 17940 50322 17966 50446
rect 18008 50322 18034 50446
rect 18634 50746 18686 50922
rect 19304 50746 19330 50966
rect 18634 50610 19330 50746
rect 18634 50322 18686 50610
rect 19304 50366 19330 50610
rect 19930 50822 19956 50966
rect 19998 50822 20024 50966
rect 19930 50450 20024 50822
rect 19930 50366 19956 50450
rect 19998 50366 20024 50450
rect 20624 50366 20712 50966
rect 3366 50064 3392 50254
rect 2712 49920 3392 50064
rect 2712 49658 2764 49920
rect 2734 49600 2764 49658
rect 3366 49654 3392 49920
rect 3992 50114 4018 50254
rect 4060 50114 4086 50254
rect 3992 49746 4086 50114
rect 3992 49654 4018 49746
rect 4060 49654 4086 49746
rect 4686 50136 4712 50254
rect 4754 50136 4780 50254
rect 4686 49768 4780 50136
rect 4686 49654 4712 49768
rect 4754 49654 4780 49768
rect 5380 50106 5432 50254
rect 6040 50106 6066 50260
rect 5380 49962 6066 50106
rect 5380 49654 5432 49962
rect 6040 49660 6066 49962
rect 6666 50120 6692 50260
rect 6734 50120 6760 50260
rect 6666 49752 6760 50120
rect 6666 49660 6692 49752
rect 6734 49660 6760 49752
rect 7360 50142 7386 50260
rect 7428 50142 7454 50260
rect 7360 49774 7454 50142
rect 7360 49660 7386 49774
rect 7428 49660 7454 49774
rect 8054 50210 8106 50260
rect 8686 50210 8712 50260
rect 8054 50032 8712 50210
rect 8054 49660 8106 50032
rect 8686 49660 8712 50032
rect 9312 50120 9338 50260
rect 9380 50120 9406 50260
rect 9312 49752 9406 50120
rect 9312 49660 9338 49752
rect 9380 49660 9406 49752
rect 10006 50142 10032 50260
rect 10074 50142 10100 50260
rect 10006 49774 10100 50142
rect 10006 49660 10032 49774
rect 10074 49660 10100 49774
rect 10700 50104 10752 50260
rect 13376 50254 13406 50312
rect 16030 50260 16060 50318
rect 18656 50264 18686 50322
rect 20644 50308 20712 50366
rect 11340 50104 11366 50254
rect 10700 49926 11366 50104
rect 10700 49660 10752 49926
rect 698 49000 724 49600
rect 1324 49452 1350 49600
rect 1392 49452 1418 49600
rect 1324 49084 1418 49452
rect 1324 49000 1350 49084
rect 1392 49000 1418 49084
rect 2018 49438 2044 49600
rect 2086 49438 2112 49600
rect 2018 49070 2112 49438
rect 2018 49000 2044 49070
rect 2086 49000 2112 49070
rect 2712 49490 2764 49600
rect 5402 49596 5432 49654
rect 8076 49602 8106 49660
rect 10722 49602 10752 49660
rect 11340 49654 11366 49926
rect 11966 50114 11992 50254
rect 12034 50114 12060 50254
rect 11966 49746 12060 50114
rect 11966 49654 11992 49746
rect 12034 49654 12060 49746
rect 12660 50136 12686 50254
rect 12728 50136 12754 50254
rect 12660 49768 12754 50136
rect 12660 49654 12686 49768
rect 12728 49654 12754 49768
rect 13354 50074 13406 50254
rect 13994 50074 14020 50260
rect 13354 49896 14020 50074
rect 13354 49654 13406 49896
rect 13994 49660 14020 49896
rect 14620 50120 14646 50260
rect 14688 50120 14714 50260
rect 14620 49752 14714 50120
rect 14620 49660 14646 49752
rect 14688 49660 14714 49752
rect 15314 50142 15340 50260
rect 15382 50142 15408 50260
rect 15314 49774 15408 50142
rect 15314 49660 15340 49774
rect 15382 49660 15408 49774
rect 16008 50052 16060 50260
rect 16620 50052 16646 50264
rect 16008 49894 16646 50052
rect 16008 49660 16060 49894
rect 16620 49664 16646 49894
rect 17246 50124 17272 50264
rect 17314 50124 17340 50264
rect 17246 49756 17340 50124
rect 17246 49664 17272 49756
rect 17314 49664 17340 49756
rect 17940 50146 17966 50264
rect 18008 50146 18034 50264
rect 17940 49778 18034 50146
rect 17940 49664 17966 49778
rect 18008 49664 18034 49778
rect 18634 50124 18686 50264
rect 19304 50124 19330 50308
rect 18634 49988 19330 50124
rect 18634 49664 18686 49988
rect 19304 49708 19330 49988
rect 19930 50192 19956 50308
rect 19998 50192 20024 50308
rect 19930 49820 20024 50192
rect 19930 49708 19956 49820
rect 19998 49708 20024 49820
rect 20624 49708 20712 50308
rect 3366 49490 3392 49596
rect 2712 49346 3392 49490
rect 2712 49000 2764 49346
rect 2734 48942 2764 49000
rect 3366 48996 3392 49346
rect 3992 49448 4018 49596
rect 4060 49448 4086 49596
rect 3992 49080 4086 49448
rect 3992 48996 4018 49080
rect 4060 48996 4086 49080
rect 4686 49434 4712 49596
rect 4754 49434 4780 49596
rect 4686 49066 4780 49434
rect 4686 48996 4712 49066
rect 4754 48996 4780 49066
rect 5380 49402 5432 49596
rect 6040 49402 6066 49602
rect 5380 49258 6066 49402
rect 5380 48996 5432 49258
rect 6040 49002 6066 49258
rect 6666 49454 6692 49602
rect 6734 49454 6760 49602
rect 6666 49086 6760 49454
rect 6666 49002 6692 49086
rect 6734 49002 6760 49086
rect 7360 49440 7386 49602
rect 7428 49440 7454 49602
rect 7360 49072 7454 49440
rect 7360 49002 7386 49072
rect 7428 49002 7454 49072
rect 8054 49468 8106 49602
rect 8686 49468 8712 49602
rect 8054 49290 8712 49468
rect 8054 49002 8106 49290
rect 8686 49002 8712 49290
rect 9312 49454 9338 49602
rect 9380 49454 9406 49602
rect 9312 49086 9406 49454
rect 9312 49002 9338 49086
rect 9380 49002 9406 49086
rect 10006 49440 10032 49602
rect 10074 49440 10100 49602
rect 10006 49072 10100 49440
rect 10006 49002 10032 49072
rect 10074 49002 10100 49072
rect 10700 49474 10752 49602
rect 13376 49596 13406 49654
rect 16030 49602 16060 49660
rect 18656 49606 18686 49664
rect 20644 49650 20712 49708
rect 11340 49474 11366 49596
rect 10700 49296 11366 49474
rect 10700 49002 10752 49296
rect 698 48342 724 48942
rect 1324 48780 1350 48942
rect 1392 48780 1418 48942
rect 1324 48412 1418 48780
rect 1324 48342 1350 48412
rect 1392 48342 1418 48412
rect 2018 48784 2044 48942
rect 2086 48784 2112 48942
rect 2018 48416 2112 48784
rect 2018 48342 2044 48416
rect 2086 48342 2112 48416
rect 2712 48866 2764 48942
rect 5402 48938 5432 48996
rect 8076 48944 8106 49002
rect 10722 48944 10752 49002
rect 11340 48996 11366 49296
rect 11966 49448 11992 49596
rect 12034 49448 12060 49596
rect 11966 49080 12060 49448
rect 11966 48996 11992 49080
rect 12034 48996 12060 49080
rect 12660 49434 12686 49596
rect 12728 49434 12754 49596
rect 12660 49066 12754 49434
rect 12660 48996 12686 49066
rect 12728 48996 12754 49066
rect 13354 49464 13406 49596
rect 13994 49464 14020 49602
rect 13354 49286 14020 49464
rect 13354 48996 13406 49286
rect 13994 49002 14020 49286
rect 14620 49454 14646 49602
rect 14688 49454 14714 49602
rect 14620 49086 14714 49454
rect 14620 49002 14646 49086
rect 14688 49002 14714 49086
rect 15314 49440 15340 49602
rect 15382 49440 15408 49602
rect 15314 49072 15408 49440
rect 15314 49002 15340 49072
rect 15382 49002 15408 49072
rect 16008 49388 16060 49602
rect 16620 49388 16646 49606
rect 16008 49230 16646 49388
rect 16008 49002 16060 49230
rect 16620 49006 16646 49230
rect 17246 49458 17272 49606
rect 17314 49458 17340 49606
rect 17246 49090 17340 49458
rect 17246 49006 17272 49090
rect 17314 49006 17340 49090
rect 17940 49444 17966 49606
rect 18008 49444 18034 49606
rect 17940 49076 18034 49444
rect 17940 49006 17966 49076
rect 18008 49006 18034 49076
rect 18634 49418 18686 49606
rect 19304 49418 19330 49650
rect 18634 49282 19330 49418
rect 18634 49006 18686 49282
rect 19304 49050 19330 49282
rect 19930 49528 19956 49650
rect 19998 49528 20024 49650
rect 19930 49156 20024 49528
rect 19930 49050 19956 49156
rect 19998 49050 20024 49156
rect 20624 49050 20712 49650
rect 3366 48866 3392 48938
rect 2712 48722 3392 48866
rect 2712 48342 2764 48722
rect 2734 48284 2764 48342
rect 3366 48338 3392 48722
rect 3992 48776 4018 48938
rect 4060 48776 4086 48938
rect 3992 48408 4086 48776
rect 3992 48338 4018 48408
rect 4060 48338 4086 48408
rect 4686 48780 4712 48938
rect 4754 48780 4780 48938
rect 4686 48412 4780 48780
rect 4686 48338 4712 48412
rect 4754 48338 4780 48412
rect 5380 48838 5432 48938
rect 6040 48838 6066 48944
rect 5380 48694 6066 48838
rect 5380 48338 5432 48694
rect 6040 48344 6066 48694
rect 6666 48782 6692 48944
rect 6734 48782 6760 48944
rect 6666 48414 6760 48782
rect 6666 48344 6692 48414
rect 6734 48344 6760 48414
rect 7360 48786 7386 48944
rect 7428 48786 7454 48944
rect 7360 48418 7454 48786
rect 7360 48344 7386 48418
rect 7428 48344 7454 48418
rect 8054 48838 8106 48944
rect 8686 48838 8712 48944
rect 8054 48660 8712 48838
rect 8054 48344 8106 48660
rect 8686 48344 8712 48660
rect 9312 48782 9338 48944
rect 9380 48782 9406 48944
rect 9312 48414 9406 48782
rect 9312 48344 9338 48414
rect 9380 48344 9406 48414
rect 10006 48786 10032 48944
rect 10074 48786 10100 48944
rect 10006 48418 10100 48786
rect 10006 48344 10032 48418
rect 10074 48344 10100 48418
rect 10700 48826 10752 48944
rect 13376 48938 13406 48996
rect 16030 48944 16060 49002
rect 18656 48948 18686 49006
rect 20644 48992 20712 49050
rect 11340 48826 11366 48938
rect 10700 48648 11366 48826
rect 10700 48344 10752 48648
rect 698 47684 724 48284
rect 1324 48156 1350 48284
rect 1392 48156 1418 48284
rect 1324 47802 1418 48156
rect 1324 47684 1350 47802
rect 1392 47684 1418 47802
rect 2018 48144 2044 48284
rect 2086 48144 2112 48284
rect 2018 47790 2112 48144
rect 2018 47684 2044 47790
rect 2086 47684 2112 47790
rect 2712 47980 2764 48284
rect 5402 48280 5432 48338
rect 8076 48286 8106 48344
rect 10722 48286 10752 48344
rect 11340 48338 11366 48648
rect 11966 48776 11992 48938
rect 12034 48776 12060 48938
rect 11966 48408 12060 48776
rect 11966 48338 11992 48408
rect 12034 48338 12060 48408
rect 12660 48780 12686 48938
rect 12728 48780 12754 48938
rect 12660 48412 12754 48780
rect 12660 48338 12686 48412
rect 12728 48338 12754 48412
rect 13354 48796 13406 48938
rect 13994 48796 14020 48944
rect 13354 48618 14020 48796
rect 13354 48338 13406 48618
rect 13994 48344 14020 48618
rect 14620 48782 14646 48944
rect 14688 48782 14714 48944
rect 14620 48414 14714 48782
rect 14620 48344 14646 48414
rect 14688 48344 14714 48414
rect 15314 48786 15340 48944
rect 15382 48786 15408 48944
rect 15314 48418 15408 48786
rect 15314 48344 15340 48418
rect 15382 48344 15408 48418
rect 16008 48784 16060 48944
rect 16620 48784 16646 48948
rect 16008 48626 16646 48784
rect 16008 48344 16060 48626
rect 16620 48348 16646 48626
rect 17246 48786 17272 48948
rect 17314 48786 17340 48948
rect 17246 48418 17340 48786
rect 17246 48348 17272 48418
rect 17314 48348 17340 48418
rect 17940 48790 17966 48948
rect 18008 48790 18034 48948
rect 17940 48422 18034 48790
rect 17940 48348 17966 48422
rect 18008 48348 18034 48422
rect 18634 48804 18686 48948
rect 19304 48804 19330 48992
rect 18634 48668 19330 48804
rect 18634 48348 18686 48668
rect 19304 48392 19330 48668
rect 19930 48862 19956 48992
rect 19998 48862 20024 48992
rect 19930 48490 20024 48862
rect 19930 48392 19956 48490
rect 19998 48392 20024 48490
rect 20624 48854 20712 48992
rect 20624 48742 20780 48854
rect 20624 48690 20678 48742
rect 20750 48690 20780 48742
rect 20624 48594 20780 48690
rect 20624 48392 20712 48594
rect 3366 47980 3392 48280
rect 2712 47836 3392 47980
rect 2712 47720 2764 47836
rect 2712 47684 2738 47720
rect 3366 47680 3392 47836
rect 3992 48152 4018 48280
rect 4060 48152 4086 48280
rect 3992 47798 4086 48152
rect 3992 47680 4018 47798
rect 4060 47680 4086 47798
rect 4686 48140 4712 48280
rect 4754 48140 4780 48280
rect 4686 47786 4780 48140
rect 4686 47680 4712 47786
rect 4754 47680 4780 47786
rect 5380 47954 5432 48280
rect 6040 47954 6066 48286
rect 5380 47810 6066 47954
rect 5380 47716 5432 47810
rect 5380 47680 5406 47716
rect 6040 47686 6066 47810
rect 6666 48158 6692 48286
rect 6734 48158 6760 48286
rect 6666 47804 6760 48158
rect 6666 47686 6692 47804
rect 6734 47686 6760 47804
rect 7360 48146 7386 48286
rect 7428 48146 7454 48286
rect 7360 47792 7454 48146
rect 7360 47686 7386 47792
rect 7428 47686 7454 47792
rect 8054 47988 8106 48286
rect 8686 47988 8712 48286
rect 8054 47810 8712 47988
rect 8054 47722 8106 47810
rect 8054 47686 8080 47722
rect 8686 47686 8712 47810
rect 9312 48158 9338 48286
rect 9380 48158 9406 48286
rect 9312 47804 9406 48158
rect 9312 47686 9338 47804
rect 9380 47686 9406 47804
rect 10006 48146 10032 48286
rect 10074 48146 10100 48286
rect 10006 47792 10100 48146
rect 10006 47686 10032 47792
rect 10074 47686 10100 47792
rect 10700 47988 10752 48286
rect 13376 48280 13406 48338
rect 16030 48286 16060 48344
rect 18656 48290 18686 48348
rect 20644 48334 20712 48392
rect 11340 47988 11366 48280
rect 10700 47810 11366 47988
rect 10700 47722 10752 47810
rect 10700 47686 10726 47722
rect 11340 47680 11366 47810
rect 11966 48152 11992 48280
rect 12034 48152 12060 48280
rect 11966 47798 12060 48152
rect 11966 47680 11992 47798
rect 12034 47680 12060 47798
rect 12660 48140 12686 48280
rect 12728 48140 12754 48280
rect 12660 47786 12754 48140
rect 12660 47680 12686 47786
rect 12728 47680 12754 47786
rect 13354 47966 13406 48280
rect 13994 47966 14020 48286
rect 13354 47788 14020 47966
rect 13354 47716 13406 47788
rect 13354 47680 13380 47716
rect 13994 47686 14020 47788
rect 14620 48158 14646 48286
rect 14688 48158 14714 48286
rect 14620 47804 14714 48158
rect 14620 47686 14646 47804
rect 14688 47686 14714 47804
rect 15314 48146 15340 48286
rect 15382 48146 15408 48286
rect 15314 47792 15408 48146
rect 15314 47686 15340 47792
rect 15382 47686 15408 47792
rect 16008 47978 16060 48286
rect 16620 47978 16646 48290
rect 16008 47834 16646 47978
rect 16008 47722 16060 47834
rect 16008 47686 16034 47722
rect 16620 47690 16646 47834
rect 17246 48162 17272 48290
rect 17314 48162 17340 48290
rect 17246 47808 17340 48162
rect 17246 47690 17272 47808
rect 17314 47690 17340 47808
rect 17940 48150 17966 48290
rect 18008 48150 18034 48290
rect 17940 47796 18034 48150
rect 17940 47690 17966 47796
rect 18008 47690 18034 47796
rect 18634 48060 18686 48290
rect 19304 48060 19330 48334
rect 18634 47924 19330 48060
rect 18634 47726 18686 47924
rect 19304 47734 19330 47924
rect 19930 48250 19956 48334
rect 19998 48250 20024 48334
rect 19930 47878 20024 48250
rect 19930 47734 19956 47878
rect 19998 47734 20024 47878
rect 20624 47814 20712 48334
rect 20624 47734 20650 47814
rect 18634 47690 18660 47726
rect 75216 68918 75816 68944
rect 75874 68918 76474 68944
rect 76532 68918 77132 68944
rect 77190 68918 77790 68944
rect 75276 68876 75700 68918
rect 76014 68876 76438 68918
rect 76596 68876 77020 68918
rect 77268 68876 77692 68918
rect 75216 68850 75816 68876
rect 75874 68850 76474 68876
rect 76532 68850 77132 68876
rect 77190 68850 77790 68876
rect 75216 68224 75816 68250
rect 75874 68224 76474 68250
rect 76532 68224 77132 68250
rect 77190 68224 77790 68250
rect 75270 68182 75694 68224
rect 75982 68182 76406 68224
rect 76592 68182 77016 68224
rect 77308 68182 77732 68224
rect 75216 68156 75816 68182
rect 75874 68156 76474 68182
rect 76532 68156 77132 68182
rect 77190 68156 77790 68182
rect 75216 67530 75816 67556
rect 75874 67530 76474 67556
rect 76532 67530 77132 67556
rect 77190 67530 77790 67556
rect 75256 67488 75680 67530
rect 76002 67488 76426 67530
rect 76630 67488 77054 67530
rect 77266 67488 77690 67530
rect 75216 67462 75816 67488
rect 75874 67462 76474 67488
rect 76532 67462 77132 67488
rect 77190 67462 77790 67488
rect 75216 66836 75816 66862
rect 75874 66836 76474 66862
rect 76532 66836 77132 66862
rect 77190 66836 77790 66862
rect 75252 66794 75676 66836
rect 76032 66794 76456 66836
rect 76582 66794 77006 66836
rect 77300 66794 77724 66836
rect 75216 66768 75816 66794
rect 75874 66768 76474 66794
rect 76532 66768 77132 66794
rect 77190 66768 77790 66794
rect 71352 66162 71952 66188
rect 72010 66162 72610 66188
rect 72668 66162 73268 66188
rect 73326 66162 73926 66188
rect 79066 68932 79666 68958
rect 79724 68932 80324 68958
rect 80382 68932 80982 68958
rect 81040 68932 81640 68958
rect 79126 68890 79550 68932
rect 79864 68890 80288 68932
rect 80446 68890 80870 68932
rect 81118 68890 81542 68932
rect 79066 68864 79666 68890
rect 79724 68864 80324 68890
rect 80382 68864 80982 68890
rect 81040 68864 81640 68890
rect 79066 68238 79666 68264
rect 79724 68238 80324 68264
rect 80382 68238 80982 68264
rect 81040 68238 81640 68264
rect 79120 68196 79544 68238
rect 79832 68196 80256 68238
rect 80442 68196 80866 68238
rect 81158 68196 81582 68238
rect 79066 68170 79666 68196
rect 79724 68170 80324 68196
rect 80382 68170 80982 68196
rect 81040 68170 81640 68196
rect 79066 67544 79666 67570
rect 79724 67544 80324 67570
rect 80382 67544 80982 67570
rect 81040 67544 81640 67570
rect 79106 67502 79530 67544
rect 79852 67502 80276 67544
rect 80480 67502 80904 67544
rect 81116 67502 81540 67544
rect 79066 67476 79666 67502
rect 79724 67476 80324 67502
rect 80382 67476 80982 67502
rect 81040 67476 81640 67502
rect 79066 66850 79666 66876
rect 79724 66850 80324 66876
rect 80382 66850 80982 66876
rect 81040 66850 81640 66876
rect 79102 66808 79526 66850
rect 79882 66808 80306 66850
rect 80432 66808 80856 66850
rect 81150 66808 81574 66850
rect 79066 66782 79666 66808
rect 79724 66782 80324 66808
rect 80382 66782 80982 66808
rect 81040 66782 81640 66808
rect 71738 65886 71844 66162
rect 72172 65886 72278 66162
rect 72892 65886 72998 66162
rect 73476 65886 73582 66162
rect 75216 66142 75816 66168
rect 75874 66142 76474 66168
rect 76532 66142 77132 66168
rect 77190 66142 77790 66168
rect 79066 66156 79666 66182
rect 79724 66156 80324 66182
rect 80382 66156 80982 66182
rect 81040 66156 81640 66182
rect 71698 65820 73788 65886
rect 75602 65866 75708 66142
rect 76036 65866 76142 66142
rect 76756 65866 76862 66142
rect 77340 65866 77446 66142
rect 79452 65880 79558 66156
rect 79886 65880 79992 66156
rect 80606 65880 80712 66156
rect 81190 65880 81296 66156
rect 71352 65816 73926 65820
rect 71352 65794 71952 65816
rect 72010 65794 72610 65816
rect 72668 65794 73268 65816
rect 73326 65794 73926 65816
rect 75562 65800 77652 65866
rect 79412 65814 81502 65880
rect 79066 65810 81640 65814
rect 75216 65796 77790 65800
rect 42150 64424 42176 64510
rect 41738 64334 42176 64424
rect 41738 64098 41814 64334
rect 42072 64098 42176 64334
rect 41738 64030 42176 64098
rect 42150 63910 42176 64030
rect 42776 64432 42802 64510
rect 42844 64432 42870 64510
rect 42776 63992 42870 64432
rect 42776 63910 42802 63992
rect 42844 63910 42870 63992
rect 43470 64430 43496 64510
rect 43538 64430 43564 64510
rect 43470 63990 43564 64430
rect 43470 63910 43496 63990
rect 43538 63910 43564 63990
rect 44164 64444 44190 64510
rect 44232 64444 44258 64510
rect 44164 64004 44258 64444
rect 44164 63910 44190 64004
rect 44232 63910 44258 64004
rect 44858 64424 44884 64510
rect 44926 64424 44952 64510
rect 44858 63978 44952 64424
rect 44858 63910 44884 63978
rect 44926 63910 44952 63978
rect 45552 64264 45578 64510
rect 45552 64240 45640 64264
rect 46158 64240 46184 64508
rect 45552 64006 46184 64240
rect 45552 63910 45640 64006
rect 45570 63852 45640 63910
rect 46158 63908 46184 64006
rect 46784 64430 46810 64508
rect 46852 64430 46878 64508
rect 46784 63990 46878 64430
rect 46784 63908 46810 63990
rect 46852 63908 46878 63990
rect 47478 64428 47504 64508
rect 47546 64428 47572 64508
rect 47478 63988 47572 64428
rect 47478 63908 47504 63988
rect 47546 63908 47572 63988
rect 48172 64442 48198 64508
rect 48240 64442 48266 64508
rect 48172 64002 48266 64442
rect 48172 63908 48198 64002
rect 48240 63908 48266 64002
rect 48866 64422 48892 64508
rect 48934 64422 48960 64508
rect 48866 63976 48960 64422
rect 48866 63908 48892 63976
rect 48934 63908 48960 63976
rect 49560 64262 49586 64508
rect 49560 64244 49648 64262
rect 50170 64244 50196 64508
rect 49560 64010 50196 64244
rect 49560 63908 49648 64010
rect 50170 63908 50196 64010
rect 50796 64430 50822 64508
rect 50864 64430 50890 64508
rect 50796 63990 50890 64430
rect 50796 63908 50822 63990
rect 50864 63908 50890 63990
rect 51490 64428 51516 64508
rect 51558 64428 51584 64508
rect 51490 63988 51584 64428
rect 51490 63908 51516 63988
rect 51558 63908 51584 63988
rect 52184 64442 52210 64508
rect 52252 64442 52278 64508
rect 52184 64002 52278 64442
rect 52184 63908 52210 64002
rect 52252 63908 52278 64002
rect 52878 64422 52904 64508
rect 52946 64422 52972 64508
rect 52878 63976 52972 64422
rect 52878 63908 52904 63976
rect 52946 63908 52972 63976
rect 53572 64262 53598 64508
rect 53572 64234 53660 64262
rect 54180 64234 54206 64508
rect 53572 64000 54206 64234
rect 53572 63908 53660 64000
rect 54180 63908 54206 64000
rect 54806 64430 54832 64508
rect 54874 64430 54900 64508
rect 54806 63990 54900 64430
rect 54806 63908 54832 63990
rect 54874 63908 54900 63990
rect 55500 64428 55526 64508
rect 55568 64428 55594 64508
rect 55500 63988 55594 64428
rect 55500 63908 55526 63988
rect 55568 63908 55594 63988
rect 56194 64442 56220 64508
rect 56262 64442 56288 64508
rect 56194 64002 56288 64442
rect 56194 63908 56220 64002
rect 56262 63908 56288 64002
rect 56888 64422 56914 64508
rect 56956 64422 56982 64508
rect 56888 63976 56982 64422
rect 56888 63908 56914 63976
rect 56956 63908 56982 63976
rect 57582 64262 57608 64508
rect 57582 63908 57670 64262
rect 42150 63252 42176 63852
rect 42776 63762 42802 63852
rect 42844 63762 42870 63852
rect 42776 63322 42870 63762
rect 42776 63252 42802 63322
rect 42844 63252 42870 63322
rect 43470 63786 43496 63852
rect 43538 63786 43564 63852
rect 43470 63346 43564 63786
rect 43470 63252 43496 63346
rect 43538 63252 43564 63346
rect 44164 63770 44190 63852
rect 44232 63770 44258 63852
rect 44164 63330 44258 63770
rect 44164 63252 44190 63330
rect 44232 63252 44258 63330
rect 44858 63782 44884 63852
rect 44926 63782 44952 63852
rect 44858 63342 44952 63782
rect 44858 63252 44884 63342
rect 44926 63252 44952 63342
rect 45552 63734 45640 63852
rect 49578 63850 49648 63908
rect 53590 63850 53660 63908
rect 57600 63850 57670 63908
rect 46158 63734 46184 63850
rect 45552 63500 46184 63734
rect 45552 63252 45640 63500
rect 45570 63194 45640 63252
rect 46158 63250 46184 63500
rect 46784 63760 46810 63850
rect 46852 63760 46878 63850
rect 46784 63320 46878 63760
rect 46784 63250 46810 63320
rect 46852 63250 46878 63320
rect 47478 63784 47504 63850
rect 47546 63784 47572 63850
rect 47478 63344 47572 63784
rect 47478 63250 47504 63344
rect 47546 63250 47572 63344
rect 48172 63768 48198 63850
rect 48240 63768 48266 63850
rect 48172 63328 48266 63768
rect 48172 63250 48198 63328
rect 48240 63250 48266 63328
rect 48866 63780 48892 63850
rect 48934 63780 48960 63850
rect 48866 63340 48960 63780
rect 48866 63250 48892 63340
rect 48934 63250 48960 63340
rect 49560 63734 49648 63850
rect 50170 63734 50196 63850
rect 49560 63500 50196 63734
rect 49560 63250 49648 63500
rect 50170 63250 50196 63500
rect 50796 63760 50822 63850
rect 50864 63760 50890 63850
rect 50796 63320 50890 63760
rect 50796 63250 50822 63320
rect 50864 63250 50890 63320
rect 51490 63784 51516 63850
rect 51558 63784 51584 63850
rect 51490 63344 51584 63784
rect 51490 63250 51516 63344
rect 51558 63250 51584 63344
rect 52184 63768 52210 63850
rect 52252 63768 52278 63850
rect 52184 63328 52278 63768
rect 52184 63250 52210 63328
rect 52252 63250 52278 63328
rect 52878 63780 52904 63850
rect 52946 63780 52972 63850
rect 52878 63340 52972 63780
rect 52878 63250 52904 63340
rect 52946 63250 52972 63340
rect 53572 63776 53660 63850
rect 54180 63776 54206 63850
rect 53572 63542 54206 63776
rect 53572 63250 53660 63542
rect 54180 63250 54206 63542
rect 54806 63760 54832 63850
rect 54874 63760 54900 63850
rect 54806 63320 54900 63760
rect 54806 63250 54832 63320
rect 54874 63250 54900 63320
rect 55500 63784 55526 63850
rect 55568 63784 55594 63850
rect 55500 63344 55594 63784
rect 55500 63250 55526 63344
rect 55568 63250 55594 63344
rect 56194 63768 56220 63850
rect 56262 63768 56288 63850
rect 56194 63328 56288 63768
rect 56194 63250 56220 63328
rect 56262 63250 56288 63328
rect 56888 63780 56914 63850
rect 56956 63780 56982 63850
rect 56888 63340 56982 63780
rect 56888 63250 56914 63340
rect 56956 63250 56982 63340
rect 57582 63250 57670 63850
rect 42150 62594 42176 63194
rect 42776 63086 42802 63194
rect 42844 63086 42870 63194
rect 42776 62646 42870 63086
rect 42776 62594 42802 62646
rect 42844 62594 42870 62646
rect 43470 63098 43496 63194
rect 43538 63098 43564 63194
rect 43470 62658 43564 63098
rect 43470 62594 43496 62658
rect 43538 62594 43564 62658
rect 44164 63076 44190 63194
rect 44232 63076 44258 63194
rect 44164 62636 44258 63076
rect 44164 62594 44190 62636
rect 44232 62594 44258 62636
rect 44858 63048 44884 63194
rect 44926 63048 44952 63194
rect 44858 62608 44952 63048
rect 44858 62594 44884 62608
rect 44926 62594 44952 62608
rect 45552 63056 45640 63194
rect 49578 63192 49648 63250
rect 53590 63192 53660 63250
rect 57600 63192 57670 63250
rect 46158 63056 46184 63192
rect 45552 62822 46184 63056
rect 45552 62594 45640 62822
rect 45570 62536 45640 62594
rect 46158 62592 46184 62822
rect 46784 63084 46810 63192
rect 46852 63084 46878 63192
rect 46784 62644 46878 63084
rect 46784 62592 46810 62644
rect 46852 62592 46878 62644
rect 47478 63096 47504 63192
rect 47546 63096 47572 63192
rect 47478 62656 47572 63096
rect 47478 62592 47504 62656
rect 47546 62592 47572 62656
rect 48172 63074 48198 63192
rect 48240 63074 48266 63192
rect 48172 62634 48266 63074
rect 48172 62592 48198 62634
rect 48240 62592 48266 62634
rect 48866 63046 48892 63192
rect 48934 63046 48960 63192
rect 48866 62606 48960 63046
rect 48866 62592 48892 62606
rect 48934 62592 48960 62606
rect 49560 63062 49648 63192
rect 50170 63062 50196 63192
rect 49560 62828 50196 63062
rect 49560 62592 49648 62828
rect 50170 62592 50196 62828
rect 50796 63084 50822 63192
rect 50864 63084 50890 63192
rect 50796 62644 50890 63084
rect 50796 62592 50822 62644
rect 50864 62592 50890 62644
rect 51490 63096 51516 63192
rect 51558 63096 51584 63192
rect 51490 62656 51584 63096
rect 51490 62592 51516 62656
rect 51558 62592 51584 62656
rect 52184 63074 52210 63192
rect 52252 63074 52278 63192
rect 52184 62634 52278 63074
rect 52184 62592 52210 62634
rect 52252 62592 52278 62634
rect 52878 63046 52904 63192
rect 52946 63046 52972 63192
rect 52878 62606 52972 63046
rect 52878 62592 52904 62606
rect 52946 62592 52972 62606
rect 53572 63046 53660 63192
rect 54180 63046 54206 63192
rect 53572 62812 54206 63046
rect 53572 62592 53660 62812
rect 54180 62592 54206 62812
rect 54806 63084 54832 63192
rect 54874 63084 54900 63192
rect 54806 62644 54900 63084
rect 54806 62592 54832 62644
rect 54874 62592 54900 62644
rect 55500 63096 55526 63192
rect 55568 63096 55594 63192
rect 55500 62656 55594 63096
rect 55500 62592 55526 62656
rect 55568 62592 55594 62656
rect 56194 63074 56220 63192
rect 56262 63074 56288 63192
rect 56194 62634 56288 63074
rect 56194 62592 56220 62634
rect 56262 62592 56288 62634
rect 56888 63046 56914 63192
rect 56956 63046 56982 63192
rect 56888 62606 56982 63046
rect 56888 62592 56914 62606
rect 56956 62592 56982 62606
rect 57582 62592 57670 63192
rect 42150 61936 42176 62536
rect 42776 62454 42802 62536
rect 42844 62454 42870 62536
rect 42776 62014 42870 62454
rect 42776 61936 42802 62014
rect 42844 61936 42870 62014
rect 43470 62476 43496 62536
rect 43538 62476 43564 62536
rect 43470 62036 43564 62476
rect 43470 61936 43496 62036
rect 43538 61936 43564 62036
rect 44164 62476 44190 62536
rect 44232 62476 44258 62536
rect 44164 62036 44258 62476
rect 44164 61936 44190 62036
rect 44232 61936 44258 62036
rect 44858 62464 44884 62536
rect 44926 62464 44952 62536
rect 44858 62024 44952 62464
rect 44858 61936 44884 62024
rect 44926 61936 44952 62024
rect 45552 62454 45640 62536
rect 49578 62534 49648 62592
rect 53590 62534 53660 62592
rect 57600 62534 57670 62592
rect 46158 62454 46184 62534
rect 45552 62220 46184 62454
rect 45552 61936 45640 62220
rect 45570 61878 45640 61936
rect 46158 61934 46184 62220
rect 46784 62452 46810 62534
rect 46852 62452 46878 62534
rect 46784 62012 46878 62452
rect 46784 61934 46810 62012
rect 46852 61934 46878 62012
rect 47478 62474 47504 62534
rect 47546 62474 47572 62534
rect 47478 62034 47572 62474
rect 47478 61934 47504 62034
rect 47546 61934 47572 62034
rect 48172 62474 48198 62534
rect 48240 62474 48266 62534
rect 48172 62034 48266 62474
rect 48172 61934 48198 62034
rect 48240 61934 48266 62034
rect 48866 62462 48892 62534
rect 48934 62462 48960 62534
rect 48866 62022 48960 62462
rect 48866 61934 48892 62022
rect 48934 61934 48960 62022
rect 49560 62420 49648 62534
rect 50170 62420 50196 62534
rect 49560 62186 50196 62420
rect 49560 61934 49648 62186
rect 50170 61934 50196 62186
rect 50796 62452 50822 62534
rect 50864 62452 50890 62534
rect 50796 62012 50890 62452
rect 50796 61934 50822 62012
rect 50864 61934 50890 62012
rect 51490 62474 51516 62534
rect 51558 62474 51584 62534
rect 51490 62034 51584 62474
rect 51490 61934 51516 62034
rect 51558 61934 51584 62034
rect 52184 62474 52210 62534
rect 52252 62474 52278 62534
rect 52184 62034 52278 62474
rect 52184 61934 52210 62034
rect 52252 61934 52278 62034
rect 52878 62462 52904 62534
rect 52946 62462 52972 62534
rect 52878 62022 52972 62462
rect 52878 61934 52904 62022
rect 52946 61934 52972 62022
rect 53572 62444 53660 62534
rect 54180 62444 54206 62534
rect 53572 62210 54206 62444
rect 53572 61934 53660 62210
rect 54180 61934 54206 62210
rect 54806 62452 54832 62534
rect 54874 62452 54900 62534
rect 54806 62012 54900 62452
rect 54806 61934 54832 62012
rect 54874 61934 54900 62012
rect 55500 62474 55526 62534
rect 55568 62474 55594 62534
rect 55500 62034 55594 62474
rect 55500 61934 55526 62034
rect 55568 61934 55594 62034
rect 56194 62474 56220 62534
rect 56262 62474 56288 62534
rect 56194 62034 56288 62474
rect 56194 61934 56220 62034
rect 56262 61934 56288 62034
rect 56888 62462 56914 62534
rect 56956 62462 56982 62534
rect 56888 62022 56982 62462
rect 56888 61934 56914 62022
rect 56956 61934 56982 62022
rect 57582 61952 57670 62534
rect 75216 65774 75816 65796
rect 75874 65774 76474 65796
rect 76532 65774 77132 65796
rect 77190 65774 77790 65796
rect 79066 65788 79666 65810
rect 79724 65788 80324 65810
rect 80382 65788 80982 65810
rect 81040 65788 81640 65810
rect 71352 65168 71952 65194
rect 72010 65168 72610 65194
rect 72668 65168 73268 65194
rect 73326 65168 73926 65194
rect 71412 65126 71836 65168
rect 72150 65126 72574 65168
rect 72732 65126 73156 65168
rect 73404 65126 73828 65168
rect 71352 65100 71952 65126
rect 72010 65100 72610 65126
rect 72668 65100 73268 65126
rect 73326 65100 73926 65126
rect 71352 64474 71952 64500
rect 72010 64474 72610 64500
rect 72668 64474 73268 64500
rect 73326 64474 73926 64500
rect 71406 64432 71830 64474
rect 72118 64432 72542 64474
rect 72728 64432 73152 64474
rect 73444 64432 73868 64474
rect 71352 64406 71952 64432
rect 72010 64406 72610 64432
rect 72668 64406 73268 64432
rect 73326 64406 73926 64432
rect 71352 63780 71952 63806
rect 72010 63780 72610 63806
rect 72668 63780 73268 63806
rect 73326 63780 73926 63806
rect 71392 63738 71816 63780
rect 72138 63738 72562 63780
rect 72766 63738 73190 63780
rect 73402 63738 73826 63780
rect 71352 63712 71952 63738
rect 72010 63712 72610 63738
rect 72668 63712 73268 63738
rect 73326 63712 73926 63738
rect 71352 63086 71952 63112
rect 72010 63086 72610 63112
rect 72668 63086 73268 63112
rect 73326 63086 73926 63112
rect 71388 63044 71812 63086
rect 72168 63044 72592 63086
rect 72718 63044 73142 63086
rect 73436 63044 73860 63086
rect 71352 63018 71952 63044
rect 72010 63018 72610 63044
rect 72668 63018 73268 63044
rect 73326 63018 73926 63044
rect 57582 61934 57860 61952
rect 42150 61278 42176 61878
rect 42776 61746 42802 61878
rect 42844 61746 42870 61878
rect 42776 61306 42870 61746
rect 42776 61278 42802 61306
rect 42844 61278 42870 61306
rect 43470 61788 43496 61878
rect 43538 61788 43564 61878
rect 43470 61348 43564 61788
rect 43470 61278 43496 61348
rect 43538 61278 43564 61348
rect 44164 61800 44190 61878
rect 44232 61800 44258 61878
rect 44164 61360 44258 61800
rect 44164 61278 44190 61360
rect 44232 61278 44258 61360
rect 44858 61826 44884 61878
rect 44926 61826 44952 61878
rect 44858 61386 44952 61826
rect 44858 61278 44884 61386
rect 44926 61278 44952 61386
rect 45552 61852 45640 61878
rect 49578 61876 49648 61934
rect 53590 61876 53660 61934
rect 57600 61876 57860 61934
rect 46158 61852 46184 61876
rect 45552 61618 46184 61852
rect 45552 61598 45640 61618
rect 45552 61278 45578 61598
rect 46158 61276 46184 61618
rect 46784 61744 46810 61876
rect 46852 61744 46878 61876
rect 46784 61304 46878 61744
rect 46784 61276 46810 61304
rect 46852 61276 46878 61304
rect 47478 61786 47504 61876
rect 47546 61786 47572 61876
rect 47478 61346 47572 61786
rect 47478 61276 47504 61346
rect 47546 61276 47572 61346
rect 48172 61798 48198 61876
rect 48240 61798 48266 61876
rect 48172 61358 48266 61798
rect 48172 61276 48198 61358
rect 48240 61276 48266 61358
rect 48866 61824 48892 61876
rect 48934 61824 48960 61876
rect 48866 61384 48960 61824
rect 48866 61276 48892 61384
rect 48934 61276 48960 61384
rect 49560 61828 49648 61876
rect 50170 61828 50196 61876
rect 49560 61594 50196 61828
rect 49560 61276 49586 61594
rect 50170 61276 50196 61594
rect 50796 61744 50822 61876
rect 50864 61744 50890 61876
rect 50796 61304 50890 61744
rect 50796 61276 50822 61304
rect 50864 61276 50890 61304
rect 51490 61786 51516 61876
rect 51558 61786 51584 61876
rect 51490 61346 51584 61786
rect 51490 61276 51516 61346
rect 51558 61276 51584 61346
rect 52184 61798 52210 61876
rect 52252 61798 52278 61876
rect 52184 61358 52278 61798
rect 52184 61276 52210 61358
rect 52252 61276 52278 61358
rect 52878 61824 52904 61876
rect 52946 61824 52972 61876
rect 52878 61384 52972 61824
rect 52878 61276 52904 61384
rect 52946 61276 52972 61384
rect 53572 61872 53660 61876
rect 54180 61872 54206 61876
rect 53572 61638 54206 61872
rect 53572 61596 53660 61638
rect 53572 61276 53598 61596
rect 54180 61276 54206 61638
rect 54806 61744 54832 61876
rect 54874 61744 54900 61876
rect 54806 61304 54900 61744
rect 54806 61276 54832 61304
rect 54874 61276 54900 61304
rect 55500 61786 55526 61876
rect 55568 61786 55594 61876
rect 55500 61346 55594 61786
rect 55500 61276 55526 61346
rect 55568 61276 55594 61346
rect 56194 61798 56220 61876
rect 56262 61798 56288 61876
rect 56194 61358 56288 61798
rect 56194 61276 56220 61358
rect 56262 61276 56288 61358
rect 56888 61824 56914 61876
rect 56956 61824 56982 61876
rect 56888 61384 56982 61824
rect 56888 61276 56914 61384
rect 56956 61276 56982 61384
rect 57582 61596 57860 61876
rect 57582 61276 57608 61596
rect 57658 61502 57860 61596
rect 75216 65148 75816 65174
rect 75874 65148 76474 65174
rect 76532 65148 77132 65174
rect 77190 65148 77790 65174
rect 75276 65106 75700 65148
rect 76014 65106 76438 65148
rect 76596 65106 77020 65148
rect 77268 65106 77692 65148
rect 75216 65080 75816 65106
rect 75874 65080 76474 65106
rect 76532 65080 77132 65106
rect 77190 65080 77790 65106
rect 75216 64454 75816 64480
rect 75874 64454 76474 64480
rect 76532 64454 77132 64480
rect 77190 64454 77790 64480
rect 75270 64412 75694 64454
rect 75982 64412 76406 64454
rect 76592 64412 77016 64454
rect 77308 64412 77732 64454
rect 75216 64386 75816 64412
rect 75874 64386 76474 64412
rect 76532 64386 77132 64412
rect 77190 64386 77790 64412
rect 75216 63760 75816 63786
rect 75874 63760 76474 63786
rect 76532 63760 77132 63786
rect 77190 63760 77790 63786
rect 75256 63718 75680 63760
rect 76002 63718 76426 63760
rect 76630 63718 77054 63760
rect 77266 63718 77690 63760
rect 75216 63692 75816 63718
rect 75874 63692 76474 63718
rect 76532 63692 77132 63718
rect 77190 63692 77790 63718
rect 75216 63066 75816 63092
rect 75874 63066 76474 63092
rect 76532 63066 77132 63092
rect 77190 63066 77790 63092
rect 75252 63024 75676 63066
rect 76032 63024 76456 63066
rect 76582 63024 77006 63066
rect 77300 63024 77724 63066
rect 75216 62998 75816 63024
rect 75874 62998 76474 63024
rect 76532 62998 77132 63024
rect 77190 62998 77790 63024
rect 71352 62392 71952 62418
rect 72010 62392 72610 62418
rect 72668 62392 73268 62418
rect 73326 62392 73926 62418
rect 79066 65162 79666 65188
rect 79724 65162 80324 65188
rect 80382 65162 80982 65188
rect 81040 65162 81640 65188
rect 79126 65120 79550 65162
rect 79864 65120 80288 65162
rect 80446 65120 80870 65162
rect 81118 65120 81542 65162
rect 79066 65094 79666 65120
rect 79724 65094 80324 65120
rect 80382 65094 80982 65120
rect 81040 65094 81640 65120
rect 79066 64468 79666 64494
rect 79724 64468 80324 64494
rect 80382 64468 80982 64494
rect 81040 64468 81640 64494
rect 79120 64426 79544 64468
rect 79832 64426 80256 64468
rect 80442 64426 80866 64468
rect 81158 64426 81582 64468
rect 79066 64400 79666 64426
rect 79724 64400 80324 64426
rect 80382 64400 80982 64426
rect 81040 64400 81640 64426
rect 79066 63774 79666 63800
rect 79724 63774 80324 63800
rect 80382 63774 80982 63800
rect 81040 63774 81640 63800
rect 79106 63732 79530 63774
rect 79852 63732 80276 63774
rect 80480 63732 80904 63774
rect 81116 63732 81540 63774
rect 79066 63706 79666 63732
rect 79724 63706 80324 63732
rect 80382 63706 80982 63732
rect 81040 63706 81640 63732
rect 79066 63080 79666 63106
rect 79724 63080 80324 63106
rect 80382 63080 80982 63106
rect 81040 63080 81640 63106
rect 79102 63038 79526 63080
rect 79882 63038 80306 63080
rect 80432 63038 80856 63080
rect 81150 63038 81574 63080
rect 79066 63012 79666 63038
rect 79724 63012 80324 63038
rect 80382 63012 80982 63038
rect 81040 63012 81640 63038
rect 71708 62122 71814 62392
rect 72082 62122 72188 62392
rect 72854 62122 72960 62392
rect 73472 62122 73578 62392
rect 75216 62372 75816 62398
rect 75874 62372 76474 62398
rect 76532 62372 77132 62398
rect 77190 62372 77790 62398
rect 79066 62386 79666 62412
rect 79724 62386 80324 62412
rect 80382 62386 80982 62412
rect 81040 62386 81640 62412
rect 71698 62056 73788 62122
rect 75572 62102 75678 62372
rect 75946 62102 76052 62372
rect 76718 62102 76824 62372
rect 77336 62102 77442 62372
rect 79422 62116 79528 62386
rect 79796 62116 79902 62386
rect 80568 62116 80674 62386
rect 81186 62116 81292 62386
rect 71352 62052 73926 62056
rect 71352 62030 71952 62052
rect 72010 62030 72610 62052
rect 72668 62030 73268 62052
rect 73326 62030 73926 62052
rect 75562 62036 77652 62102
rect 79412 62050 81502 62116
rect 79066 62046 81640 62050
rect 75216 62032 77790 62036
rect 57658 61190 58102 61502
rect 57658 60506 57780 61190
rect 57972 60506 58102 61190
rect 42142 59712 42168 60312
rect 42768 60234 42794 60312
rect 42836 60234 42862 60312
rect 42768 59794 42862 60234
rect 42768 59712 42794 59794
rect 42836 59712 42862 59794
rect 43462 60232 43488 60312
rect 43530 60232 43556 60312
rect 43462 59792 43556 60232
rect 43462 59712 43488 59792
rect 43530 59712 43556 59792
rect 44156 60246 44182 60312
rect 44224 60246 44250 60312
rect 44156 59806 44250 60246
rect 44156 59712 44182 59806
rect 44224 59712 44250 59806
rect 44850 60226 44876 60312
rect 44918 60226 44944 60312
rect 44850 59780 44944 60226
rect 44850 59712 44876 59780
rect 44918 59712 44944 59780
rect 45544 60066 45570 60312
rect 45544 60030 45632 60066
rect 46136 60030 46162 60312
rect 45544 59794 46162 60030
rect 45544 59712 45632 59794
rect 46136 59712 46162 59794
rect 46762 60234 46788 60312
rect 46830 60234 46856 60312
rect 46762 59794 46856 60234
rect 46762 59712 46788 59794
rect 46830 59712 46856 59794
rect 47456 60232 47482 60312
rect 47524 60232 47550 60312
rect 47456 59792 47550 60232
rect 47456 59712 47482 59792
rect 47524 59712 47550 59792
rect 48150 60246 48176 60312
rect 48218 60246 48244 60312
rect 48150 59806 48244 60246
rect 48150 59712 48176 59806
rect 48218 59712 48244 59806
rect 48844 60226 48870 60312
rect 48912 60226 48938 60312
rect 48844 59780 48938 60226
rect 48844 59712 48870 59780
rect 48912 59712 48938 59780
rect 49538 60066 49564 60312
rect 49538 60026 49626 60066
rect 50158 60026 50184 60312
rect 49538 59790 50184 60026
rect 49538 59712 49626 59790
rect 50158 59712 50184 59790
rect 50784 60234 50810 60312
rect 50852 60234 50878 60312
rect 50784 59794 50878 60234
rect 50784 59712 50810 59794
rect 50852 59712 50878 59794
rect 51478 60232 51504 60312
rect 51546 60232 51572 60312
rect 51478 59792 51572 60232
rect 51478 59712 51504 59792
rect 51546 59712 51572 59792
rect 52172 60246 52198 60312
rect 52240 60246 52266 60312
rect 52172 59806 52266 60246
rect 52172 59712 52198 59806
rect 52240 59712 52266 59806
rect 52866 60226 52892 60312
rect 52934 60226 52960 60312
rect 52866 59780 52960 60226
rect 52866 59712 52892 59780
rect 52934 59712 52960 59780
rect 53560 60066 53586 60312
rect 53560 60026 53648 60066
rect 54180 60026 54206 60312
rect 53560 59790 54206 60026
rect 53560 59712 53648 59790
rect 54180 59712 54206 59790
rect 54806 60234 54832 60312
rect 54874 60234 54900 60312
rect 54806 59794 54900 60234
rect 54806 59712 54832 59794
rect 54874 59712 54900 59794
rect 55500 60232 55526 60312
rect 55568 60232 55594 60312
rect 55500 59792 55594 60232
rect 55500 59712 55526 59792
rect 55568 59712 55594 59792
rect 56194 60246 56220 60312
rect 56262 60246 56288 60312
rect 56194 59806 56288 60246
rect 56194 59712 56220 59806
rect 56262 59712 56288 59806
rect 56888 60226 56914 60312
rect 56956 60226 56982 60312
rect 56888 59780 56982 60226
rect 56888 59712 56914 59780
rect 56956 59712 56982 59780
rect 57582 60066 57608 60312
rect 57658 60248 58102 60506
rect 57658 60066 57860 60248
rect 57582 59834 57860 60066
rect 57582 59712 57670 59834
rect 45562 59654 45632 59712
rect 49556 59654 49626 59712
rect 53578 59654 53648 59712
rect 57600 59654 57670 59712
rect 42142 59054 42168 59654
rect 42768 59564 42794 59654
rect 42836 59564 42862 59654
rect 42768 59124 42862 59564
rect 42768 59054 42794 59124
rect 42836 59054 42862 59124
rect 43462 59588 43488 59654
rect 43530 59588 43556 59654
rect 43462 59148 43556 59588
rect 43462 59054 43488 59148
rect 43530 59054 43556 59148
rect 44156 59572 44182 59654
rect 44224 59572 44250 59654
rect 44156 59132 44250 59572
rect 44156 59054 44182 59132
rect 44224 59054 44250 59132
rect 44850 59584 44876 59654
rect 44918 59584 44944 59654
rect 44850 59144 44944 59584
rect 44850 59054 44876 59144
rect 44918 59054 44944 59144
rect 45544 59534 45632 59654
rect 46136 59534 46162 59654
rect 45544 59298 46162 59534
rect 45544 59054 45632 59298
rect 46136 59054 46162 59298
rect 46762 59564 46788 59654
rect 46830 59564 46856 59654
rect 46762 59124 46856 59564
rect 46762 59054 46788 59124
rect 46830 59054 46856 59124
rect 47456 59588 47482 59654
rect 47524 59588 47550 59654
rect 47456 59148 47550 59588
rect 47456 59054 47482 59148
rect 47524 59054 47550 59148
rect 48150 59572 48176 59654
rect 48218 59572 48244 59654
rect 48150 59132 48244 59572
rect 48150 59054 48176 59132
rect 48218 59054 48244 59132
rect 48844 59584 48870 59654
rect 48912 59584 48938 59654
rect 48844 59144 48938 59584
rect 48844 59054 48870 59144
rect 48912 59054 48938 59144
rect 49538 59494 49626 59654
rect 50158 59494 50184 59654
rect 49538 59258 50184 59494
rect 49538 59054 49626 59258
rect 50158 59054 50184 59258
rect 50784 59564 50810 59654
rect 50852 59564 50878 59654
rect 50784 59124 50878 59564
rect 50784 59054 50810 59124
rect 50852 59054 50878 59124
rect 51478 59588 51504 59654
rect 51546 59588 51572 59654
rect 51478 59148 51572 59588
rect 51478 59054 51504 59148
rect 51546 59054 51572 59148
rect 52172 59572 52198 59654
rect 52240 59572 52266 59654
rect 52172 59132 52266 59572
rect 52172 59054 52198 59132
rect 52240 59054 52266 59132
rect 52866 59584 52892 59654
rect 52934 59584 52960 59654
rect 52866 59144 52960 59584
rect 52866 59054 52892 59144
rect 52934 59054 52960 59144
rect 53560 59504 53648 59654
rect 54180 59504 54206 59654
rect 53560 59268 54206 59504
rect 53560 59054 53648 59268
rect 54180 59054 54206 59268
rect 54806 59564 54832 59654
rect 54874 59564 54900 59654
rect 54806 59124 54900 59564
rect 54806 59054 54832 59124
rect 54874 59054 54900 59124
rect 55500 59588 55526 59654
rect 55568 59588 55594 59654
rect 55500 59148 55594 59588
rect 55500 59054 55526 59148
rect 55568 59054 55594 59148
rect 56194 59572 56220 59654
rect 56262 59572 56288 59654
rect 56194 59132 56288 59572
rect 56194 59054 56220 59132
rect 56262 59054 56288 59132
rect 56888 59584 56914 59654
rect 56956 59584 56982 59654
rect 56888 59144 56982 59584
rect 56888 59054 56914 59144
rect 56956 59054 56982 59144
rect 57582 59054 57670 59654
rect 45562 58996 45632 59054
rect 49556 58996 49626 59054
rect 53578 58996 53648 59054
rect 57600 58996 57670 59054
rect 42142 58396 42168 58996
rect 42768 58888 42794 58996
rect 42836 58888 42862 58996
rect 42768 58448 42862 58888
rect 42768 58396 42794 58448
rect 42836 58396 42862 58448
rect 43462 58900 43488 58996
rect 43530 58900 43556 58996
rect 43462 58460 43556 58900
rect 43462 58396 43488 58460
rect 43530 58396 43556 58460
rect 44156 58878 44182 58996
rect 44224 58878 44250 58996
rect 44156 58438 44250 58878
rect 44156 58396 44182 58438
rect 44224 58396 44250 58438
rect 44850 58850 44876 58996
rect 44918 58850 44944 58996
rect 44850 58410 44944 58850
rect 44850 58396 44876 58410
rect 44918 58396 44944 58410
rect 45544 58854 45632 58996
rect 46136 58854 46162 58996
rect 45544 58618 46162 58854
rect 45544 58396 45632 58618
rect 46136 58396 46162 58618
rect 46762 58888 46788 58996
rect 46830 58888 46856 58996
rect 46762 58448 46856 58888
rect 46762 58396 46788 58448
rect 46830 58396 46856 58448
rect 47456 58900 47482 58996
rect 47524 58900 47550 58996
rect 47456 58460 47550 58900
rect 47456 58396 47482 58460
rect 47524 58396 47550 58460
rect 48150 58878 48176 58996
rect 48218 58878 48244 58996
rect 48150 58438 48244 58878
rect 48150 58396 48176 58438
rect 48218 58396 48244 58438
rect 48844 58850 48870 58996
rect 48912 58850 48938 58996
rect 48844 58410 48938 58850
rect 48844 58396 48870 58410
rect 48912 58396 48938 58410
rect 49538 58802 49626 58996
rect 50158 58802 50184 58996
rect 49538 58566 50184 58802
rect 49538 58396 49626 58566
rect 50158 58396 50184 58566
rect 50784 58888 50810 58996
rect 50852 58888 50878 58996
rect 50784 58448 50878 58888
rect 50784 58396 50810 58448
rect 50852 58396 50878 58448
rect 51478 58900 51504 58996
rect 51546 58900 51572 58996
rect 51478 58460 51572 58900
rect 51478 58396 51504 58460
rect 51546 58396 51572 58460
rect 52172 58878 52198 58996
rect 52240 58878 52266 58996
rect 52172 58438 52266 58878
rect 52172 58396 52198 58438
rect 52240 58396 52266 58438
rect 52866 58850 52892 58996
rect 52934 58850 52960 58996
rect 52866 58410 52960 58850
rect 52866 58396 52892 58410
rect 52934 58396 52960 58410
rect 53560 58854 53648 58996
rect 54180 58854 54206 58996
rect 53560 58618 54206 58854
rect 53560 58396 53648 58618
rect 54180 58396 54206 58618
rect 54806 58888 54832 58996
rect 54874 58888 54900 58996
rect 54806 58448 54900 58888
rect 54806 58396 54832 58448
rect 54874 58396 54900 58448
rect 55500 58900 55526 58996
rect 55568 58900 55594 58996
rect 55500 58460 55594 58900
rect 55500 58396 55526 58460
rect 55568 58396 55594 58460
rect 56194 58878 56220 58996
rect 56262 58878 56288 58996
rect 56194 58438 56288 58878
rect 56194 58396 56220 58438
rect 56262 58396 56288 58438
rect 56888 58850 56914 58996
rect 56956 58850 56982 58996
rect 56888 58410 56982 58850
rect 56888 58396 56914 58410
rect 56956 58396 56982 58410
rect 57582 58396 57670 58996
rect 45562 58338 45632 58396
rect 49556 58338 49626 58396
rect 53578 58338 53648 58396
rect 57600 58338 57670 58396
rect 42142 57738 42168 58338
rect 42768 58256 42794 58338
rect 42836 58256 42862 58338
rect 42768 57816 42862 58256
rect 42768 57738 42794 57816
rect 42836 57738 42862 57816
rect 43462 58278 43488 58338
rect 43530 58278 43556 58338
rect 43462 57838 43556 58278
rect 43462 57738 43488 57838
rect 43530 57738 43556 57838
rect 44156 58278 44182 58338
rect 44224 58278 44250 58338
rect 44156 57838 44250 58278
rect 44156 57738 44182 57838
rect 44224 57738 44250 57838
rect 44850 58266 44876 58338
rect 44918 58266 44944 58338
rect 44850 57826 44944 58266
rect 44850 57738 44876 57826
rect 44918 57738 44944 57826
rect 45544 58160 45632 58338
rect 46136 58160 46162 58338
rect 45544 57924 46162 58160
rect 45544 57738 45632 57924
rect 46136 57738 46162 57924
rect 46762 58256 46788 58338
rect 46830 58256 46856 58338
rect 46762 57816 46856 58256
rect 46762 57738 46788 57816
rect 46830 57738 46856 57816
rect 47456 58278 47482 58338
rect 47524 58278 47550 58338
rect 47456 57838 47550 58278
rect 47456 57738 47482 57838
rect 47524 57738 47550 57838
rect 48150 58278 48176 58338
rect 48218 58278 48244 58338
rect 48150 57838 48244 58278
rect 48150 57738 48176 57838
rect 48218 57738 48244 57838
rect 48844 58266 48870 58338
rect 48912 58266 48938 58338
rect 48844 57826 48938 58266
rect 48844 57738 48870 57826
rect 48912 57738 48938 57826
rect 49538 58160 49626 58338
rect 50158 58160 50184 58338
rect 49538 57924 50184 58160
rect 49538 57738 49626 57924
rect 50158 57738 50184 57924
rect 50784 58256 50810 58338
rect 50852 58256 50878 58338
rect 50784 57816 50878 58256
rect 50784 57738 50810 57816
rect 50852 57738 50878 57816
rect 51478 58278 51504 58338
rect 51546 58278 51572 58338
rect 51478 57838 51572 58278
rect 51478 57738 51504 57838
rect 51546 57738 51572 57838
rect 52172 58278 52198 58338
rect 52240 58278 52266 58338
rect 52172 57838 52266 58278
rect 52172 57738 52198 57838
rect 52240 57738 52266 57838
rect 52866 58266 52892 58338
rect 52934 58266 52960 58338
rect 52866 57826 52960 58266
rect 52866 57738 52892 57826
rect 52934 57738 52960 57826
rect 53560 58266 53648 58338
rect 54180 58266 54206 58338
rect 53560 58030 54206 58266
rect 53560 57738 53648 58030
rect 54180 57738 54206 58030
rect 54806 58256 54832 58338
rect 54874 58256 54900 58338
rect 54806 57816 54900 58256
rect 54806 57738 54832 57816
rect 54874 57738 54900 57816
rect 55500 58278 55526 58338
rect 55568 58278 55594 58338
rect 55500 57838 55594 58278
rect 55500 57738 55526 57838
rect 55568 57738 55594 57838
rect 56194 58278 56220 58338
rect 56262 58278 56288 58338
rect 56194 57838 56288 58278
rect 56194 57738 56220 57838
rect 56262 57738 56288 57838
rect 56888 58266 56914 58338
rect 56956 58266 56982 58338
rect 56888 57826 56982 58266
rect 56888 57738 56914 57826
rect 56956 57738 56982 57826
rect 57582 57738 57670 58338
rect 45562 57680 45632 57738
rect 49556 57680 49626 57738
rect 53578 57680 53648 57738
rect 57600 57680 57670 57738
rect 23394 56834 23420 57434
rect 24020 57232 24046 57434
rect 24088 57232 24114 57434
rect 24020 56968 24114 57232
rect 24020 56834 24046 56968
rect 24088 56834 24114 56968
rect 24714 57202 24740 57434
rect 24782 57202 24808 57434
rect 24714 56938 24808 57202
rect 24714 56834 24740 56938
rect 24782 56834 24808 56938
rect 25408 57214 25434 57434
rect 25476 57214 25502 57434
rect 25408 56950 25502 57214
rect 25408 56834 25434 56950
rect 25476 56834 25502 56950
rect 26102 57228 26128 57434
rect 26170 57228 26196 57434
rect 26102 56964 26196 57228
rect 26102 56834 26128 56964
rect 26170 56834 26196 56964
rect 26796 57230 26822 57434
rect 26864 57230 26890 57434
rect 26796 56966 26890 57230
rect 26796 56834 26822 56966
rect 26864 56834 26890 56966
rect 27490 57258 27516 57434
rect 27558 57258 27584 57434
rect 27490 56994 27584 57258
rect 27490 56834 27516 56994
rect 27558 56834 27584 56994
rect 28184 57272 28210 57434
rect 28252 57272 28278 57434
rect 28184 57008 28278 57272
rect 28184 56834 28210 57008
rect 28252 56834 28278 57008
rect 28878 57256 28904 57434
rect 28946 57256 28972 57434
rect 28878 56992 28972 57256
rect 28878 56834 28904 56992
rect 28946 56834 28972 56992
rect 29572 57278 29598 57434
rect 29640 57278 29666 57434
rect 29572 57014 29666 57278
rect 29572 56834 29598 57014
rect 29640 56834 29666 57014
rect 30266 57086 30292 57434
rect 30266 56854 30406 57086
rect 30266 56834 30340 56854
rect 30284 56776 30340 56834
rect 23394 56176 23420 56776
rect 24020 56532 24046 56776
rect 24088 56532 24114 56776
rect 24020 56268 24114 56532
rect 24020 56176 24046 56268
rect 24088 56176 24114 56268
rect 24714 56554 24740 56776
rect 24782 56554 24808 56776
rect 24714 56290 24808 56554
rect 24714 56176 24740 56290
rect 24782 56176 24808 56290
rect 25408 56500 25434 56776
rect 25476 56500 25502 56776
rect 25408 56236 25502 56500
rect 25408 56176 25434 56236
rect 25476 56176 25502 56236
rect 26102 56526 26128 56776
rect 26170 56526 26196 56776
rect 26102 56262 26196 56526
rect 26102 56176 26128 56262
rect 26170 56176 26196 56262
rect 26796 56508 26822 56776
rect 26864 56508 26890 56776
rect 26796 56244 26890 56508
rect 26796 56176 26822 56244
rect 26864 56176 26890 56244
rect 27490 56472 27516 56776
rect 27558 56472 27584 56776
rect 27490 56208 27584 56472
rect 27490 56176 27516 56208
rect 27558 56176 27584 56208
rect 28184 56522 28210 56776
rect 28252 56522 28278 56776
rect 28184 56258 28278 56522
rect 28184 56176 28210 56258
rect 28252 56176 28278 56258
rect 28878 56530 28904 56776
rect 28946 56530 28972 56776
rect 28878 56266 28972 56530
rect 28878 56176 28904 56266
rect 28946 56176 28972 56266
rect 29572 56586 29598 56776
rect 29640 56586 29666 56776
rect 29572 56322 29666 56586
rect 29572 56176 29598 56322
rect 29640 56176 29666 56322
rect 30266 56768 30340 56776
rect 30394 56768 30406 56854
rect 30266 56534 30406 56768
rect 30266 56530 30356 56534
rect 30266 56176 30292 56530
rect 23400 54944 23426 55544
rect 24026 55342 24052 55544
rect 24094 55342 24120 55544
rect 24026 55078 24120 55342
rect 24026 54944 24052 55078
rect 24094 54944 24120 55078
rect 24720 55312 24746 55544
rect 24788 55312 24814 55544
rect 24720 55048 24814 55312
rect 24720 54944 24746 55048
rect 24788 54944 24814 55048
rect 25414 55324 25440 55544
rect 25482 55324 25508 55544
rect 25414 55060 25508 55324
rect 25414 54944 25440 55060
rect 25482 54944 25508 55060
rect 26108 55338 26134 55544
rect 26176 55338 26202 55544
rect 26108 55074 26202 55338
rect 26108 54944 26134 55074
rect 26176 54944 26202 55074
rect 26802 55340 26828 55544
rect 26870 55340 26896 55544
rect 26802 55076 26896 55340
rect 26802 54944 26828 55076
rect 26870 54944 26896 55076
rect 27496 55368 27522 55544
rect 27564 55368 27590 55544
rect 27496 55104 27590 55368
rect 27496 54944 27522 55104
rect 27564 54944 27590 55104
rect 28190 55382 28216 55544
rect 28258 55382 28284 55544
rect 28190 55118 28284 55382
rect 28190 54944 28216 55118
rect 28258 54944 28284 55118
rect 28884 55366 28910 55544
rect 28952 55366 28978 55544
rect 28884 55102 28978 55366
rect 28884 54944 28910 55102
rect 28952 54944 28978 55102
rect 29578 55388 29604 55544
rect 29646 55388 29672 55544
rect 29578 55124 29672 55388
rect 29578 54944 29604 55124
rect 29646 54944 29672 55124
rect 30272 55196 30298 55544
rect 30272 55098 30362 55196
rect 30272 54944 30454 55098
rect 30290 54886 30454 54944
rect 23400 54810 23426 54886
rect 23258 54734 23426 54810
rect 23258 54418 23294 54734
rect 23382 54418 23426 54734
rect 23258 54332 23426 54418
rect 23400 54286 23426 54332
rect 24026 54642 24052 54886
rect 24094 54642 24120 54886
rect 24026 54378 24120 54642
rect 24026 54286 24052 54378
rect 24094 54286 24120 54378
rect 24720 54664 24746 54886
rect 24788 54664 24814 54886
rect 24720 54400 24814 54664
rect 24720 54286 24746 54400
rect 24788 54286 24814 54400
rect 25414 54610 25440 54886
rect 25482 54610 25508 54886
rect 25414 54346 25508 54610
rect 25414 54286 25440 54346
rect 25482 54286 25508 54346
rect 26108 54636 26134 54886
rect 26176 54636 26202 54886
rect 26108 54372 26202 54636
rect 26108 54286 26134 54372
rect 26176 54286 26202 54372
rect 26802 54618 26828 54886
rect 26870 54618 26896 54886
rect 26802 54354 26896 54618
rect 26802 54286 26828 54354
rect 26870 54286 26896 54354
rect 27496 54582 27522 54886
rect 27564 54582 27590 54886
rect 27496 54318 27590 54582
rect 27496 54286 27522 54318
rect 27564 54286 27590 54318
rect 28190 54632 28216 54886
rect 28258 54632 28284 54886
rect 28190 54368 28284 54632
rect 28190 54286 28216 54368
rect 28258 54286 28284 54368
rect 28884 54640 28910 54886
rect 28952 54640 28978 54886
rect 28884 54376 28978 54640
rect 28884 54286 28910 54376
rect 28952 54286 28978 54376
rect 29578 54696 29604 54886
rect 29646 54696 29672 54886
rect 29578 54432 29672 54696
rect 29578 54286 29604 54432
rect 29646 54286 29672 54432
rect 30272 54688 30454 54886
rect 30272 54640 30362 54688
rect 30272 54286 30298 54640
rect 23416 53002 23442 53602
rect 24042 53400 24068 53602
rect 24110 53400 24136 53602
rect 24042 53136 24136 53400
rect 24042 53002 24068 53136
rect 24110 53002 24136 53136
rect 24736 53370 24762 53602
rect 24804 53370 24830 53602
rect 24736 53106 24830 53370
rect 24736 53002 24762 53106
rect 24804 53002 24830 53106
rect 25430 53382 25456 53602
rect 25498 53382 25524 53602
rect 25430 53118 25524 53382
rect 25430 53002 25456 53118
rect 25498 53002 25524 53118
rect 26124 53396 26150 53602
rect 26192 53396 26218 53602
rect 26124 53132 26218 53396
rect 26124 53002 26150 53132
rect 26192 53002 26218 53132
rect 26818 53398 26844 53602
rect 26886 53398 26912 53602
rect 26818 53134 26912 53398
rect 26818 53002 26844 53134
rect 26886 53002 26912 53134
rect 27512 53426 27538 53602
rect 27580 53426 27606 53602
rect 27512 53162 27606 53426
rect 27512 53002 27538 53162
rect 27580 53002 27606 53162
rect 28206 53440 28232 53602
rect 28274 53440 28300 53602
rect 28206 53176 28300 53440
rect 28206 53002 28232 53176
rect 28274 53002 28300 53176
rect 28900 53424 28926 53602
rect 28968 53424 28994 53602
rect 28900 53160 28994 53424
rect 28900 53002 28926 53160
rect 28968 53002 28994 53160
rect 29594 53446 29620 53602
rect 29662 53446 29688 53602
rect 29594 53182 29688 53446
rect 29594 53002 29620 53182
rect 29662 53002 29688 53182
rect 30288 53254 30314 53602
rect 30288 53250 30378 53254
rect 30288 53076 30492 53250
rect 30288 53002 30374 53076
rect 30306 52944 30374 53002
rect 23416 52344 23442 52944
rect 24042 52700 24068 52944
rect 24110 52700 24136 52944
rect 24042 52436 24136 52700
rect 24042 52344 24068 52436
rect 24110 52344 24136 52436
rect 24736 52722 24762 52944
rect 24804 52722 24830 52944
rect 24736 52458 24830 52722
rect 24736 52344 24762 52458
rect 24804 52344 24830 52458
rect 25430 52668 25456 52944
rect 25498 52668 25524 52944
rect 25430 52404 25524 52668
rect 25430 52344 25456 52404
rect 25498 52344 25524 52404
rect 26124 52694 26150 52944
rect 26192 52694 26218 52944
rect 26124 52430 26218 52694
rect 26124 52344 26150 52430
rect 26192 52344 26218 52430
rect 26818 52676 26844 52944
rect 26886 52676 26912 52944
rect 26818 52412 26912 52676
rect 26818 52344 26844 52412
rect 26886 52344 26912 52412
rect 27512 52640 27538 52944
rect 27580 52640 27606 52944
rect 27512 52376 27606 52640
rect 27512 52344 27538 52376
rect 27580 52344 27606 52376
rect 28206 52690 28232 52944
rect 28274 52690 28300 52944
rect 28206 52426 28300 52690
rect 28206 52344 28232 52426
rect 28274 52344 28300 52426
rect 28900 52698 28926 52944
rect 28968 52698 28994 52944
rect 28900 52434 28994 52698
rect 28900 52344 28926 52434
rect 28968 52344 28994 52434
rect 29594 52754 29620 52944
rect 29662 52754 29688 52944
rect 29594 52490 29688 52754
rect 29594 52344 29620 52490
rect 29662 52344 29688 52490
rect 30288 52928 30374 52944
rect 30470 52928 30492 53076
rect 30288 52712 30492 52928
rect 30288 52698 30378 52712
rect 30288 52344 30314 52698
rect 42142 57080 42168 57680
rect 42768 57548 42794 57680
rect 42836 57548 42862 57680
rect 42768 57108 42862 57548
rect 42768 57080 42794 57108
rect 42836 57080 42862 57108
rect 43462 57590 43488 57680
rect 43530 57590 43556 57680
rect 43462 57150 43556 57590
rect 43462 57080 43488 57150
rect 43530 57080 43556 57150
rect 44156 57602 44182 57680
rect 44224 57602 44250 57680
rect 44156 57162 44250 57602
rect 44156 57080 44182 57162
rect 44224 57080 44250 57162
rect 44850 57628 44876 57680
rect 44918 57628 44944 57680
rect 44850 57188 44944 57628
rect 44850 57080 44876 57188
rect 44918 57080 44944 57188
rect 45544 57650 45632 57680
rect 46136 57650 46162 57680
rect 45544 57414 46162 57650
rect 45544 57400 45632 57414
rect 45544 57080 45570 57400
rect 46136 57080 46162 57414
rect 46762 57548 46788 57680
rect 46830 57548 46856 57680
rect 46762 57108 46856 57548
rect 46762 57080 46788 57108
rect 46830 57080 46856 57108
rect 47456 57590 47482 57680
rect 47524 57590 47550 57680
rect 47456 57150 47550 57590
rect 47456 57080 47482 57150
rect 47524 57080 47550 57150
rect 48150 57602 48176 57680
rect 48218 57602 48244 57680
rect 48150 57162 48244 57602
rect 48150 57080 48176 57162
rect 48218 57080 48244 57162
rect 48844 57628 48870 57680
rect 48912 57628 48938 57680
rect 48844 57188 48938 57628
rect 48844 57080 48870 57188
rect 48912 57080 48938 57188
rect 49538 57634 49626 57680
rect 50158 57634 50184 57680
rect 49538 57398 50184 57634
rect 49538 57080 49564 57398
rect 50158 57080 50184 57398
rect 50784 57548 50810 57680
rect 50852 57548 50878 57680
rect 50784 57108 50878 57548
rect 50784 57080 50810 57108
rect 50852 57080 50878 57108
rect 51478 57590 51504 57680
rect 51546 57590 51572 57680
rect 51478 57150 51572 57590
rect 51478 57080 51504 57150
rect 51546 57080 51572 57150
rect 52172 57602 52198 57680
rect 52240 57602 52266 57680
rect 52172 57162 52266 57602
rect 52172 57080 52198 57162
rect 52240 57080 52266 57162
rect 52866 57628 52892 57680
rect 52934 57628 52960 57680
rect 52866 57188 52960 57628
rect 52866 57080 52892 57188
rect 52934 57080 52960 57188
rect 53560 57664 53648 57680
rect 54180 57664 54206 57680
rect 53560 57428 54206 57664
rect 53560 57400 53648 57428
rect 53560 57080 53586 57400
rect 54180 57080 54206 57428
rect 54806 57548 54832 57680
rect 54874 57548 54900 57680
rect 54806 57108 54900 57548
rect 54806 57080 54832 57108
rect 54874 57080 54900 57108
rect 55500 57590 55526 57680
rect 55568 57590 55594 57680
rect 55500 57150 55594 57590
rect 55500 57080 55526 57150
rect 55568 57080 55594 57150
rect 56194 57602 56220 57680
rect 56262 57602 56288 57680
rect 56194 57162 56288 57602
rect 56194 57080 56220 57162
rect 56262 57080 56288 57162
rect 56888 57628 56914 57680
rect 56956 57628 56982 57680
rect 56888 57188 56982 57628
rect 56888 57080 56914 57188
rect 56956 57080 56982 57188
rect 57582 57400 57670 57680
rect 75216 62010 75816 62032
rect 75874 62010 76474 62032
rect 76532 62010 77132 62032
rect 77190 62010 77790 62032
rect 79066 62024 79666 62046
rect 79724 62024 80324 62046
rect 80382 62024 80982 62046
rect 81040 62024 81640 62046
rect 71352 61404 71952 61430
rect 72010 61404 72610 61430
rect 72668 61404 73268 61430
rect 73326 61404 73926 61430
rect 71412 61362 71836 61404
rect 72150 61362 72574 61404
rect 72732 61362 73156 61404
rect 73404 61362 73828 61404
rect 71352 61336 71952 61362
rect 72010 61336 72610 61362
rect 72668 61336 73268 61362
rect 73326 61336 73926 61362
rect 71352 60710 71952 60736
rect 72010 60710 72610 60736
rect 72668 60710 73268 60736
rect 73326 60710 73926 60736
rect 71406 60668 71830 60710
rect 72118 60668 72542 60710
rect 72728 60668 73152 60710
rect 73444 60668 73868 60710
rect 71352 60642 71952 60668
rect 72010 60642 72610 60668
rect 72668 60642 73268 60668
rect 73326 60642 73926 60668
rect 71352 60016 71952 60042
rect 72010 60016 72610 60042
rect 72668 60016 73268 60042
rect 73326 60016 73926 60042
rect 71392 59974 71816 60016
rect 72138 59974 72562 60016
rect 72766 59974 73190 60016
rect 73402 59974 73826 60016
rect 71352 59948 71952 59974
rect 72010 59948 72610 59974
rect 72668 59948 73268 59974
rect 73326 59948 73926 59974
rect 71352 59322 71952 59348
rect 72010 59322 72610 59348
rect 72668 59322 73268 59348
rect 73326 59322 73926 59348
rect 71388 59280 71812 59322
rect 72168 59280 72592 59322
rect 72718 59280 73142 59322
rect 73436 59280 73860 59322
rect 71352 59254 71952 59280
rect 72010 59254 72610 59280
rect 72668 59254 73268 59280
rect 73326 59254 73926 59280
rect 75216 61384 75816 61410
rect 75874 61384 76474 61410
rect 76532 61384 77132 61410
rect 77190 61384 77790 61410
rect 75276 61342 75700 61384
rect 76014 61342 76438 61384
rect 76596 61342 77020 61384
rect 77268 61342 77692 61384
rect 75216 61316 75816 61342
rect 75874 61316 76474 61342
rect 76532 61316 77132 61342
rect 77190 61316 77790 61342
rect 75216 60690 75816 60716
rect 75874 60690 76474 60716
rect 76532 60690 77132 60716
rect 77190 60690 77790 60716
rect 75270 60648 75694 60690
rect 75982 60648 76406 60690
rect 76592 60648 77016 60690
rect 77308 60648 77732 60690
rect 75216 60622 75816 60648
rect 75874 60622 76474 60648
rect 76532 60622 77132 60648
rect 77190 60622 77790 60648
rect 75216 59996 75816 60022
rect 75874 59996 76474 60022
rect 76532 59996 77132 60022
rect 77190 59996 77790 60022
rect 75256 59954 75680 59996
rect 76002 59954 76426 59996
rect 76630 59954 77054 59996
rect 77266 59954 77690 59996
rect 75216 59928 75816 59954
rect 75874 59928 76474 59954
rect 76532 59928 77132 59954
rect 77190 59928 77790 59954
rect 75216 59302 75816 59328
rect 75874 59302 76474 59328
rect 76532 59302 77132 59328
rect 77190 59302 77790 59328
rect 75252 59260 75676 59302
rect 76032 59260 76456 59302
rect 76582 59260 77006 59302
rect 77300 59260 77724 59302
rect 75216 59234 75816 59260
rect 75874 59234 76474 59260
rect 76532 59234 77132 59260
rect 77190 59234 77790 59260
rect 71352 58628 71952 58654
rect 72010 58628 72610 58654
rect 72668 58628 73268 58654
rect 73326 58628 73926 58654
rect 79066 61398 79666 61424
rect 79724 61398 80324 61424
rect 80382 61398 80982 61424
rect 81040 61398 81640 61424
rect 79126 61356 79550 61398
rect 79864 61356 80288 61398
rect 80446 61356 80870 61398
rect 81118 61356 81542 61398
rect 79066 61330 79666 61356
rect 79724 61330 80324 61356
rect 80382 61330 80982 61356
rect 81040 61330 81640 61356
rect 79066 60704 79666 60730
rect 79724 60704 80324 60730
rect 80382 60704 80982 60730
rect 81040 60704 81640 60730
rect 79120 60662 79544 60704
rect 79832 60662 80256 60704
rect 80442 60662 80866 60704
rect 81158 60662 81582 60704
rect 79066 60636 79666 60662
rect 79724 60636 80324 60662
rect 80382 60636 80982 60662
rect 81040 60636 81640 60662
rect 79066 60010 79666 60036
rect 79724 60010 80324 60036
rect 80382 60010 80982 60036
rect 81040 60010 81640 60036
rect 79106 59968 79530 60010
rect 79852 59968 80276 60010
rect 80480 59968 80904 60010
rect 81116 59968 81540 60010
rect 79066 59942 79666 59968
rect 79724 59942 80324 59968
rect 80382 59942 80982 59968
rect 81040 59942 81640 59968
rect 79066 59316 79666 59342
rect 79724 59316 80324 59342
rect 80382 59316 80982 59342
rect 81040 59316 81640 59342
rect 79102 59274 79526 59316
rect 79882 59274 80306 59316
rect 80432 59274 80856 59316
rect 81150 59274 81574 59316
rect 79066 59248 79666 59274
rect 79724 59248 80324 59274
rect 80382 59248 80982 59274
rect 81040 59248 81640 59274
rect 71722 58346 71818 58628
rect 72190 58346 72286 58628
rect 72800 58346 72896 58628
rect 73490 58346 73586 58628
rect 75216 58608 75816 58634
rect 75874 58608 76474 58634
rect 76532 58608 77132 58634
rect 77190 58608 77790 58634
rect 79066 58622 79666 58648
rect 79724 58622 80324 58648
rect 80382 58622 80982 58648
rect 81040 58622 81640 58648
rect 71698 58280 73788 58346
rect 75586 58326 75682 58608
rect 76054 58326 76150 58608
rect 76664 58326 76760 58608
rect 77354 58326 77450 58608
rect 79436 58340 79532 58622
rect 79904 58340 80000 58622
rect 80514 58340 80610 58622
rect 81204 58340 81300 58622
rect 71352 58276 73926 58280
rect 71352 58254 71952 58276
rect 72010 58254 72610 58276
rect 72668 58254 73268 58276
rect 73326 58254 73926 58276
rect 75562 58260 77652 58326
rect 79412 58274 81502 58340
rect 79066 58270 81640 58274
rect 75216 58256 77790 58260
rect 57582 57080 57608 57400
rect 42094 55322 42120 55922
rect 42720 55844 42746 55922
rect 42788 55844 42814 55922
rect 42720 55404 42814 55844
rect 42720 55322 42746 55404
rect 42788 55322 42814 55404
rect 43414 55842 43440 55922
rect 43482 55842 43508 55922
rect 43414 55402 43508 55842
rect 43414 55322 43440 55402
rect 43482 55322 43508 55402
rect 44108 55856 44134 55922
rect 44176 55856 44202 55922
rect 44108 55416 44202 55856
rect 44108 55322 44134 55416
rect 44176 55322 44202 55416
rect 44802 55836 44828 55922
rect 44870 55836 44896 55922
rect 44802 55390 44896 55836
rect 44802 55322 44828 55390
rect 44870 55322 44896 55390
rect 45496 55676 45522 55922
rect 45496 55652 45584 55676
rect 46102 55652 46128 55920
rect 45496 55418 46128 55652
rect 45496 55322 45584 55418
rect 45514 55264 45584 55322
rect 46102 55320 46128 55418
rect 46728 55842 46754 55920
rect 46796 55842 46822 55920
rect 46728 55402 46822 55842
rect 46728 55320 46754 55402
rect 46796 55320 46822 55402
rect 47422 55840 47448 55920
rect 47490 55840 47516 55920
rect 47422 55400 47516 55840
rect 47422 55320 47448 55400
rect 47490 55320 47516 55400
rect 48116 55854 48142 55920
rect 48184 55854 48210 55920
rect 48116 55414 48210 55854
rect 48116 55320 48142 55414
rect 48184 55320 48210 55414
rect 48810 55834 48836 55920
rect 48878 55834 48904 55920
rect 48810 55388 48904 55834
rect 48810 55320 48836 55388
rect 48878 55320 48904 55388
rect 49504 55674 49530 55920
rect 49504 55656 49592 55674
rect 50114 55656 50140 55920
rect 49504 55422 50140 55656
rect 49504 55320 49592 55422
rect 50114 55320 50140 55422
rect 50740 55842 50766 55920
rect 50808 55842 50834 55920
rect 50740 55402 50834 55842
rect 50740 55320 50766 55402
rect 50808 55320 50834 55402
rect 51434 55840 51460 55920
rect 51502 55840 51528 55920
rect 51434 55400 51528 55840
rect 51434 55320 51460 55400
rect 51502 55320 51528 55400
rect 52128 55854 52154 55920
rect 52196 55854 52222 55920
rect 52128 55414 52222 55854
rect 52128 55320 52154 55414
rect 52196 55320 52222 55414
rect 52822 55834 52848 55920
rect 52890 55834 52916 55920
rect 52822 55388 52916 55834
rect 52822 55320 52848 55388
rect 52890 55320 52916 55388
rect 53516 55674 53542 55920
rect 53516 55646 53604 55674
rect 54124 55646 54150 55920
rect 53516 55412 54150 55646
rect 53516 55320 53604 55412
rect 54124 55320 54150 55412
rect 54750 55842 54776 55920
rect 54818 55842 54844 55920
rect 54750 55402 54844 55842
rect 54750 55320 54776 55402
rect 54818 55320 54844 55402
rect 55444 55840 55470 55920
rect 55512 55840 55538 55920
rect 55444 55400 55538 55840
rect 55444 55320 55470 55400
rect 55512 55320 55538 55400
rect 56138 55854 56164 55920
rect 56206 55854 56232 55920
rect 56138 55414 56232 55854
rect 56138 55320 56164 55414
rect 56206 55320 56232 55414
rect 56832 55834 56858 55920
rect 56900 55834 56926 55920
rect 56832 55388 56926 55834
rect 56832 55320 56858 55388
rect 56900 55320 56926 55388
rect 57526 55674 57552 55920
rect 57526 55320 57614 55674
rect 42094 54664 42120 55264
rect 42720 55174 42746 55264
rect 42788 55174 42814 55264
rect 42720 54734 42814 55174
rect 42720 54664 42746 54734
rect 42788 54664 42814 54734
rect 43414 55198 43440 55264
rect 43482 55198 43508 55264
rect 43414 54758 43508 55198
rect 43414 54664 43440 54758
rect 43482 54664 43508 54758
rect 44108 55182 44134 55264
rect 44176 55182 44202 55264
rect 44108 54742 44202 55182
rect 44108 54664 44134 54742
rect 44176 54664 44202 54742
rect 44802 55194 44828 55264
rect 44870 55194 44896 55264
rect 44802 54754 44896 55194
rect 44802 54664 44828 54754
rect 44870 54664 44896 54754
rect 45496 55146 45584 55264
rect 49522 55262 49592 55320
rect 53534 55262 53604 55320
rect 57544 55262 57614 55320
rect 46102 55146 46128 55262
rect 45496 54912 46128 55146
rect 45496 54664 45584 54912
rect 45514 54606 45584 54664
rect 46102 54662 46128 54912
rect 46728 55172 46754 55262
rect 46796 55172 46822 55262
rect 46728 54732 46822 55172
rect 46728 54662 46754 54732
rect 46796 54662 46822 54732
rect 47422 55196 47448 55262
rect 47490 55196 47516 55262
rect 47422 54756 47516 55196
rect 47422 54662 47448 54756
rect 47490 54662 47516 54756
rect 48116 55180 48142 55262
rect 48184 55180 48210 55262
rect 48116 54740 48210 55180
rect 48116 54662 48142 54740
rect 48184 54662 48210 54740
rect 48810 55192 48836 55262
rect 48878 55192 48904 55262
rect 48810 54752 48904 55192
rect 48810 54662 48836 54752
rect 48878 54662 48904 54752
rect 49504 55146 49592 55262
rect 50114 55146 50140 55262
rect 49504 54912 50140 55146
rect 49504 54662 49592 54912
rect 50114 54662 50140 54912
rect 50740 55172 50766 55262
rect 50808 55172 50834 55262
rect 50740 54732 50834 55172
rect 50740 54662 50766 54732
rect 50808 54662 50834 54732
rect 51434 55196 51460 55262
rect 51502 55196 51528 55262
rect 51434 54756 51528 55196
rect 51434 54662 51460 54756
rect 51502 54662 51528 54756
rect 52128 55180 52154 55262
rect 52196 55180 52222 55262
rect 52128 54740 52222 55180
rect 52128 54662 52154 54740
rect 52196 54662 52222 54740
rect 52822 55192 52848 55262
rect 52890 55192 52916 55262
rect 52822 54752 52916 55192
rect 52822 54662 52848 54752
rect 52890 54662 52916 54752
rect 53516 55188 53604 55262
rect 54124 55188 54150 55262
rect 53516 54954 54150 55188
rect 53516 54662 53604 54954
rect 54124 54662 54150 54954
rect 54750 55172 54776 55262
rect 54818 55172 54844 55262
rect 54750 54732 54844 55172
rect 54750 54662 54776 54732
rect 54818 54662 54844 54732
rect 55444 55196 55470 55262
rect 55512 55196 55538 55262
rect 55444 54756 55538 55196
rect 55444 54662 55470 54756
rect 55512 54662 55538 54756
rect 56138 55180 56164 55262
rect 56206 55180 56232 55262
rect 56138 54740 56232 55180
rect 56138 54662 56164 54740
rect 56206 54662 56232 54740
rect 56832 55192 56858 55262
rect 56900 55192 56926 55262
rect 56832 54752 56926 55192
rect 56832 54662 56858 54752
rect 56900 54662 56926 54752
rect 57526 54662 57614 55262
rect 42094 54006 42120 54606
rect 42720 54498 42746 54606
rect 42788 54498 42814 54606
rect 42720 54058 42814 54498
rect 42720 54006 42746 54058
rect 42788 54006 42814 54058
rect 43414 54510 43440 54606
rect 43482 54510 43508 54606
rect 43414 54070 43508 54510
rect 43414 54006 43440 54070
rect 43482 54006 43508 54070
rect 44108 54488 44134 54606
rect 44176 54488 44202 54606
rect 44108 54048 44202 54488
rect 44108 54006 44134 54048
rect 44176 54006 44202 54048
rect 44802 54460 44828 54606
rect 44870 54460 44896 54606
rect 44802 54020 44896 54460
rect 44802 54006 44828 54020
rect 44870 54006 44896 54020
rect 45496 54468 45584 54606
rect 49522 54604 49592 54662
rect 53534 54604 53604 54662
rect 57544 54604 57614 54662
rect 46102 54468 46128 54604
rect 45496 54234 46128 54468
rect 45496 54006 45584 54234
rect 45514 53948 45584 54006
rect 46102 54004 46128 54234
rect 46728 54496 46754 54604
rect 46796 54496 46822 54604
rect 46728 54056 46822 54496
rect 46728 54004 46754 54056
rect 46796 54004 46822 54056
rect 47422 54508 47448 54604
rect 47490 54508 47516 54604
rect 47422 54068 47516 54508
rect 47422 54004 47448 54068
rect 47490 54004 47516 54068
rect 48116 54486 48142 54604
rect 48184 54486 48210 54604
rect 48116 54046 48210 54486
rect 48116 54004 48142 54046
rect 48184 54004 48210 54046
rect 48810 54458 48836 54604
rect 48878 54458 48904 54604
rect 48810 54018 48904 54458
rect 48810 54004 48836 54018
rect 48878 54004 48904 54018
rect 49504 54474 49592 54604
rect 50114 54474 50140 54604
rect 49504 54240 50140 54474
rect 49504 54004 49592 54240
rect 50114 54004 50140 54240
rect 50740 54496 50766 54604
rect 50808 54496 50834 54604
rect 50740 54056 50834 54496
rect 50740 54004 50766 54056
rect 50808 54004 50834 54056
rect 51434 54508 51460 54604
rect 51502 54508 51528 54604
rect 51434 54068 51528 54508
rect 51434 54004 51460 54068
rect 51502 54004 51528 54068
rect 52128 54486 52154 54604
rect 52196 54486 52222 54604
rect 52128 54046 52222 54486
rect 52128 54004 52154 54046
rect 52196 54004 52222 54046
rect 52822 54458 52848 54604
rect 52890 54458 52916 54604
rect 52822 54018 52916 54458
rect 52822 54004 52848 54018
rect 52890 54004 52916 54018
rect 53516 54458 53604 54604
rect 54124 54458 54150 54604
rect 53516 54224 54150 54458
rect 53516 54004 53604 54224
rect 54124 54004 54150 54224
rect 54750 54496 54776 54604
rect 54818 54496 54844 54604
rect 54750 54056 54844 54496
rect 54750 54004 54776 54056
rect 54818 54004 54844 54056
rect 55444 54508 55470 54604
rect 55512 54508 55538 54604
rect 55444 54068 55538 54508
rect 55444 54004 55470 54068
rect 55512 54004 55538 54068
rect 56138 54486 56164 54604
rect 56206 54486 56232 54604
rect 56138 54046 56232 54486
rect 56138 54004 56164 54046
rect 56206 54004 56232 54046
rect 56832 54458 56858 54604
rect 56900 54458 56926 54604
rect 56832 54018 56926 54458
rect 56832 54004 56858 54018
rect 56900 54004 56926 54018
rect 57526 54004 57614 54604
rect 42094 53348 42120 53948
rect 42720 53866 42746 53948
rect 42788 53866 42814 53948
rect 42720 53426 42814 53866
rect 42720 53348 42746 53426
rect 42788 53348 42814 53426
rect 43414 53888 43440 53948
rect 43482 53888 43508 53948
rect 43414 53448 43508 53888
rect 43414 53348 43440 53448
rect 43482 53348 43508 53448
rect 44108 53888 44134 53948
rect 44176 53888 44202 53948
rect 44108 53448 44202 53888
rect 44108 53348 44134 53448
rect 44176 53348 44202 53448
rect 44802 53876 44828 53948
rect 44870 53876 44896 53948
rect 44802 53436 44896 53876
rect 44802 53348 44828 53436
rect 44870 53348 44896 53436
rect 45496 53866 45584 53948
rect 49522 53946 49592 54004
rect 53534 53946 53604 54004
rect 57544 53946 57614 54004
rect 46102 53866 46128 53946
rect 45496 53632 46128 53866
rect 45496 53348 45584 53632
rect 45514 53290 45584 53348
rect 46102 53346 46128 53632
rect 46728 53864 46754 53946
rect 46796 53864 46822 53946
rect 46728 53424 46822 53864
rect 46728 53346 46754 53424
rect 46796 53346 46822 53424
rect 47422 53886 47448 53946
rect 47490 53886 47516 53946
rect 47422 53446 47516 53886
rect 47422 53346 47448 53446
rect 47490 53346 47516 53446
rect 48116 53886 48142 53946
rect 48184 53886 48210 53946
rect 48116 53446 48210 53886
rect 48116 53346 48142 53446
rect 48184 53346 48210 53446
rect 48810 53874 48836 53946
rect 48878 53874 48904 53946
rect 48810 53434 48904 53874
rect 48810 53346 48836 53434
rect 48878 53346 48904 53434
rect 49504 53832 49592 53946
rect 50114 53832 50140 53946
rect 49504 53598 50140 53832
rect 49504 53346 49592 53598
rect 50114 53346 50140 53598
rect 50740 53864 50766 53946
rect 50808 53864 50834 53946
rect 50740 53424 50834 53864
rect 50740 53346 50766 53424
rect 50808 53346 50834 53424
rect 51434 53886 51460 53946
rect 51502 53886 51528 53946
rect 51434 53446 51528 53886
rect 51434 53346 51460 53446
rect 51502 53346 51528 53446
rect 52128 53886 52154 53946
rect 52196 53886 52222 53946
rect 52128 53446 52222 53886
rect 52128 53346 52154 53446
rect 52196 53346 52222 53446
rect 52822 53874 52848 53946
rect 52890 53874 52916 53946
rect 52822 53434 52916 53874
rect 52822 53346 52848 53434
rect 52890 53346 52916 53434
rect 53516 53856 53604 53946
rect 54124 53856 54150 53946
rect 53516 53622 54150 53856
rect 53516 53346 53604 53622
rect 54124 53346 54150 53622
rect 54750 53864 54776 53946
rect 54818 53864 54844 53946
rect 54750 53424 54844 53864
rect 54750 53346 54776 53424
rect 54818 53346 54844 53424
rect 55444 53886 55470 53946
rect 55512 53886 55538 53946
rect 55444 53446 55538 53886
rect 55444 53346 55470 53446
rect 55512 53346 55538 53446
rect 56138 53886 56164 53946
rect 56206 53886 56232 53946
rect 56138 53446 56232 53886
rect 56138 53346 56164 53446
rect 56206 53346 56232 53446
rect 56832 53874 56858 53946
rect 56900 53874 56926 53946
rect 56832 53434 56926 53874
rect 56832 53346 56858 53434
rect 56900 53346 56926 53434
rect 57526 53364 57614 53946
rect 75216 58234 75816 58256
rect 75874 58234 76474 58256
rect 76532 58234 77132 58256
rect 77190 58234 77790 58256
rect 79066 58248 79666 58270
rect 79724 58248 80324 58270
rect 80382 58248 80982 58270
rect 81040 58248 81640 58270
rect 71352 57628 71952 57654
rect 72010 57628 72610 57654
rect 72668 57628 73268 57654
rect 73326 57628 73926 57654
rect 71412 57586 71836 57628
rect 72150 57586 72574 57628
rect 72732 57586 73156 57628
rect 73404 57586 73828 57628
rect 71352 57560 71952 57586
rect 72010 57560 72610 57586
rect 72668 57560 73268 57586
rect 73326 57560 73926 57586
rect 71352 56934 71952 56960
rect 72010 56934 72610 56960
rect 72668 56934 73268 56960
rect 73326 56934 73926 56960
rect 71406 56892 71830 56934
rect 72118 56892 72542 56934
rect 72728 56892 73152 56934
rect 73444 56892 73868 56934
rect 71352 56866 71952 56892
rect 72010 56866 72610 56892
rect 72668 56866 73268 56892
rect 73326 56866 73926 56892
rect 71352 56240 71952 56266
rect 72010 56240 72610 56266
rect 72668 56240 73268 56266
rect 73326 56240 73926 56266
rect 71392 56198 71816 56240
rect 72138 56198 72562 56240
rect 72766 56198 73190 56240
rect 73402 56198 73826 56240
rect 71352 56172 71952 56198
rect 72010 56172 72610 56198
rect 72668 56172 73268 56198
rect 73326 56172 73926 56198
rect 71352 55546 71952 55572
rect 72010 55546 72610 55572
rect 72668 55546 73268 55572
rect 73326 55546 73926 55572
rect 71388 55504 71812 55546
rect 72168 55504 72592 55546
rect 72718 55504 73142 55546
rect 73436 55504 73860 55546
rect 71352 55478 71952 55504
rect 72010 55478 72610 55504
rect 72668 55478 73268 55504
rect 73326 55478 73926 55504
rect 75216 57608 75816 57634
rect 75874 57608 76474 57634
rect 76532 57608 77132 57634
rect 77190 57608 77790 57634
rect 75276 57566 75700 57608
rect 76014 57566 76438 57608
rect 76596 57566 77020 57608
rect 77268 57566 77692 57608
rect 75216 57540 75816 57566
rect 75874 57540 76474 57566
rect 76532 57540 77132 57566
rect 77190 57540 77790 57566
rect 75216 56914 75816 56940
rect 75874 56914 76474 56940
rect 76532 56914 77132 56940
rect 77190 56914 77790 56940
rect 75270 56872 75694 56914
rect 75982 56872 76406 56914
rect 76592 56872 77016 56914
rect 77308 56872 77732 56914
rect 75216 56846 75816 56872
rect 75874 56846 76474 56872
rect 76532 56846 77132 56872
rect 77190 56846 77790 56872
rect 75216 56220 75816 56246
rect 75874 56220 76474 56246
rect 76532 56220 77132 56246
rect 77190 56220 77790 56246
rect 75256 56178 75680 56220
rect 76002 56178 76426 56220
rect 76630 56178 77054 56220
rect 77266 56178 77690 56220
rect 75216 56152 75816 56178
rect 75874 56152 76474 56178
rect 76532 56152 77132 56178
rect 77190 56152 77790 56178
rect 75216 55526 75816 55552
rect 75874 55526 76474 55552
rect 76532 55526 77132 55552
rect 77190 55526 77790 55552
rect 75252 55484 75676 55526
rect 76032 55484 76456 55526
rect 76582 55484 77006 55526
rect 77300 55484 77724 55526
rect 75216 55458 75816 55484
rect 75874 55458 76474 55484
rect 76532 55458 77132 55484
rect 77190 55458 77790 55484
rect 71352 54852 71952 54878
rect 72010 54852 72610 54878
rect 72668 54852 73268 54878
rect 73326 54852 73926 54878
rect 79066 57622 79666 57648
rect 79724 57622 80324 57648
rect 80382 57622 80982 57648
rect 81040 57622 81640 57648
rect 79126 57580 79550 57622
rect 79864 57580 80288 57622
rect 80446 57580 80870 57622
rect 81118 57580 81542 57622
rect 79066 57554 79666 57580
rect 79724 57554 80324 57580
rect 80382 57554 80982 57580
rect 81040 57554 81640 57580
rect 79066 56928 79666 56954
rect 79724 56928 80324 56954
rect 80382 56928 80982 56954
rect 81040 56928 81640 56954
rect 79120 56886 79544 56928
rect 79832 56886 80256 56928
rect 80442 56886 80866 56928
rect 81158 56886 81582 56928
rect 79066 56860 79666 56886
rect 79724 56860 80324 56886
rect 80382 56860 80982 56886
rect 81040 56860 81640 56886
rect 79066 56234 79666 56260
rect 79724 56234 80324 56260
rect 80382 56234 80982 56260
rect 81040 56234 81640 56260
rect 79106 56192 79530 56234
rect 79852 56192 80276 56234
rect 80480 56192 80904 56234
rect 81116 56192 81540 56234
rect 79066 56166 79666 56192
rect 79724 56166 80324 56192
rect 80382 56166 80982 56192
rect 81040 56166 81640 56192
rect 79066 55540 79666 55566
rect 79724 55540 80324 55566
rect 80382 55540 80982 55566
rect 81040 55540 81640 55566
rect 79102 55498 79526 55540
rect 79882 55498 80306 55540
rect 80432 55498 80856 55540
rect 81150 55498 81574 55540
rect 79066 55472 79666 55498
rect 79724 55472 80324 55498
rect 80382 55472 80982 55498
rect 81040 55472 81640 55498
rect 71746 54574 71842 54852
rect 72174 54574 72270 54852
rect 72850 54574 72946 54852
rect 73512 54574 73608 54852
rect 75216 54832 75816 54858
rect 75874 54832 76474 54858
rect 76532 54832 77132 54858
rect 77190 54832 77790 54858
rect 79066 54846 79666 54872
rect 79724 54846 80324 54872
rect 80382 54846 80982 54872
rect 81040 54846 81640 54872
rect 71702 54508 73792 54574
rect 75610 54554 75706 54832
rect 76038 54554 76134 54832
rect 76714 54554 76810 54832
rect 77376 54554 77472 54832
rect 79460 54568 79556 54846
rect 79888 54568 79984 54846
rect 80564 54568 80660 54846
rect 81226 54568 81322 54846
rect 71356 54504 73930 54508
rect 71356 54482 71956 54504
rect 72014 54482 72614 54504
rect 72672 54482 73272 54504
rect 73330 54482 73930 54504
rect 75566 54488 77656 54554
rect 79416 54502 81506 54568
rect 79070 54498 81644 54502
rect 75220 54484 77794 54488
rect 57526 53346 57804 53364
rect 42094 52690 42120 53290
rect 42720 53158 42746 53290
rect 42788 53158 42814 53290
rect 42720 52718 42814 53158
rect 42720 52690 42746 52718
rect 42788 52690 42814 52718
rect 43414 53200 43440 53290
rect 43482 53200 43508 53290
rect 43414 52760 43508 53200
rect 43414 52690 43440 52760
rect 43482 52690 43508 52760
rect 44108 53212 44134 53290
rect 44176 53212 44202 53290
rect 44108 52772 44202 53212
rect 44108 52690 44134 52772
rect 44176 52690 44202 52772
rect 44802 53238 44828 53290
rect 44870 53238 44896 53290
rect 44802 52798 44896 53238
rect 44802 52690 44828 52798
rect 44870 52690 44896 52798
rect 45496 53264 45584 53290
rect 49522 53288 49592 53346
rect 53534 53288 53604 53346
rect 57544 53288 57804 53346
rect 46102 53264 46128 53288
rect 45496 53030 46128 53264
rect 45496 53010 45584 53030
rect 45496 52690 45522 53010
rect 46102 52688 46128 53030
rect 46728 53156 46754 53288
rect 46796 53156 46822 53288
rect 46728 52716 46822 53156
rect 46728 52688 46754 52716
rect 46796 52688 46822 52716
rect 47422 53198 47448 53288
rect 47490 53198 47516 53288
rect 47422 52758 47516 53198
rect 47422 52688 47448 52758
rect 47490 52688 47516 52758
rect 48116 53210 48142 53288
rect 48184 53210 48210 53288
rect 48116 52770 48210 53210
rect 48116 52688 48142 52770
rect 48184 52688 48210 52770
rect 48810 53236 48836 53288
rect 48878 53236 48904 53288
rect 48810 52796 48904 53236
rect 48810 52688 48836 52796
rect 48878 52688 48904 52796
rect 49504 53240 49592 53288
rect 50114 53240 50140 53288
rect 49504 53006 50140 53240
rect 49504 52688 49530 53006
rect 50114 52688 50140 53006
rect 50740 53156 50766 53288
rect 50808 53156 50834 53288
rect 50740 52716 50834 53156
rect 50740 52688 50766 52716
rect 50808 52688 50834 52716
rect 51434 53198 51460 53288
rect 51502 53198 51528 53288
rect 51434 52758 51528 53198
rect 51434 52688 51460 52758
rect 51502 52688 51528 52758
rect 52128 53210 52154 53288
rect 52196 53210 52222 53288
rect 52128 52770 52222 53210
rect 52128 52688 52154 52770
rect 52196 52688 52222 52770
rect 52822 53236 52848 53288
rect 52890 53236 52916 53288
rect 52822 52796 52916 53236
rect 52822 52688 52848 52796
rect 52890 52688 52916 52796
rect 53516 53284 53604 53288
rect 54124 53284 54150 53288
rect 53516 53050 54150 53284
rect 53516 53008 53604 53050
rect 53516 52688 53542 53008
rect 54124 52688 54150 53050
rect 54750 53156 54776 53288
rect 54818 53156 54844 53288
rect 54750 52716 54844 53156
rect 54750 52688 54776 52716
rect 54818 52688 54844 52716
rect 55444 53198 55470 53288
rect 55512 53198 55538 53288
rect 55444 52758 55538 53198
rect 55444 52688 55470 52758
rect 55512 52688 55538 52758
rect 56138 53210 56164 53288
rect 56206 53210 56232 53288
rect 56138 52770 56232 53210
rect 56138 52688 56164 52770
rect 56206 52688 56232 52770
rect 56832 53236 56858 53288
rect 56900 53236 56926 53288
rect 56832 52796 56926 53236
rect 56832 52688 56858 52796
rect 56900 52688 56926 52796
rect 57526 53008 57804 53288
rect 57526 52688 57552 53008
rect 57602 52376 57804 53008
rect 57602 51974 57626 52376
rect 57772 51974 57804 52376
rect 42086 51124 42112 51724
rect 42712 51646 42738 51724
rect 42780 51646 42806 51724
rect 42712 51206 42806 51646
rect 42712 51124 42738 51206
rect 42780 51124 42806 51206
rect 43406 51644 43432 51724
rect 43474 51644 43500 51724
rect 43406 51204 43500 51644
rect 43406 51124 43432 51204
rect 43474 51124 43500 51204
rect 44100 51658 44126 51724
rect 44168 51658 44194 51724
rect 44100 51218 44194 51658
rect 44100 51124 44126 51218
rect 44168 51124 44194 51218
rect 44794 51638 44820 51724
rect 44862 51638 44888 51724
rect 44794 51192 44888 51638
rect 44794 51124 44820 51192
rect 44862 51124 44888 51192
rect 45488 51478 45514 51724
rect 45488 51442 45576 51478
rect 46080 51442 46106 51724
rect 45488 51206 46106 51442
rect 45488 51124 45576 51206
rect 46080 51124 46106 51206
rect 46706 51646 46732 51724
rect 46774 51646 46800 51724
rect 46706 51206 46800 51646
rect 46706 51124 46732 51206
rect 46774 51124 46800 51206
rect 47400 51644 47426 51724
rect 47468 51644 47494 51724
rect 47400 51204 47494 51644
rect 47400 51124 47426 51204
rect 47468 51124 47494 51204
rect 48094 51658 48120 51724
rect 48162 51658 48188 51724
rect 48094 51218 48188 51658
rect 48094 51124 48120 51218
rect 48162 51124 48188 51218
rect 48788 51638 48814 51724
rect 48856 51638 48882 51724
rect 48788 51192 48882 51638
rect 48788 51124 48814 51192
rect 48856 51124 48882 51192
rect 49482 51478 49508 51724
rect 49482 51438 49570 51478
rect 50102 51438 50128 51724
rect 49482 51202 50128 51438
rect 49482 51124 49570 51202
rect 50102 51124 50128 51202
rect 50728 51646 50754 51724
rect 50796 51646 50822 51724
rect 50728 51206 50822 51646
rect 50728 51124 50754 51206
rect 50796 51124 50822 51206
rect 51422 51644 51448 51724
rect 51490 51644 51516 51724
rect 51422 51204 51516 51644
rect 51422 51124 51448 51204
rect 51490 51124 51516 51204
rect 52116 51658 52142 51724
rect 52184 51658 52210 51724
rect 52116 51218 52210 51658
rect 52116 51124 52142 51218
rect 52184 51124 52210 51218
rect 52810 51638 52836 51724
rect 52878 51638 52904 51724
rect 52810 51192 52904 51638
rect 52810 51124 52836 51192
rect 52878 51124 52904 51192
rect 53504 51478 53530 51724
rect 53504 51438 53592 51478
rect 54124 51438 54150 51724
rect 53504 51202 54150 51438
rect 53504 51124 53592 51202
rect 54124 51124 54150 51202
rect 54750 51646 54776 51724
rect 54818 51646 54844 51724
rect 54750 51206 54844 51646
rect 54750 51124 54776 51206
rect 54818 51124 54844 51206
rect 55444 51644 55470 51724
rect 55512 51644 55538 51724
rect 55444 51204 55538 51644
rect 55444 51124 55470 51204
rect 55512 51124 55538 51204
rect 56138 51658 56164 51724
rect 56206 51658 56232 51724
rect 56138 51218 56232 51658
rect 56138 51124 56164 51218
rect 56206 51124 56232 51218
rect 56832 51638 56858 51724
rect 56900 51638 56926 51724
rect 56832 51192 56926 51638
rect 56832 51124 56858 51192
rect 56900 51124 56926 51192
rect 57526 51478 57552 51724
rect 57602 51478 57804 51974
rect 57526 51246 57804 51478
rect 75220 54462 75820 54484
rect 75878 54462 76478 54484
rect 76536 54462 77136 54484
rect 77194 54462 77794 54484
rect 79070 54476 79670 54498
rect 79728 54476 80328 54498
rect 80386 54476 80986 54498
rect 81044 54476 81644 54498
rect 71356 53856 71956 53882
rect 72014 53856 72614 53882
rect 72672 53856 73272 53882
rect 73330 53856 73930 53882
rect 71416 53814 71840 53856
rect 72154 53814 72578 53856
rect 72736 53814 73160 53856
rect 73408 53814 73832 53856
rect 71356 53788 71956 53814
rect 72014 53788 72614 53814
rect 72672 53788 73272 53814
rect 73330 53788 73930 53814
rect 71356 53162 71956 53188
rect 72014 53162 72614 53188
rect 72672 53162 73272 53188
rect 73330 53162 73930 53188
rect 71410 53120 71834 53162
rect 72122 53120 72546 53162
rect 72732 53120 73156 53162
rect 73448 53120 73872 53162
rect 71356 53094 71956 53120
rect 72014 53094 72614 53120
rect 72672 53094 73272 53120
rect 73330 53094 73930 53120
rect 71356 52468 71956 52494
rect 72014 52468 72614 52494
rect 72672 52468 73272 52494
rect 73330 52468 73930 52494
rect 71396 52426 71820 52468
rect 72142 52426 72566 52468
rect 72770 52426 73194 52468
rect 73406 52426 73830 52468
rect 71356 52400 71956 52426
rect 72014 52400 72614 52426
rect 72672 52400 73272 52426
rect 73330 52400 73930 52426
rect 71356 51774 71956 51800
rect 72014 51774 72614 51800
rect 72672 51774 73272 51800
rect 73330 51774 73930 51800
rect 71392 51732 71816 51774
rect 72172 51732 72596 51774
rect 72722 51732 73146 51774
rect 73440 51732 73864 51774
rect 71356 51706 71956 51732
rect 72014 51706 72614 51732
rect 72672 51706 73272 51732
rect 73330 51706 73930 51732
rect 57526 51124 57614 51246
rect 45506 51066 45576 51124
rect 49500 51066 49570 51124
rect 53522 51066 53592 51124
rect 57544 51066 57614 51124
rect 42086 50466 42112 51066
rect 42712 50976 42738 51066
rect 42780 50976 42806 51066
rect 42712 50536 42806 50976
rect 42712 50466 42738 50536
rect 42780 50466 42806 50536
rect 43406 51000 43432 51066
rect 43474 51000 43500 51066
rect 43406 50560 43500 51000
rect 43406 50466 43432 50560
rect 43474 50466 43500 50560
rect 44100 50984 44126 51066
rect 44168 50984 44194 51066
rect 44100 50544 44194 50984
rect 44100 50466 44126 50544
rect 44168 50466 44194 50544
rect 44794 50996 44820 51066
rect 44862 50996 44888 51066
rect 44794 50556 44888 50996
rect 44794 50466 44820 50556
rect 44862 50466 44888 50556
rect 45488 50946 45576 51066
rect 46080 50946 46106 51066
rect 45488 50710 46106 50946
rect 45488 50466 45576 50710
rect 46080 50466 46106 50710
rect 46706 50976 46732 51066
rect 46774 50976 46800 51066
rect 46706 50536 46800 50976
rect 46706 50466 46732 50536
rect 46774 50466 46800 50536
rect 47400 51000 47426 51066
rect 47468 51000 47494 51066
rect 47400 50560 47494 51000
rect 47400 50466 47426 50560
rect 47468 50466 47494 50560
rect 48094 50984 48120 51066
rect 48162 50984 48188 51066
rect 48094 50544 48188 50984
rect 48094 50466 48120 50544
rect 48162 50466 48188 50544
rect 48788 50996 48814 51066
rect 48856 50996 48882 51066
rect 48788 50556 48882 50996
rect 48788 50466 48814 50556
rect 48856 50466 48882 50556
rect 49482 50906 49570 51066
rect 50102 50906 50128 51066
rect 49482 50670 50128 50906
rect 49482 50466 49570 50670
rect 50102 50466 50128 50670
rect 50728 50976 50754 51066
rect 50796 50976 50822 51066
rect 50728 50536 50822 50976
rect 50728 50466 50754 50536
rect 50796 50466 50822 50536
rect 51422 51000 51448 51066
rect 51490 51000 51516 51066
rect 51422 50560 51516 51000
rect 51422 50466 51448 50560
rect 51490 50466 51516 50560
rect 52116 50984 52142 51066
rect 52184 50984 52210 51066
rect 52116 50544 52210 50984
rect 52116 50466 52142 50544
rect 52184 50466 52210 50544
rect 52810 50996 52836 51066
rect 52878 50996 52904 51066
rect 52810 50556 52904 50996
rect 52810 50466 52836 50556
rect 52878 50466 52904 50556
rect 53504 50916 53592 51066
rect 54124 50916 54150 51066
rect 53504 50680 54150 50916
rect 53504 50466 53592 50680
rect 54124 50466 54150 50680
rect 54750 50976 54776 51066
rect 54818 50976 54844 51066
rect 54750 50536 54844 50976
rect 54750 50466 54776 50536
rect 54818 50466 54844 50536
rect 55444 51000 55470 51066
rect 55512 51000 55538 51066
rect 55444 50560 55538 51000
rect 55444 50466 55470 50560
rect 55512 50466 55538 50560
rect 56138 50984 56164 51066
rect 56206 50984 56232 51066
rect 56138 50544 56232 50984
rect 56138 50466 56164 50544
rect 56206 50466 56232 50544
rect 56832 50996 56858 51066
rect 56900 50996 56926 51066
rect 56832 50556 56926 50996
rect 56832 50466 56858 50556
rect 56900 50466 56926 50556
rect 57526 50466 57614 51066
rect 75220 53836 75820 53862
rect 75878 53836 76478 53862
rect 76536 53836 77136 53862
rect 77194 53836 77794 53862
rect 75280 53794 75704 53836
rect 76018 53794 76442 53836
rect 76600 53794 77024 53836
rect 77272 53794 77696 53836
rect 75220 53768 75820 53794
rect 75878 53768 76478 53794
rect 76536 53768 77136 53794
rect 77194 53768 77794 53794
rect 75220 53142 75820 53168
rect 75878 53142 76478 53168
rect 76536 53142 77136 53168
rect 77194 53142 77794 53168
rect 75274 53100 75698 53142
rect 75986 53100 76410 53142
rect 76596 53100 77020 53142
rect 77312 53100 77736 53142
rect 75220 53074 75820 53100
rect 75878 53074 76478 53100
rect 76536 53074 77136 53100
rect 77194 53074 77794 53100
rect 75220 52448 75820 52474
rect 75878 52448 76478 52474
rect 76536 52448 77136 52474
rect 77194 52448 77794 52474
rect 75260 52406 75684 52448
rect 76006 52406 76430 52448
rect 76634 52406 77058 52448
rect 77270 52406 77694 52448
rect 75220 52380 75820 52406
rect 75878 52380 76478 52406
rect 76536 52380 77136 52406
rect 77194 52380 77794 52406
rect 75220 51754 75820 51780
rect 75878 51754 76478 51780
rect 76536 51754 77136 51780
rect 77194 51754 77794 51780
rect 75256 51712 75680 51754
rect 76036 51712 76460 51754
rect 76586 51712 77010 51754
rect 77304 51712 77728 51754
rect 75220 51686 75820 51712
rect 75878 51686 76478 51712
rect 76536 51686 77136 51712
rect 77194 51686 77794 51712
rect 71356 51080 71956 51106
rect 72014 51080 72614 51106
rect 72672 51080 73272 51106
rect 73330 51080 73930 51106
rect 79070 53850 79670 53876
rect 79728 53850 80328 53876
rect 80386 53850 80986 53876
rect 81044 53850 81644 53876
rect 79130 53808 79554 53850
rect 79868 53808 80292 53850
rect 80450 53808 80874 53850
rect 81122 53808 81546 53850
rect 79070 53782 79670 53808
rect 79728 53782 80328 53808
rect 80386 53782 80986 53808
rect 81044 53782 81644 53808
rect 79070 53156 79670 53182
rect 79728 53156 80328 53182
rect 80386 53156 80986 53182
rect 81044 53156 81644 53182
rect 79124 53114 79548 53156
rect 79836 53114 80260 53156
rect 80446 53114 80870 53156
rect 81162 53114 81586 53156
rect 79070 53088 79670 53114
rect 79728 53088 80328 53114
rect 80386 53088 80986 53114
rect 81044 53088 81644 53114
rect 79070 52462 79670 52488
rect 79728 52462 80328 52488
rect 80386 52462 80986 52488
rect 81044 52462 81644 52488
rect 79110 52420 79534 52462
rect 79856 52420 80280 52462
rect 80484 52420 80908 52462
rect 81120 52420 81544 52462
rect 79070 52394 79670 52420
rect 79728 52394 80328 52420
rect 80386 52394 80986 52420
rect 81044 52394 81644 52420
rect 79070 51768 79670 51794
rect 79728 51768 80328 51794
rect 80386 51768 80986 51794
rect 81044 51768 81644 51794
rect 79106 51726 79530 51768
rect 79886 51726 80310 51768
rect 80436 51726 80860 51768
rect 81154 51726 81578 51768
rect 79070 51700 79670 51726
rect 79728 51700 80328 51726
rect 80386 51700 80986 51726
rect 81044 51700 81644 51726
rect 84891 54011 84991 54037
rect 85047 54011 85147 54037
rect 86161 54011 86261 54037
rect 83781 53984 83881 54010
rect 83937 53984 84037 54010
rect 84093 53984 84193 54010
rect 84249 53984 84349 54010
rect 84391 53984 84491 54010
rect 84563 53984 84663 54010
rect 83355 53955 83455 53981
rect 83511 53955 83611 53981
rect 83355 53641 83455 53805
rect 83511 53779 83611 53805
rect 83511 53757 83615 53779
rect 83511 53723 83536 53757
rect 83570 53723 83615 53757
rect 83511 53689 83615 53723
rect 83511 53655 83536 53689
rect 83570 53655 83615 53689
rect 83355 53621 83459 53641
rect 83511 53635 83615 53655
rect 83355 53587 83400 53621
rect 83434 53587 83459 53621
rect 83355 53553 83459 53587
rect 83355 53519 83400 53553
rect 83434 53519 83459 53553
rect 83355 53485 83459 53519
rect 83359 53459 83459 53485
rect 83515 53459 83615 53635
rect 83781 53730 83881 53900
rect 83937 53878 84037 53900
rect 83937 53778 84051 53878
rect 84093 53852 84193 53900
rect 84093 53818 84123 53852
rect 84157 53818 84193 53852
rect 84093 53802 84193 53818
rect 84249 53852 84349 53900
rect 84249 53818 84284 53852
rect 84318 53818 84349 53852
rect 84249 53802 84349 53818
rect 83781 53710 83909 53730
rect 83781 53676 83827 53710
rect 83861 53676 83909 53710
rect 83781 53642 83909 53676
rect 83781 53608 83827 53642
rect 83861 53608 83909 53642
rect 83781 53547 83909 53608
rect 83809 53525 83909 53547
rect 83951 53673 84051 53778
rect 84235 53760 84349 53802
rect 84391 53874 84491 53900
rect 84563 53874 84663 53900
rect 84391 53774 84510 53874
rect 83951 53639 83971 53673
rect 84005 53639 84051 53673
rect 83951 53605 84051 53639
rect 83951 53571 83971 53605
rect 84005 53571 84051 53605
rect 83951 53525 84051 53571
rect 84107 53725 84349 53760
rect 84405 53736 84510 53774
rect 84107 53683 84221 53725
rect 84405 53702 84456 53736
rect 84490 53702 84510 53736
rect 84107 53525 84207 53683
rect 84263 53667 84363 53683
rect 84263 53633 84283 53667
rect 84317 53633 84363 53667
rect 84263 53599 84363 53633
rect 84263 53565 84283 53599
rect 84317 53565 84363 53599
rect 84263 53525 84363 53565
rect 84405 53668 84510 53702
rect 84405 53634 84456 53668
rect 84490 53634 84510 53668
rect 84405 53547 84510 53634
rect 84552 53667 84663 53874
rect 85226 53895 85326 53921
rect 85368 53895 85468 53921
rect 85545 53895 85645 53921
rect 85701 53895 85801 53921
rect 85986 53861 86086 53887
rect 84552 53633 84609 53667
rect 84643 53633 84663 53667
rect 84891 53647 84991 53811
rect 85047 53785 85147 53811
rect 85047 53763 85138 53785
rect 85047 53729 85088 53763
rect 85122 53729 85138 53763
rect 85226 53755 85326 53811
rect 85047 53695 85138 53729
rect 85047 53661 85088 53695
rect 85122 53661 85138 53695
rect 84552 53613 84663 53633
rect 84405 53525 84505 53547
rect 84552 53525 84652 53613
rect 84824 53597 85005 53647
rect 85047 53641 85138 53661
rect 85180 53739 85326 53755
rect 85180 53705 85213 53739
rect 85247 53705 85326 53739
rect 85180 53685 85326 53705
rect 85368 53785 85468 53811
rect 85368 53685 85503 53785
rect 85180 53599 85223 53685
rect 85403 53664 85503 53685
rect 85403 53630 85449 53664
rect 85483 53630 85503 53664
rect 84824 53563 84844 53597
rect 84878 53563 85005 53597
rect 84824 53547 85005 53563
rect 84905 53525 85005 53547
rect 85061 53547 85223 53599
rect 85265 53603 85361 53623
rect 85265 53569 85281 53603
rect 85315 53569 85361 53603
rect 85061 53525 85161 53547
rect 85265 53535 85361 53569
rect 83809 53415 83909 53441
rect 83951 53415 84051 53441
rect 84107 53415 84207 53441
rect 84263 53415 84363 53441
rect 84405 53415 84505 53441
rect 84552 53415 84652 53441
rect 85265 53505 85281 53535
rect 85261 53501 85281 53505
rect 85315 53501 85361 53535
rect 85261 53459 85361 53501
rect 85403 53596 85503 53630
rect 85403 53562 85449 53596
rect 85483 53562 85503 53596
rect 85403 53459 85503 53562
rect 85545 53619 85645 53811
rect 85701 53739 85801 53811
rect 85701 53705 85721 53739
rect 85755 53705 85801 53739
rect 85701 53685 85801 53705
rect 85986 53685 86086 53711
rect 86161 53685 86261 53711
rect 85545 53599 85659 53619
rect 85545 53565 85579 53599
rect 85613 53565 85659 53599
rect 85545 53531 85659 53565
rect 85545 53497 85579 53531
rect 85613 53497 85659 53531
rect 85545 53481 85659 53497
rect 85559 53459 85659 53481
rect 85701 53585 86086 53685
rect 86146 53653 86261 53685
rect 86146 53619 86166 53653
rect 86200 53619 86261 53653
rect 86146 53585 86261 53619
rect 85701 53459 85801 53585
rect 85978 53559 86078 53585
rect 86157 53559 86257 53585
rect 85978 53449 86078 53475
rect 86157 53383 86257 53409
rect 83359 53349 83459 53375
rect 83515 53349 83615 53375
rect 84905 53349 85005 53375
rect 85061 53349 85161 53375
rect 85261 53349 85361 53375
rect 85403 53349 85503 53375
rect 85559 53349 85659 53375
rect 85701 53349 85801 53375
rect 75220 51060 75820 51086
rect 75878 51060 76478 51086
rect 76536 51060 77136 51086
rect 77194 51060 77794 51086
rect 79070 51074 79670 51100
rect 79728 51074 80328 51100
rect 80386 51074 80986 51100
rect 81044 51074 81644 51100
rect 77304 51022 77728 51060
rect 77304 50826 77348 51022
rect 77656 50826 77728 51022
rect 77304 50774 77728 50826
rect 45506 50408 45576 50466
rect 49500 50408 49570 50466
rect 53522 50408 53592 50466
rect 57544 50408 57614 50466
rect 42086 49808 42112 50408
rect 42712 50300 42738 50408
rect 42780 50300 42806 50408
rect 42712 49860 42806 50300
rect 42712 49808 42738 49860
rect 42780 49808 42806 49860
rect 43406 50312 43432 50408
rect 43474 50312 43500 50408
rect 43406 49872 43500 50312
rect 43406 49808 43432 49872
rect 43474 49808 43500 49872
rect 44100 50290 44126 50408
rect 44168 50290 44194 50408
rect 44100 49850 44194 50290
rect 44100 49808 44126 49850
rect 44168 49808 44194 49850
rect 44794 50262 44820 50408
rect 44862 50262 44888 50408
rect 44794 49822 44888 50262
rect 44794 49808 44820 49822
rect 44862 49808 44888 49822
rect 45488 50266 45576 50408
rect 46080 50266 46106 50408
rect 45488 50030 46106 50266
rect 45488 49808 45576 50030
rect 46080 49808 46106 50030
rect 46706 50300 46732 50408
rect 46774 50300 46800 50408
rect 46706 49860 46800 50300
rect 46706 49808 46732 49860
rect 46774 49808 46800 49860
rect 47400 50312 47426 50408
rect 47468 50312 47494 50408
rect 47400 49872 47494 50312
rect 47400 49808 47426 49872
rect 47468 49808 47494 49872
rect 48094 50290 48120 50408
rect 48162 50290 48188 50408
rect 48094 49850 48188 50290
rect 48094 49808 48120 49850
rect 48162 49808 48188 49850
rect 48788 50262 48814 50408
rect 48856 50262 48882 50408
rect 48788 49822 48882 50262
rect 48788 49808 48814 49822
rect 48856 49808 48882 49822
rect 49482 50214 49570 50408
rect 50102 50214 50128 50408
rect 49482 49978 50128 50214
rect 49482 49808 49570 49978
rect 50102 49808 50128 49978
rect 50728 50300 50754 50408
rect 50796 50300 50822 50408
rect 50728 49860 50822 50300
rect 50728 49808 50754 49860
rect 50796 49808 50822 49860
rect 51422 50312 51448 50408
rect 51490 50312 51516 50408
rect 51422 49872 51516 50312
rect 51422 49808 51448 49872
rect 51490 49808 51516 49872
rect 52116 50290 52142 50408
rect 52184 50290 52210 50408
rect 52116 49850 52210 50290
rect 52116 49808 52142 49850
rect 52184 49808 52210 49850
rect 52810 50262 52836 50408
rect 52878 50262 52904 50408
rect 52810 49822 52904 50262
rect 52810 49808 52836 49822
rect 52878 49808 52904 49822
rect 53504 50266 53592 50408
rect 54124 50266 54150 50408
rect 53504 50030 54150 50266
rect 53504 49808 53592 50030
rect 54124 49808 54150 50030
rect 54750 50300 54776 50408
rect 54818 50300 54844 50408
rect 54750 49860 54844 50300
rect 54750 49808 54776 49860
rect 54818 49808 54844 49860
rect 55444 50312 55470 50408
rect 55512 50312 55538 50408
rect 55444 49872 55538 50312
rect 55444 49808 55470 49872
rect 55512 49808 55538 49872
rect 56138 50290 56164 50408
rect 56206 50290 56232 50408
rect 56138 49850 56232 50290
rect 56138 49808 56164 49850
rect 56206 49808 56232 49850
rect 56832 50262 56858 50408
rect 56900 50262 56926 50408
rect 56832 49822 56926 50262
rect 56832 49808 56858 49822
rect 56900 49808 56926 49822
rect 57526 49808 57614 50408
rect 45506 49750 45576 49808
rect 49500 49750 49570 49808
rect 53522 49750 53592 49808
rect 57544 49750 57614 49808
rect 42086 49150 42112 49750
rect 42712 49668 42738 49750
rect 42780 49668 42806 49750
rect 42712 49228 42806 49668
rect 42712 49150 42738 49228
rect 42780 49150 42806 49228
rect 43406 49690 43432 49750
rect 43474 49690 43500 49750
rect 43406 49250 43500 49690
rect 43406 49150 43432 49250
rect 43474 49150 43500 49250
rect 44100 49690 44126 49750
rect 44168 49690 44194 49750
rect 44100 49250 44194 49690
rect 44100 49150 44126 49250
rect 44168 49150 44194 49250
rect 44794 49678 44820 49750
rect 44862 49678 44888 49750
rect 44794 49238 44888 49678
rect 44794 49150 44820 49238
rect 44862 49150 44888 49238
rect 45488 49572 45576 49750
rect 46080 49572 46106 49750
rect 45488 49336 46106 49572
rect 45488 49150 45576 49336
rect 46080 49150 46106 49336
rect 46706 49668 46732 49750
rect 46774 49668 46800 49750
rect 46706 49228 46800 49668
rect 46706 49150 46732 49228
rect 46774 49150 46800 49228
rect 47400 49690 47426 49750
rect 47468 49690 47494 49750
rect 47400 49250 47494 49690
rect 47400 49150 47426 49250
rect 47468 49150 47494 49250
rect 48094 49690 48120 49750
rect 48162 49690 48188 49750
rect 48094 49250 48188 49690
rect 48094 49150 48120 49250
rect 48162 49150 48188 49250
rect 48788 49678 48814 49750
rect 48856 49678 48882 49750
rect 48788 49238 48882 49678
rect 48788 49150 48814 49238
rect 48856 49150 48882 49238
rect 49482 49572 49570 49750
rect 50102 49572 50128 49750
rect 49482 49336 50128 49572
rect 49482 49150 49570 49336
rect 50102 49150 50128 49336
rect 50728 49668 50754 49750
rect 50796 49668 50822 49750
rect 50728 49228 50822 49668
rect 50728 49150 50754 49228
rect 50796 49150 50822 49228
rect 51422 49690 51448 49750
rect 51490 49690 51516 49750
rect 51422 49250 51516 49690
rect 51422 49150 51448 49250
rect 51490 49150 51516 49250
rect 52116 49690 52142 49750
rect 52184 49690 52210 49750
rect 52116 49250 52210 49690
rect 52116 49150 52142 49250
rect 52184 49150 52210 49250
rect 52810 49678 52836 49750
rect 52878 49678 52904 49750
rect 52810 49238 52904 49678
rect 52810 49150 52836 49238
rect 52878 49150 52904 49238
rect 53504 49678 53592 49750
rect 54124 49678 54150 49750
rect 53504 49442 54150 49678
rect 53504 49150 53592 49442
rect 54124 49150 54150 49442
rect 54750 49668 54776 49750
rect 54818 49668 54844 49750
rect 54750 49228 54844 49668
rect 54750 49150 54776 49228
rect 54818 49150 54844 49228
rect 55444 49690 55470 49750
rect 55512 49690 55538 49750
rect 55444 49250 55538 49690
rect 55444 49150 55470 49250
rect 55512 49150 55538 49250
rect 56138 49690 56164 49750
rect 56206 49690 56232 49750
rect 56138 49250 56232 49690
rect 56138 49150 56164 49250
rect 56206 49150 56232 49250
rect 56832 49678 56858 49750
rect 56900 49678 56926 49750
rect 56832 49238 56926 49678
rect 56832 49150 56858 49238
rect 56900 49150 56926 49238
rect 57526 49150 57614 49750
rect 45506 49092 45576 49150
rect 49500 49092 49570 49150
rect 53522 49092 53592 49150
rect 57544 49092 57614 49150
rect 42086 48492 42112 49092
rect 42712 48960 42738 49092
rect 42780 48960 42806 49092
rect 42712 48520 42806 48960
rect 42712 48492 42738 48520
rect 42780 48492 42806 48520
rect 43406 49002 43432 49092
rect 43474 49002 43500 49092
rect 43406 48562 43500 49002
rect 43406 48492 43432 48562
rect 43474 48492 43500 48562
rect 44100 49014 44126 49092
rect 44168 49014 44194 49092
rect 44100 48574 44194 49014
rect 44100 48492 44126 48574
rect 44168 48492 44194 48574
rect 44794 49040 44820 49092
rect 44862 49040 44888 49092
rect 44794 48600 44888 49040
rect 44794 48492 44820 48600
rect 44862 48492 44888 48600
rect 45488 49062 45576 49092
rect 46080 49062 46106 49092
rect 45488 48826 46106 49062
rect 45488 48812 45576 48826
rect 45488 48492 45514 48812
rect 46080 48492 46106 48826
rect 46706 48960 46732 49092
rect 46774 48960 46800 49092
rect 46706 48520 46800 48960
rect 46706 48492 46732 48520
rect 46774 48492 46800 48520
rect 47400 49002 47426 49092
rect 47468 49002 47494 49092
rect 47400 48562 47494 49002
rect 47400 48492 47426 48562
rect 47468 48492 47494 48562
rect 48094 49014 48120 49092
rect 48162 49014 48188 49092
rect 48094 48574 48188 49014
rect 48094 48492 48120 48574
rect 48162 48492 48188 48574
rect 48788 49040 48814 49092
rect 48856 49040 48882 49092
rect 48788 48600 48882 49040
rect 48788 48492 48814 48600
rect 48856 48492 48882 48600
rect 49482 49046 49570 49092
rect 50102 49046 50128 49092
rect 49482 48810 50128 49046
rect 49482 48492 49508 48810
rect 50102 48492 50128 48810
rect 50728 48960 50754 49092
rect 50796 48960 50822 49092
rect 50728 48520 50822 48960
rect 50728 48492 50754 48520
rect 50796 48492 50822 48520
rect 51422 49002 51448 49092
rect 51490 49002 51516 49092
rect 51422 48562 51516 49002
rect 51422 48492 51448 48562
rect 51490 48492 51516 48562
rect 52116 49014 52142 49092
rect 52184 49014 52210 49092
rect 52116 48574 52210 49014
rect 52116 48492 52142 48574
rect 52184 48492 52210 48574
rect 52810 49040 52836 49092
rect 52878 49040 52904 49092
rect 52810 48600 52904 49040
rect 52810 48492 52836 48600
rect 52878 48492 52904 48600
rect 53504 49076 53592 49092
rect 54124 49076 54150 49092
rect 53504 48840 54150 49076
rect 53504 48812 53592 48840
rect 53504 48492 53530 48812
rect 54124 48492 54150 48840
rect 54750 48960 54776 49092
rect 54818 48960 54844 49092
rect 54750 48520 54844 48960
rect 54750 48492 54776 48520
rect 54818 48492 54844 48520
rect 55444 49002 55470 49092
rect 55512 49002 55538 49092
rect 55444 48562 55538 49002
rect 55444 48492 55470 48562
rect 55512 48492 55538 48562
rect 56138 49014 56164 49092
rect 56206 49014 56232 49092
rect 56138 48574 56232 49014
rect 56138 48492 56164 48574
rect 56206 48492 56232 48574
rect 56832 49040 56858 49092
rect 56900 49040 56926 49092
rect 56832 48600 56926 49040
rect 56832 48492 56858 48600
rect 56900 48492 56926 48600
rect 57526 48812 57614 49092
rect 57526 48492 57552 48812
rect 30102 43998 31230 44070
rect 23908 43890 37838 43998
rect 42918 43936 56848 44042
rect 23908 43868 38042 43890
rect 42918 43878 49550 43936
rect 6158 43736 16898 43822
rect 6158 43698 11050 43736
rect 5524 43606 11050 43698
rect 11240 43698 16898 43736
rect 23476 43702 38042 43868
rect 11240 43606 17462 43698
rect 5524 43600 17462 43606
rect 5524 43474 6560 43600
rect 10630 43482 11666 43600
rect 16426 43490 17462 43600
rect 2454 43432 7080 43474
rect 8968 43440 13594 43482
rect 15474 43448 20100 43490
rect 23476 43474 24556 43702
rect 30106 43490 31186 43702
rect 36962 43496 38042 43702
rect 42490 43746 49550 43878
rect 42490 43496 43570 43746
rect 49214 43672 49550 43746
rect 49974 43922 56848 43936
rect 49974 43746 57470 43922
rect 49974 43672 50294 43746
rect 49214 43518 50294 43672
rect 56390 43532 57470 43746
rect 15024 43442 20256 43448
rect 8518 43434 13750 43440
rect 2004 43426 7236 43432
rect 2004 43406 3004 43426
rect 3062 43406 4062 43426
rect 4120 43406 5120 43426
rect 5178 43406 6178 43426
rect 6236 43406 7236 43426
rect 8518 43414 9518 43434
rect 9576 43414 10576 43434
rect 10634 43414 11634 43434
rect 11692 43414 12692 43434
rect 12750 43414 13750 43434
rect 15024 43422 16024 43442
rect 16082 43422 17082 43442
rect 17140 43422 18140 43442
rect 18198 43422 19198 43442
rect 19256 43422 20256 43442
rect 21964 43432 26590 43474
rect 28486 43448 33112 43490
rect 34996 43454 39622 43496
rect 41486 43454 46112 43496
rect 48074 43476 52700 43518
rect 54588 43490 59214 43532
rect 54138 43484 59370 43490
rect 47624 43470 52856 43476
rect 34546 43448 39778 43454
rect 28036 43442 33268 43448
rect 21514 43426 26746 43432
rect 21514 43406 22514 43426
rect 22572 43406 23572 43426
rect 23630 43406 24630 43426
rect 24688 43406 25688 43426
rect 25746 43406 26746 43426
rect 28036 43422 29036 43442
rect 29094 43422 30094 43442
rect 30152 43422 31152 43442
rect 31210 43422 32210 43442
rect 32268 43422 33268 43442
rect 34546 43428 35546 43448
rect 35604 43428 36604 43448
rect 36662 43428 37662 43448
rect 37720 43428 38720 43448
rect 38778 43428 39778 43448
rect 41036 43448 46268 43454
rect 47624 43450 48624 43470
rect 48682 43450 49682 43470
rect 49740 43450 50740 43470
rect 50798 43450 51798 43470
rect 51856 43450 52856 43470
rect 54138 43464 55138 43484
rect 55196 43464 56196 43484
rect 56254 43464 57254 43484
rect 57312 43464 58312 43484
rect 58370 43464 59370 43484
rect 41036 43428 42036 43448
rect 42094 43428 43094 43448
rect 43152 43428 44152 43448
rect 44210 43428 45210 43448
rect 45268 43428 46268 43448
rect 2004 42380 3004 42406
rect 3062 42380 4062 42406
rect 4120 42380 5120 42406
rect 5178 42380 6178 42406
rect 6236 42380 7236 42406
rect 8518 42388 9518 42414
rect 9576 42388 10576 42414
rect 10634 42388 11634 42414
rect 11692 42388 12692 42414
rect 12750 42388 13750 42414
rect 15024 42396 16024 42422
rect 16082 42396 17082 42422
rect 17140 42396 18140 42422
rect 18198 42396 19198 42422
rect 19256 42396 20256 42422
rect 2256 42338 2790 42380
rect 3294 42338 3828 42380
rect 4412 42338 4946 42380
rect 5428 42338 5962 42380
rect 6494 42338 7028 42380
rect 8770 42346 9304 42388
rect 9808 42346 10342 42388
rect 10926 42346 11460 42388
rect 11942 42346 12476 42388
rect 13008 42346 13542 42388
rect 15276 42354 15810 42396
rect 16314 42354 16848 42396
rect 17432 42354 17966 42396
rect 18448 42354 18982 42396
rect 19514 42354 20048 42396
rect 21514 42380 22514 42406
rect 22572 42380 23572 42406
rect 23630 42380 24630 42406
rect 24688 42380 25688 42406
rect 25746 42380 26746 42406
rect 28036 42396 29036 42422
rect 29094 42396 30094 42422
rect 30152 42396 31152 42422
rect 31210 42396 32210 42422
rect 32268 42396 33268 42422
rect 34546 42402 35546 42428
rect 35604 42402 36604 42428
rect 36662 42402 37662 42428
rect 37720 42402 38720 42428
rect 38778 42402 39778 42428
rect 41036 42402 42036 42428
rect 42094 42402 43094 42428
rect 43152 42402 44152 42428
rect 44210 42402 45210 42428
rect 45268 42402 46268 42428
rect 47624 42424 48624 42450
rect 48682 42424 49682 42450
rect 49740 42424 50740 42450
rect 50798 42424 51798 42450
rect 51856 42424 52856 42450
rect 54138 42438 55138 42464
rect 55196 42438 56196 42464
rect 56254 42438 57254 42464
rect 57312 42438 58312 42464
rect 58370 42438 59370 42464
rect 2004 42312 3004 42338
rect 3062 42312 4062 42338
rect 4120 42312 5120 42338
rect 5178 42312 6178 42338
rect 6236 42312 7236 42338
rect 8518 42320 9518 42346
rect 9576 42320 10576 42346
rect 10634 42320 11634 42346
rect 11692 42320 12692 42346
rect 12750 42320 13750 42346
rect 15024 42328 16024 42354
rect 16082 42328 17082 42354
rect 17140 42328 18140 42354
rect 18198 42328 19198 42354
rect 19256 42328 20256 42354
rect 21766 42338 22300 42380
rect 22804 42338 23338 42380
rect 23922 42338 24456 42380
rect 24938 42338 25472 42380
rect 26004 42338 26538 42380
rect 28288 42354 28822 42396
rect 29326 42354 29860 42396
rect 30444 42354 30978 42396
rect 31460 42354 31994 42396
rect 32526 42354 33060 42396
rect 34798 42360 35332 42402
rect 35836 42360 36370 42402
rect 36954 42360 37488 42402
rect 37970 42360 38504 42402
rect 39036 42360 39570 42402
rect 41288 42360 41822 42402
rect 42326 42360 42860 42402
rect 43444 42360 43978 42402
rect 44460 42360 44994 42402
rect 45526 42360 46060 42402
rect 47876 42382 48410 42424
rect 48914 42382 49448 42424
rect 50032 42382 50566 42424
rect 51048 42382 51582 42424
rect 52114 42382 52648 42424
rect 54390 42396 54924 42438
rect 55428 42396 55962 42438
rect 56546 42396 57080 42438
rect 57562 42396 58096 42438
rect 58628 42396 59162 42438
rect 2004 41286 3004 41312
rect 3062 41286 4062 41312
rect 4120 41286 5120 41312
rect 5178 41286 6178 41312
rect 6236 41286 7236 41312
rect 2292 41244 2826 41286
rect 3248 41244 3782 41286
rect 4356 41244 4890 41286
rect 5462 41244 5996 41286
rect 6492 41244 7026 41286
rect 2004 41218 3004 41244
rect 3062 41218 4062 41244
rect 4120 41218 5120 41244
rect 5178 41218 6178 41244
rect 6236 41218 7236 41244
rect 8518 41294 9518 41320
rect 9576 41294 10576 41320
rect 10634 41294 11634 41320
rect 11692 41294 12692 41320
rect 12750 41294 13750 41320
rect 8806 41252 9340 41294
rect 9762 41252 10296 41294
rect 10870 41252 11404 41294
rect 11976 41252 12510 41294
rect 13006 41252 13540 41294
rect 8518 41226 9518 41252
rect 9576 41226 10576 41252
rect 10634 41226 11634 41252
rect 11692 41226 12692 41252
rect 12750 41226 13750 41252
rect 2004 40192 3004 40218
rect 3062 40192 4062 40218
rect 4120 40192 5120 40218
rect 5178 40192 6178 40218
rect 6236 40192 7236 40218
rect 2228 40150 2762 40192
rect 3282 40150 3816 40192
rect 4334 40150 4868 40192
rect 5442 40150 5976 40192
rect 6498 40150 7032 40192
rect 2004 40124 3004 40150
rect 3062 40124 4062 40150
rect 4120 40124 5120 40150
rect 5178 40124 6178 40150
rect 6236 40124 7236 40150
rect 21514 42312 22514 42338
rect 22572 42312 23572 42338
rect 23630 42312 24630 42338
rect 24688 42312 25688 42338
rect 25746 42312 26746 42338
rect 28036 42328 29036 42354
rect 29094 42328 30094 42354
rect 30152 42328 31152 42354
rect 31210 42328 32210 42354
rect 32268 42328 33268 42354
rect 34546 42334 35546 42360
rect 35604 42334 36604 42360
rect 36662 42334 37662 42360
rect 37720 42334 38720 42360
rect 38778 42334 39778 42360
rect 41036 42334 42036 42360
rect 42094 42334 43094 42360
rect 43152 42334 44152 42360
rect 44210 42334 45210 42360
rect 45268 42334 46268 42360
rect 47624 42356 48624 42382
rect 48682 42356 49682 42382
rect 49740 42356 50740 42382
rect 50798 42356 51798 42382
rect 51856 42356 52856 42382
rect 54138 42370 55138 42396
rect 55196 42370 56196 42396
rect 56254 42370 57254 42396
rect 57312 42370 58312 42396
rect 58370 42370 59370 42396
rect 15024 41302 16024 41328
rect 16082 41302 17082 41328
rect 17140 41302 18140 41328
rect 18198 41302 19198 41328
rect 19256 41302 20256 41328
rect 15312 41260 15846 41302
rect 16268 41260 16802 41302
rect 17376 41260 17910 41302
rect 18482 41260 19016 41302
rect 19512 41260 20046 41302
rect 15024 41234 16024 41260
rect 16082 41234 17082 41260
rect 17140 41234 18140 41260
rect 18198 41234 19198 41260
rect 19256 41234 20256 41260
rect 8518 40200 9518 40226
rect 9576 40200 10576 40226
rect 10634 40200 11634 40226
rect 11692 40200 12692 40226
rect 12750 40200 13750 40226
rect 8742 40158 9276 40200
rect 9796 40158 10330 40200
rect 10848 40158 11382 40200
rect 11956 40158 12490 40200
rect 13012 40158 13546 40200
rect 8518 40132 9518 40158
rect 9576 40132 10576 40158
rect 10634 40132 11634 40158
rect 11692 40132 12692 40158
rect 12750 40132 13750 40158
rect 21514 41286 22514 41312
rect 22572 41286 23572 41312
rect 23630 41286 24630 41312
rect 24688 41286 25688 41312
rect 25746 41286 26746 41312
rect 21802 41244 22336 41286
rect 22758 41244 23292 41286
rect 23866 41244 24400 41286
rect 24972 41244 25506 41286
rect 26002 41244 26536 41286
rect 21514 41218 22514 41244
rect 22572 41218 23572 41244
rect 23630 41218 24630 41244
rect 24688 41218 25688 41244
rect 25746 41218 26746 41244
rect 15024 40208 16024 40234
rect 16082 40208 17082 40234
rect 17140 40208 18140 40234
rect 18198 40208 19198 40234
rect 19256 40208 20256 40234
rect 15248 40166 15782 40208
rect 16302 40166 16836 40208
rect 17354 40166 17888 40208
rect 18462 40166 18996 40208
rect 19518 40166 20052 40208
rect 15024 40140 16024 40166
rect 16082 40140 17082 40166
rect 17140 40140 18140 40166
rect 18198 40140 19198 40166
rect 19256 40140 20256 40166
rect 28036 41302 29036 41328
rect 29094 41302 30094 41328
rect 30152 41302 31152 41328
rect 31210 41302 32210 41328
rect 32268 41302 33268 41328
rect 28324 41260 28858 41302
rect 29280 41260 29814 41302
rect 30388 41260 30922 41302
rect 31494 41260 32028 41302
rect 32524 41260 33058 41302
rect 28036 41234 29036 41260
rect 29094 41234 30094 41260
rect 30152 41234 31152 41260
rect 31210 41234 32210 41260
rect 32268 41234 33268 41260
rect 21514 40192 22514 40218
rect 22572 40192 23572 40218
rect 23630 40192 24630 40218
rect 24688 40192 25688 40218
rect 25746 40192 26746 40218
rect 21738 40150 22272 40192
rect 22792 40150 23326 40192
rect 23844 40150 24378 40192
rect 24952 40150 25486 40192
rect 26008 40150 26542 40192
rect 21514 40124 22514 40150
rect 22572 40124 23572 40150
rect 23630 40124 24630 40150
rect 24688 40124 25688 40150
rect 25746 40124 26746 40150
rect 2004 39098 3004 39124
rect 3062 39098 4062 39124
rect 4120 39098 5120 39124
rect 5178 39098 6178 39124
rect 6236 39098 7236 39124
rect 8518 39106 9518 39132
rect 9576 39106 10576 39132
rect 10634 39106 11634 39132
rect 11692 39106 12692 39132
rect 12750 39106 13750 39132
rect 15024 39114 16024 39140
rect 16082 39114 17082 39140
rect 17140 39114 18140 39140
rect 18198 39114 19198 39140
rect 19256 39114 20256 39140
rect 34546 41308 35546 41334
rect 35604 41308 36604 41334
rect 36662 41308 37662 41334
rect 37720 41308 38720 41334
rect 38778 41308 39778 41334
rect 34834 41266 35368 41308
rect 35790 41266 36324 41308
rect 36898 41266 37432 41308
rect 38004 41266 38538 41308
rect 39034 41266 39568 41308
rect 34546 41240 35546 41266
rect 35604 41240 36604 41266
rect 36662 41240 37662 41266
rect 37720 41240 38720 41266
rect 38778 41240 39778 41266
rect 28036 40208 29036 40234
rect 29094 40208 30094 40234
rect 30152 40208 31152 40234
rect 31210 40208 32210 40234
rect 32268 40208 33268 40234
rect 28260 40166 28794 40208
rect 29314 40166 29848 40208
rect 30366 40166 30900 40208
rect 31474 40166 32008 40208
rect 32530 40166 33064 40208
rect 28036 40140 29036 40166
rect 29094 40140 30094 40166
rect 30152 40140 31152 40166
rect 31210 40140 32210 40166
rect 32268 40140 33268 40166
rect 41036 41308 42036 41334
rect 42094 41308 43094 41334
rect 43152 41308 44152 41334
rect 44210 41308 45210 41334
rect 45268 41308 46268 41334
rect 41324 41266 41858 41308
rect 42280 41266 42814 41308
rect 43388 41266 43922 41308
rect 44494 41266 45028 41308
rect 45524 41266 46058 41308
rect 41036 41240 42036 41266
rect 42094 41240 43094 41266
rect 43152 41240 44152 41266
rect 44210 41240 45210 41266
rect 45268 41240 46268 41266
rect 34546 40214 35546 40240
rect 35604 40214 36604 40240
rect 36662 40214 37662 40240
rect 37720 40214 38720 40240
rect 38778 40214 39778 40240
rect 34770 40172 35304 40214
rect 35824 40172 36358 40214
rect 36876 40172 37410 40214
rect 37984 40172 38518 40214
rect 39040 40172 39574 40214
rect 34546 40146 35546 40172
rect 35604 40146 36604 40172
rect 36662 40146 37662 40172
rect 37720 40146 38720 40172
rect 38778 40146 39778 40172
rect 47624 41330 48624 41356
rect 48682 41330 49682 41356
rect 49740 41330 50740 41356
rect 50798 41330 51798 41356
rect 51856 41330 52856 41356
rect 47912 41288 48446 41330
rect 48868 41288 49402 41330
rect 49976 41288 50510 41330
rect 51082 41288 51616 41330
rect 52112 41288 52646 41330
rect 47624 41262 48624 41288
rect 48682 41262 49682 41288
rect 49740 41262 50740 41288
rect 50798 41262 51798 41288
rect 51856 41262 52856 41288
rect 41036 40214 42036 40240
rect 42094 40214 43094 40240
rect 43152 40214 44152 40240
rect 44210 40214 45210 40240
rect 45268 40214 46268 40240
rect 41260 40172 41794 40214
rect 42314 40172 42848 40214
rect 43366 40172 43900 40214
rect 44474 40172 45008 40214
rect 45530 40172 46064 40214
rect 41036 40146 42036 40172
rect 42094 40146 43094 40172
rect 43152 40146 44152 40172
rect 44210 40146 45210 40172
rect 45268 40146 46268 40172
rect 54138 41344 55138 41370
rect 55196 41344 56196 41370
rect 56254 41344 57254 41370
rect 57312 41344 58312 41370
rect 58370 41344 59370 41370
rect 54426 41302 54960 41344
rect 55382 41302 55916 41344
rect 56490 41302 57024 41344
rect 57596 41302 58130 41344
rect 58626 41302 59160 41344
rect 54138 41276 55138 41302
rect 55196 41276 56196 41302
rect 56254 41276 57254 41302
rect 57312 41276 58312 41302
rect 58370 41276 59370 41302
rect 47624 40236 48624 40262
rect 48682 40236 49682 40262
rect 49740 40236 50740 40262
rect 50798 40236 51798 40262
rect 51856 40236 52856 40262
rect 47848 40194 48382 40236
rect 48902 40194 49436 40236
rect 49954 40194 50488 40236
rect 51062 40194 51596 40236
rect 52118 40194 52652 40236
rect 47624 40168 48624 40194
rect 48682 40168 49682 40194
rect 49740 40168 50740 40194
rect 50798 40168 51798 40194
rect 51856 40168 52856 40194
rect 54138 40250 55138 40276
rect 55196 40250 56196 40276
rect 56254 40250 57254 40276
rect 57312 40250 58312 40276
rect 58370 40250 59370 40276
rect 54362 40208 54896 40250
rect 55416 40208 55950 40250
rect 56468 40208 57002 40250
rect 57576 40208 58110 40250
rect 58632 40208 59166 40250
rect 54138 40182 55138 40208
rect 55196 40182 56196 40208
rect 56254 40182 57254 40208
rect 57312 40182 58312 40208
rect 58370 40182 59370 40208
rect 2256 39056 2790 39098
rect 3354 39056 3888 39098
rect 4382 39056 4916 39098
rect 5346 39056 5880 39098
rect 6446 39056 6980 39098
rect 8770 39064 9304 39106
rect 9868 39064 10402 39106
rect 10896 39064 11430 39106
rect 11860 39064 12394 39106
rect 12960 39064 13494 39106
rect 15276 39072 15810 39114
rect 16374 39072 16908 39114
rect 17402 39072 17936 39114
rect 18366 39072 18900 39114
rect 19466 39072 20000 39114
rect 21514 39098 22514 39124
rect 22572 39098 23572 39124
rect 23630 39098 24630 39124
rect 24688 39098 25688 39124
rect 25746 39098 26746 39124
rect 28036 39114 29036 39140
rect 29094 39114 30094 39140
rect 30152 39114 31152 39140
rect 31210 39114 32210 39140
rect 32268 39114 33268 39140
rect 34546 39120 35546 39146
rect 35604 39120 36604 39146
rect 36662 39120 37662 39146
rect 37720 39120 38720 39146
rect 38778 39120 39778 39146
rect 41036 39120 42036 39146
rect 42094 39120 43094 39146
rect 43152 39120 44152 39146
rect 44210 39120 45210 39146
rect 45268 39120 46268 39146
rect 47624 39142 48624 39168
rect 48682 39142 49682 39168
rect 49740 39142 50740 39168
rect 50798 39142 51798 39168
rect 51856 39142 52856 39168
rect 54138 39156 55138 39182
rect 55196 39156 56196 39182
rect 56254 39156 57254 39182
rect 57312 39156 58312 39182
rect 58370 39156 59370 39182
rect 2004 39030 3004 39056
rect 3062 39030 4062 39056
rect 4120 39030 5120 39056
rect 5178 39030 6178 39056
rect 6236 39030 7236 39056
rect 8518 39038 9518 39064
rect 9576 39038 10576 39064
rect 10634 39038 11634 39064
rect 11692 39038 12692 39064
rect 12750 39038 13750 39064
rect 15024 39046 16024 39072
rect 16082 39046 17082 39072
rect 17140 39046 18140 39072
rect 18198 39046 19198 39072
rect 19256 39046 20256 39072
rect 21766 39056 22300 39098
rect 22864 39056 23398 39098
rect 23892 39056 24426 39098
rect 24856 39056 25390 39098
rect 25956 39056 26490 39098
rect 28288 39072 28822 39114
rect 29386 39072 29920 39114
rect 30414 39072 30948 39114
rect 31378 39072 31912 39114
rect 32478 39072 33012 39114
rect 34798 39078 35332 39120
rect 35896 39078 36430 39120
rect 36924 39078 37458 39120
rect 37888 39078 38422 39120
rect 38988 39078 39522 39120
rect 41288 39078 41822 39120
rect 42386 39078 42920 39120
rect 43414 39078 43948 39120
rect 44378 39078 44912 39120
rect 45478 39078 46012 39120
rect 47876 39100 48410 39142
rect 48974 39100 49508 39142
rect 50002 39100 50536 39142
rect 50966 39100 51500 39142
rect 52066 39100 52600 39142
rect 54390 39114 54924 39156
rect 55488 39114 56022 39156
rect 56516 39114 57050 39156
rect 57480 39114 58014 39156
rect 58580 39114 59114 39156
rect 21514 39030 22514 39056
rect 22572 39030 23572 39056
rect 23630 39030 24630 39056
rect 24688 39030 25688 39056
rect 25746 39030 26746 39056
rect 28036 39046 29036 39072
rect 29094 39046 30094 39072
rect 30152 39046 31152 39072
rect 31210 39046 32210 39072
rect 32268 39046 33268 39072
rect 34546 39052 35546 39078
rect 35604 39052 36604 39078
rect 36662 39052 37662 39078
rect 37720 39052 38720 39078
rect 38778 39052 39778 39078
rect 41036 39052 42036 39078
rect 42094 39052 43094 39078
rect 43152 39052 44152 39078
rect 44210 39052 45210 39078
rect 45268 39052 46268 39078
rect 47624 39074 48624 39100
rect 48682 39074 49682 39100
rect 49740 39074 50740 39100
rect 50798 39074 51798 39100
rect 51856 39074 52856 39100
rect 54138 39088 55138 39114
rect 55196 39088 56196 39114
rect 56254 39088 57254 39114
rect 57312 39088 58312 39114
rect 58370 39088 59370 39114
rect 2004 38004 3004 38030
rect 3062 38004 4062 38030
rect 4120 38004 5120 38030
rect 5178 38004 6178 38030
rect 6236 38004 7236 38030
rect 8518 38018 9518 38038
rect 9576 38018 10576 38038
rect 10634 38018 11634 38038
rect 11692 38018 12692 38038
rect 12750 38018 13750 38038
rect 15024 38026 16024 38046
rect 16082 38026 17082 38046
rect 17140 38026 18140 38046
rect 18198 38026 19198 38046
rect 19256 38026 20256 38046
rect 47624 38056 48624 38074
rect 48682 38056 49682 38074
rect 49740 38056 50740 38074
rect 50798 38056 51798 38074
rect 51856 38056 52856 38074
rect 54138 38068 55138 38088
rect 55196 38068 56196 38088
rect 56254 38068 57254 38088
rect 57312 38068 58312 38088
rect 58370 38068 59370 38088
rect 54138 38062 59370 38068
rect 15024 38020 20256 38026
rect 8518 38012 13750 38018
rect 2488 37658 2654 38004
rect 3382 37658 3548 38004
rect 4412 37658 4578 38004
rect 5446 37658 5612 38004
rect 6480 37658 6646 38004
rect 8934 37954 13584 38012
rect 11152 37666 11480 37954
rect 15458 37924 19714 38020
rect 21514 38014 22514 38030
rect 22572 38014 23572 38030
rect 23630 38014 24630 38030
rect 24688 38014 25688 38030
rect 25746 38014 26746 38030
rect 28036 38028 29036 38046
rect 29094 38028 30094 38046
rect 30152 38028 31152 38046
rect 31210 38028 32210 38046
rect 32268 38028 33268 38046
rect 28036 38020 33268 38028
rect 34546 38036 35546 38052
rect 35604 38036 36604 38052
rect 36662 38036 37662 38052
rect 37720 38036 38720 38052
rect 38778 38036 39778 38052
rect 34546 38026 39778 38036
rect 41036 38034 42036 38052
rect 42094 38034 43094 38052
rect 43152 38034 44152 38052
rect 44210 38034 45210 38052
rect 45268 38034 46268 38052
rect 47624 38048 52856 38056
rect 41036 38026 46268 38034
rect 21514 38004 26746 38014
rect 18282 37674 18438 37924
rect 22014 37826 26492 38004
rect 2454 37616 7080 37658
rect 8968 37624 13594 37666
rect 15474 37632 20100 37674
rect 23596 37658 23894 37826
rect 28532 37810 32830 38020
rect 35016 37832 39506 38026
rect 41484 37834 45974 38026
rect 30074 37674 30372 37810
rect 36470 37680 36768 37832
rect 43026 37680 43324 37834
rect 48104 37782 52562 38048
rect 54564 37904 59158 38062
rect 50478 37702 50776 37782
rect 55740 37716 55966 37904
rect 15024 37626 20256 37632
rect 8518 37618 13750 37624
rect 2004 37610 7236 37616
rect 2004 37590 3004 37610
rect 3062 37590 4062 37610
rect 4120 37590 5120 37610
rect 5178 37590 6178 37610
rect 6236 37590 7236 37610
rect 8518 37598 9518 37618
rect 9576 37598 10576 37618
rect 10634 37598 11634 37618
rect 11692 37598 12692 37618
rect 12750 37598 13750 37618
rect 15024 37606 16024 37626
rect 16082 37606 17082 37626
rect 17140 37606 18140 37626
rect 18198 37606 19198 37626
rect 19256 37606 20256 37626
rect 21964 37616 26590 37658
rect 28486 37632 33112 37674
rect 34996 37638 39622 37680
rect 41486 37638 46112 37680
rect 48074 37660 52700 37702
rect 54588 37674 59214 37716
rect 54138 37668 59370 37674
rect 47624 37654 52856 37660
rect 34546 37632 39778 37638
rect 28036 37626 33268 37632
rect 21514 37610 26746 37616
rect 21514 37590 22514 37610
rect 22572 37590 23572 37610
rect 23630 37590 24630 37610
rect 24688 37590 25688 37610
rect 25746 37590 26746 37610
rect 28036 37606 29036 37626
rect 29094 37606 30094 37626
rect 30152 37606 31152 37626
rect 31210 37606 32210 37626
rect 32268 37606 33268 37626
rect 34546 37612 35546 37632
rect 35604 37612 36604 37632
rect 36662 37612 37662 37632
rect 37720 37612 38720 37632
rect 38778 37612 39778 37632
rect 41036 37632 46268 37638
rect 47624 37634 48624 37654
rect 48682 37634 49682 37654
rect 49740 37634 50740 37654
rect 50798 37634 51798 37654
rect 51856 37634 52856 37654
rect 54138 37648 55138 37668
rect 55196 37648 56196 37668
rect 56254 37648 57254 37668
rect 57312 37648 58312 37668
rect 58370 37648 59370 37668
rect 41036 37612 42036 37632
rect 42094 37628 44152 37632
rect 42094 37612 43094 37628
rect 43152 37612 44152 37628
rect 44210 37612 45210 37632
rect 45268 37612 46268 37632
rect 2004 36564 3004 36590
rect 3062 36564 4062 36590
rect 4120 36564 5120 36590
rect 5178 36564 6178 36590
rect 6236 36564 7236 36590
rect 8518 36572 9518 36598
rect 9576 36572 10576 36598
rect 10634 36572 11634 36598
rect 11692 36572 12692 36598
rect 12750 36572 13750 36598
rect 15024 36580 16024 36606
rect 16082 36580 17082 36606
rect 17140 36580 18140 36606
rect 18198 36580 19198 36606
rect 19256 36580 20256 36606
rect 2256 36522 2790 36564
rect 3294 36522 3828 36564
rect 4412 36522 4946 36564
rect 5428 36522 5962 36564
rect 6494 36522 7028 36564
rect 8770 36530 9304 36572
rect 9808 36530 10342 36572
rect 10926 36530 11460 36572
rect 11942 36530 12476 36572
rect 13008 36530 13542 36572
rect 15276 36538 15810 36580
rect 16314 36538 16848 36580
rect 17432 36538 17966 36580
rect 18448 36538 18982 36580
rect 19514 36538 20048 36580
rect 21514 36564 22514 36590
rect 22572 36564 23572 36590
rect 23630 36564 24630 36590
rect 24688 36564 25688 36590
rect 25746 36564 26746 36590
rect 28036 36580 29036 36606
rect 29094 36580 30094 36606
rect 30152 36580 31152 36606
rect 31210 36580 32210 36606
rect 32268 36580 33268 36606
rect 34546 36586 35546 36612
rect 35604 36586 36604 36612
rect 36662 36586 37662 36612
rect 37720 36586 38720 36612
rect 38778 36586 39778 36612
rect 41036 36586 42036 36612
rect 42094 36586 43094 36612
rect 43152 36586 44152 36612
rect 44210 36586 45210 36612
rect 45268 36586 46268 36612
rect 47624 36608 48624 36634
rect 48682 36608 49682 36634
rect 49740 36608 50740 36634
rect 50798 36608 51798 36634
rect 51856 36608 52856 36634
rect 54138 36622 55138 36648
rect 55196 36622 56196 36648
rect 56254 36622 57254 36648
rect 57312 36622 58312 36648
rect 58370 36622 59370 36648
rect 2004 36496 3004 36522
rect 3062 36496 4062 36522
rect 4120 36496 5120 36522
rect 5178 36496 6178 36522
rect 6236 36496 7236 36522
rect 8518 36504 9518 36530
rect 9576 36504 10576 36530
rect 10634 36504 11634 36530
rect 11692 36504 12692 36530
rect 12750 36504 13750 36530
rect 15024 36512 16024 36538
rect 16082 36512 17082 36538
rect 17140 36512 18140 36538
rect 18198 36512 19198 36538
rect 19256 36512 20256 36538
rect 21766 36522 22300 36564
rect 22804 36522 23338 36564
rect 23922 36522 24456 36564
rect 24938 36522 25472 36564
rect 26004 36522 26538 36564
rect 28288 36538 28822 36580
rect 29326 36538 29860 36580
rect 30444 36538 30978 36580
rect 31460 36538 31994 36580
rect 32526 36538 33060 36580
rect 34798 36544 35332 36586
rect 35836 36544 36370 36586
rect 36954 36544 37488 36586
rect 37970 36544 38504 36586
rect 39036 36544 39570 36586
rect 41288 36544 41822 36586
rect 42326 36544 42860 36586
rect 43444 36544 43978 36586
rect 44460 36544 44994 36586
rect 45526 36544 46060 36586
rect 47876 36566 48410 36608
rect 48914 36566 49448 36608
rect 50032 36566 50566 36608
rect 51048 36566 51582 36608
rect 52114 36566 52648 36608
rect 54390 36580 54924 36622
rect 55428 36580 55962 36622
rect 56546 36580 57080 36622
rect 57562 36580 58096 36622
rect 58628 36580 59162 36622
rect 2004 35470 3004 35496
rect 3062 35470 4062 35496
rect 4120 35470 5120 35496
rect 5178 35470 6178 35496
rect 6236 35470 7236 35496
rect 2292 35428 2826 35470
rect 3248 35428 3782 35470
rect 4356 35428 4890 35470
rect 5462 35428 5996 35470
rect 6492 35428 7026 35470
rect 2004 35402 3004 35428
rect 3062 35402 4062 35428
rect 4120 35402 5120 35428
rect 5178 35402 6178 35428
rect 6236 35402 7236 35428
rect 8518 35478 9518 35504
rect 9576 35478 10576 35504
rect 10634 35478 11634 35504
rect 11692 35478 12692 35504
rect 12750 35478 13750 35504
rect 8806 35436 9340 35478
rect 9762 35436 10296 35478
rect 10870 35436 11404 35478
rect 11976 35436 12510 35478
rect 13006 35436 13540 35478
rect 8518 35410 9518 35436
rect 9576 35410 10576 35436
rect 10634 35410 11634 35436
rect 11692 35410 12692 35436
rect 12750 35410 13750 35436
rect 2004 34376 3004 34402
rect 3062 34376 4062 34402
rect 4120 34376 5120 34402
rect 5178 34376 6178 34402
rect 6236 34376 7236 34402
rect 2228 34334 2762 34376
rect 3282 34334 3816 34376
rect 4334 34334 4868 34376
rect 5442 34334 5976 34376
rect 6498 34334 7032 34376
rect 2004 34308 3004 34334
rect 3062 34308 4062 34334
rect 4120 34308 5120 34334
rect 5178 34308 6178 34334
rect 6236 34308 7236 34334
rect 21514 36496 22514 36522
rect 22572 36496 23572 36522
rect 23630 36496 24630 36522
rect 24688 36496 25688 36522
rect 25746 36496 26746 36522
rect 28036 36512 29036 36538
rect 29094 36512 30094 36538
rect 30152 36512 31152 36538
rect 31210 36512 32210 36538
rect 32268 36512 33268 36538
rect 34546 36518 35546 36544
rect 35604 36518 36604 36544
rect 36662 36518 37662 36544
rect 37720 36518 38720 36544
rect 38778 36518 39778 36544
rect 41036 36518 42036 36544
rect 42094 36518 43094 36544
rect 43152 36518 44152 36544
rect 44210 36518 45210 36544
rect 45268 36518 46268 36544
rect 47624 36540 48624 36566
rect 48682 36540 49682 36566
rect 49740 36540 50740 36566
rect 50798 36540 51798 36566
rect 51856 36540 52856 36566
rect 54138 36554 55138 36580
rect 55196 36554 56196 36580
rect 56254 36554 57254 36580
rect 57312 36554 58312 36580
rect 58370 36554 59370 36580
rect 15024 35486 16024 35512
rect 16082 35486 17082 35512
rect 17140 35486 18140 35512
rect 18198 35486 19198 35512
rect 19256 35486 20256 35512
rect 15312 35444 15846 35486
rect 16268 35444 16802 35486
rect 17376 35444 17910 35486
rect 18482 35444 19016 35486
rect 19512 35444 20046 35486
rect 15024 35418 16024 35444
rect 16082 35418 17082 35444
rect 17140 35418 18140 35444
rect 18198 35418 19198 35444
rect 19256 35418 20256 35444
rect 8518 34384 9518 34410
rect 9576 34384 10576 34410
rect 10634 34384 11634 34410
rect 11692 34384 12692 34410
rect 12750 34384 13750 34410
rect 8742 34342 9276 34384
rect 9796 34342 10330 34384
rect 10848 34342 11382 34384
rect 11956 34342 12490 34384
rect 13012 34342 13546 34384
rect 8518 34316 9518 34342
rect 9576 34316 10576 34342
rect 10634 34316 11634 34342
rect 11692 34316 12692 34342
rect 12750 34316 13750 34342
rect 21514 35470 22514 35496
rect 22572 35470 23572 35496
rect 23630 35470 24630 35496
rect 24688 35470 25688 35496
rect 25746 35470 26746 35496
rect 21802 35428 22336 35470
rect 22758 35428 23292 35470
rect 23866 35428 24400 35470
rect 24972 35428 25506 35470
rect 26002 35428 26536 35470
rect 21514 35402 22514 35428
rect 22572 35402 23572 35428
rect 23630 35402 24630 35428
rect 24688 35402 25688 35428
rect 25746 35402 26746 35428
rect 15024 34392 16024 34418
rect 16082 34392 17082 34418
rect 17140 34392 18140 34418
rect 18198 34392 19198 34418
rect 19256 34392 20256 34418
rect 15248 34350 15782 34392
rect 16302 34350 16836 34392
rect 17354 34350 17888 34392
rect 18462 34350 18996 34392
rect 19518 34350 20052 34392
rect 15024 34324 16024 34350
rect 16082 34324 17082 34350
rect 17140 34324 18140 34350
rect 18198 34324 19198 34350
rect 19256 34324 20256 34350
rect 28036 35486 29036 35512
rect 29094 35486 30094 35512
rect 30152 35486 31152 35512
rect 31210 35486 32210 35512
rect 32268 35486 33268 35512
rect 28324 35444 28858 35486
rect 29280 35444 29814 35486
rect 30388 35444 30922 35486
rect 31494 35444 32028 35486
rect 32524 35444 33058 35486
rect 28036 35418 29036 35444
rect 29094 35418 30094 35444
rect 30152 35418 31152 35444
rect 31210 35418 32210 35444
rect 32268 35418 33268 35444
rect 21514 34376 22514 34402
rect 22572 34376 23572 34402
rect 23630 34376 24630 34402
rect 24688 34376 25688 34402
rect 25746 34376 26746 34402
rect 21738 34334 22272 34376
rect 22792 34334 23326 34376
rect 23844 34334 24378 34376
rect 24952 34334 25486 34376
rect 26008 34334 26542 34376
rect 21514 34308 22514 34334
rect 22572 34308 23572 34334
rect 23630 34308 24630 34334
rect 24688 34308 25688 34334
rect 25746 34308 26746 34334
rect 2004 33282 3004 33308
rect 3062 33282 4062 33308
rect 4120 33282 5120 33308
rect 5178 33282 6178 33308
rect 6236 33282 7236 33308
rect 8518 33290 9518 33316
rect 9576 33290 10576 33316
rect 10634 33290 11634 33316
rect 11692 33290 12692 33316
rect 12750 33290 13750 33316
rect 15024 33298 16024 33324
rect 16082 33298 17082 33324
rect 17140 33298 18140 33324
rect 18198 33298 19198 33324
rect 19256 33298 20256 33324
rect 34546 35492 35546 35518
rect 35604 35492 36604 35518
rect 36662 35492 37662 35518
rect 37720 35492 38720 35518
rect 38778 35492 39778 35518
rect 34834 35450 35368 35492
rect 35790 35450 36324 35492
rect 36898 35450 37432 35492
rect 38004 35450 38538 35492
rect 39034 35450 39568 35492
rect 34546 35424 35546 35450
rect 35604 35424 36604 35450
rect 36662 35424 37662 35450
rect 37720 35424 38720 35450
rect 38778 35424 39778 35450
rect 28036 34392 29036 34418
rect 29094 34392 30094 34418
rect 30152 34392 31152 34418
rect 31210 34392 32210 34418
rect 32268 34392 33268 34418
rect 28260 34350 28794 34392
rect 29314 34350 29848 34392
rect 30366 34350 30900 34392
rect 31474 34350 32008 34392
rect 32530 34350 33064 34392
rect 28036 34324 29036 34350
rect 29094 34324 30094 34350
rect 30152 34324 31152 34350
rect 31210 34324 32210 34350
rect 32268 34324 33268 34350
rect 41036 35492 42036 35518
rect 42094 35492 43094 35518
rect 43152 35492 44152 35518
rect 44210 35492 45210 35518
rect 45268 35492 46268 35518
rect 41324 35450 41858 35492
rect 42280 35450 42814 35492
rect 43388 35450 43922 35492
rect 44494 35450 45028 35492
rect 45524 35450 46058 35492
rect 41036 35424 42036 35450
rect 42094 35424 43094 35450
rect 43152 35424 44152 35450
rect 44210 35424 45210 35450
rect 45268 35424 46268 35450
rect 34546 34398 35546 34424
rect 35604 34398 36604 34424
rect 36662 34398 37662 34424
rect 37720 34398 38720 34424
rect 38778 34398 39778 34424
rect 34770 34356 35304 34398
rect 35824 34356 36358 34398
rect 36876 34356 37410 34398
rect 37984 34356 38518 34398
rect 39040 34356 39574 34398
rect 34546 34330 35546 34356
rect 35604 34330 36604 34356
rect 36662 34330 37662 34356
rect 37720 34330 38720 34356
rect 38778 34330 39778 34356
rect 47624 35514 48624 35540
rect 48682 35514 49682 35540
rect 49740 35514 50740 35540
rect 50798 35514 51798 35540
rect 51856 35514 52856 35540
rect 47912 35472 48446 35514
rect 48868 35472 49402 35514
rect 49976 35472 50510 35514
rect 51082 35472 51616 35514
rect 52112 35472 52646 35514
rect 47624 35446 48624 35472
rect 48682 35446 49682 35472
rect 49740 35446 50740 35472
rect 50798 35446 51798 35472
rect 51856 35446 52856 35472
rect 41036 34398 42036 34424
rect 42094 34398 43094 34424
rect 43152 34398 44152 34424
rect 44210 34398 45210 34424
rect 45268 34398 46268 34424
rect 41260 34356 41794 34398
rect 42314 34356 42848 34398
rect 43366 34356 43900 34398
rect 44474 34356 45008 34398
rect 45530 34356 46064 34398
rect 41036 34330 42036 34356
rect 42094 34330 43094 34356
rect 43152 34330 44152 34356
rect 44210 34330 45210 34356
rect 45268 34330 46268 34356
rect 63532 43632 64602 43690
rect 63532 43466 63810 43632
rect 64200 43466 64602 43632
rect 63532 43440 64602 43466
rect 67610 43584 68350 43686
rect 67610 43442 67818 43584
rect 62860 43348 65688 43440
rect 66654 43438 67818 43442
rect 68110 43442 68350 43584
rect 71304 43614 72242 43648
rect 71304 43456 71596 43614
rect 70462 43444 71596 43456
rect 71844 43456 72242 43614
rect 71844 43444 73290 43456
rect 68110 43438 69482 43442
rect 66654 43350 69482 43438
rect 70462 43364 73290 43444
rect 70156 43358 73388 43364
rect 62554 43342 65786 43348
rect 62554 43322 63154 43342
rect 63212 43322 63812 43342
rect 63870 43322 64470 43342
rect 64528 43322 65128 43342
rect 65186 43322 65786 43342
rect 66348 43344 69580 43350
rect 66348 43324 66948 43344
rect 67006 43324 67606 43344
rect 67664 43324 68264 43344
rect 68322 43324 68922 43344
rect 68980 43324 69580 43344
rect 70156 43338 70756 43358
rect 70814 43338 71414 43358
rect 71472 43338 72072 43358
rect 72130 43338 72730 43358
rect 72788 43338 73388 43358
rect 62554 42696 63154 42722
rect 63212 42696 63812 42722
rect 63870 42696 64470 42722
rect 64528 42696 65128 42722
rect 65186 42696 65786 42722
rect 62666 42654 62990 42696
rect 63332 42654 63656 42696
rect 63984 42654 64308 42696
rect 64694 42654 65018 42696
rect 65276 42654 65600 42696
rect 62554 42628 63154 42654
rect 63212 42628 63812 42654
rect 63870 42628 64470 42654
rect 64528 42628 65128 42654
rect 65186 42628 65786 42654
rect 66348 42698 66948 42724
rect 67006 42698 67606 42724
rect 67664 42698 68264 42724
rect 68322 42698 68922 42724
rect 68980 42698 69580 42724
rect 66460 42656 66784 42698
rect 67126 42656 67450 42698
rect 67778 42656 68102 42698
rect 68488 42656 68812 42698
rect 69070 42656 69394 42698
rect 62554 42002 63154 42028
rect 63212 42002 63812 42028
rect 63870 42002 64470 42028
rect 64528 42002 65128 42028
rect 65186 42002 65786 42028
rect 62672 41960 62996 42002
rect 63294 41960 63618 42002
rect 63918 41960 64242 42002
rect 64670 41960 64994 42002
rect 65240 41960 65564 42002
rect 62554 41934 63154 41960
rect 63212 41934 63812 41960
rect 63870 41934 64470 41960
rect 64528 41934 65128 41960
rect 65186 41934 65786 41960
rect 62554 41308 63154 41334
rect 63212 41308 63812 41334
rect 63870 41308 64470 41334
rect 64528 41308 65128 41334
rect 65186 41308 65786 41334
rect 62668 41266 62992 41308
rect 63360 41266 63684 41308
rect 63990 41266 64314 41308
rect 64678 41266 65002 41308
rect 65358 41266 65682 41308
rect 62554 41240 63154 41266
rect 63212 41240 63812 41266
rect 63870 41240 64470 41266
rect 64528 41240 65128 41266
rect 65186 41240 65786 41266
rect 66348 42630 66948 42656
rect 67006 42630 67606 42656
rect 67664 42630 68264 42656
rect 68322 42630 68922 42656
rect 68980 42630 69580 42656
rect 70156 42712 70756 42738
rect 70814 42712 71414 42738
rect 71472 42712 72072 42738
rect 72130 42712 72730 42738
rect 72788 42712 73388 42738
rect 70268 42670 70592 42712
rect 70934 42670 71258 42712
rect 71586 42670 71910 42712
rect 72296 42670 72620 42712
rect 72878 42670 73202 42712
rect 66348 42004 66948 42030
rect 67006 42004 67606 42030
rect 67664 42004 68264 42030
rect 68322 42004 68922 42030
rect 68980 42004 69580 42030
rect 66466 41962 66790 42004
rect 67088 41962 67412 42004
rect 67712 41962 68036 42004
rect 68464 41962 68788 42004
rect 69034 41962 69358 42004
rect 66348 41936 66948 41962
rect 67006 41936 67606 41962
rect 67664 41936 68264 41962
rect 68322 41936 68922 41962
rect 68980 41936 69580 41962
rect 66348 41310 66948 41336
rect 67006 41310 67606 41336
rect 67664 41310 68264 41336
rect 68322 41310 68922 41336
rect 68980 41310 69580 41336
rect 66462 41268 66786 41310
rect 67154 41268 67478 41310
rect 67784 41268 68108 41310
rect 68472 41268 68796 41310
rect 69152 41268 69476 41310
rect 66348 41242 66948 41268
rect 67006 41242 67606 41268
rect 67664 41242 68264 41268
rect 68322 41242 68922 41268
rect 68980 41242 69580 41268
rect 70156 42644 70756 42670
rect 70814 42644 71414 42670
rect 71472 42644 72072 42670
rect 72130 42644 72730 42670
rect 72788 42644 73388 42670
rect 70156 42018 70756 42044
rect 70814 42018 71414 42044
rect 71472 42018 72072 42044
rect 72130 42018 72730 42044
rect 72788 42018 73388 42044
rect 70274 41976 70598 42018
rect 70896 41976 71220 42018
rect 71520 41976 71844 42018
rect 72272 41976 72596 42018
rect 72842 41976 73166 42018
rect 70156 41950 70756 41976
rect 70814 41950 71414 41976
rect 71472 41950 72072 41976
rect 72130 41950 72730 41976
rect 72788 41950 73388 41976
rect 70156 41324 70756 41350
rect 70814 41324 71414 41350
rect 71472 41324 72072 41350
rect 72130 41324 72730 41350
rect 72788 41324 73388 41350
rect 70270 41282 70594 41324
rect 70962 41282 71286 41324
rect 71592 41282 71916 41324
rect 72280 41282 72604 41324
rect 72960 41282 73284 41324
rect 70156 41256 70756 41282
rect 70814 41256 71414 41282
rect 71472 41256 72072 41282
rect 72130 41256 72730 41282
rect 72788 41256 73388 41282
rect 62554 40614 63154 40640
rect 63212 40614 63812 40640
rect 63870 40614 64470 40640
rect 64528 40614 65128 40640
rect 65186 40614 65786 40640
rect 66348 40616 66948 40642
rect 67006 40616 67606 40642
rect 67664 40616 68264 40642
rect 68322 40616 68922 40642
rect 68980 40616 69580 40642
rect 70156 40630 70756 40656
rect 70814 40630 71414 40656
rect 71472 40630 72072 40656
rect 72130 40630 72730 40656
rect 72788 40630 73388 40656
rect 62646 40572 62970 40614
rect 63314 40572 63638 40614
rect 63998 40572 64322 40614
rect 64696 40572 65020 40614
rect 65322 40572 65646 40614
rect 66440 40574 66764 40616
rect 67108 40574 67432 40616
rect 67792 40574 68116 40616
rect 68490 40574 68814 40616
rect 69116 40574 69440 40616
rect 70248 40588 70572 40630
rect 70916 40588 71240 40630
rect 71600 40588 71924 40630
rect 72298 40588 72622 40630
rect 72924 40588 73248 40630
rect 62554 40546 63154 40572
rect 63212 40546 63812 40572
rect 63870 40546 64470 40572
rect 64528 40546 65128 40572
rect 65186 40546 65786 40572
rect 66348 40548 66948 40574
rect 67006 40548 67606 40574
rect 67664 40548 68264 40574
rect 68322 40548 68922 40574
rect 68980 40548 69580 40574
rect 70156 40562 70756 40588
rect 70814 40562 71414 40588
rect 71472 40562 72072 40588
rect 72130 40562 72730 40588
rect 72788 40562 73388 40588
rect 62554 39920 63154 39946
rect 63212 39920 63812 39946
rect 63870 39920 64470 39946
rect 64528 39920 65128 39946
rect 65186 39920 65786 39946
rect 66348 39922 66948 39948
rect 67006 39922 67606 39948
rect 67664 39922 68264 39948
rect 68322 39922 68922 39948
rect 68980 39922 69580 39948
rect 70156 39936 70756 39962
rect 70814 39936 71414 39962
rect 71472 39936 72072 39962
rect 72130 39936 72730 39962
rect 72788 39936 73388 39962
rect 54138 35528 55138 35554
rect 55196 35528 56196 35554
rect 56254 35528 57254 35554
rect 57312 35528 58312 35554
rect 58370 35528 59370 35554
rect 54426 35486 54960 35528
rect 55382 35486 55916 35528
rect 56490 35486 57024 35528
rect 57596 35486 58130 35528
rect 58626 35486 59160 35528
rect 54138 35460 55138 35486
rect 55196 35460 56196 35486
rect 56254 35460 57254 35486
rect 57312 35460 58312 35486
rect 58370 35460 59370 35486
rect 47624 34420 48624 34446
rect 48682 34420 49682 34446
rect 49740 34420 50740 34446
rect 50798 34420 51798 34446
rect 51856 34420 52856 34446
rect 47848 34378 48382 34420
rect 48902 34378 49436 34420
rect 49954 34378 50488 34420
rect 51062 34378 51596 34420
rect 52118 34378 52652 34420
rect 47624 34352 48624 34378
rect 48682 34352 49682 34378
rect 49740 34352 50740 34378
rect 50798 34352 51798 34378
rect 51856 34352 52856 34378
rect 54138 34434 55138 34460
rect 55196 34434 56196 34460
rect 56254 34434 57254 34460
rect 57312 34434 58312 34460
rect 58370 34434 59370 34460
rect 78392 39510 78904 39542
rect 78392 39414 78536 39510
rect 77520 39406 78536 39414
rect 78796 39414 78904 39510
rect 80846 39538 81140 39582
rect 78796 39406 79646 39414
rect 77520 39334 79646 39406
rect 80846 39410 80866 39538
rect 81116 39410 81140 39538
rect 80846 39408 81140 39410
rect 84954 39524 85480 39568
rect 84954 39412 85060 39524
rect 85316 39412 85480 39524
rect 84954 39408 85480 39412
rect 77216 39332 79790 39334
rect 77216 39308 77816 39332
rect 77874 39308 78474 39332
rect 78532 39308 79132 39332
rect 79190 39308 79790 39332
rect 80846 39328 82972 39408
rect 84156 39328 86282 39408
rect 80542 39326 83116 39328
rect 80542 39302 81142 39326
rect 81200 39302 81800 39326
rect 81858 39302 82458 39326
rect 82516 39302 83116 39326
rect 83852 39326 86426 39328
rect 83852 39302 84452 39326
rect 84510 39302 85110 39326
rect 85168 39302 85768 39326
rect 85826 39302 86426 39326
rect 77216 38682 77816 38708
rect 77874 38682 78474 38708
rect 78532 38682 79132 38708
rect 79190 38682 79790 38708
rect 77374 38640 77706 38682
rect 78020 38640 78352 38682
rect 78732 38640 79064 38682
rect 79322 38640 79654 38682
rect 77216 38614 77816 38640
rect 77874 38614 78474 38640
rect 78532 38614 79132 38640
rect 79190 38614 79790 38640
rect 77216 37988 77816 38014
rect 77874 37988 78474 38014
rect 78532 37988 79132 38014
rect 79190 37988 79790 38014
rect 77338 37946 77670 37988
rect 78044 37946 78376 37988
rect 78706 37946 79038 37988
rect 79284 37946 79616 37988
rect 77216 37920 77816 37946
rect 77874 37920 78474 37946
rect 78532 37920 79132 37946
rect 79190 37920 79790 37946
rect 77216 37294 77816 37320
rect 77874 37294 78474 37320
rect 78532 37294 79132 37320
rect 79190 37294 79790 37320
rect 77342 37252 77674 37294
rect 78046 37252 78378 37294
rect 78684 37252 79016 37294
rect 79328 37252 79660 37294
rect 77216 37226 77816 37252
rect 77874 37226 78474 37252
rect 78532 37226 79132 37252
rect 79190 37226 79790 37252
rect 77216 36600 77816 36626
rect 77874 36600 78474 36626
rect 78532 36600 79132 36626
rect 79190 36600 79790 36626
rect 77336 36558 77668 36600
rect 78016 36558 78348 36600
rect 78700 36558 79032 36600
rect 79334 36558 79666 36600
rect 77216 36532 77816 36558
rect 77874 36532 78474 36558
rect 78532 36532 79132 36558
rect 79190 36532 79790 36558
rect 77216 35906 77816 35932
rect 77874 35906 78474 35932
rect 78532 35906 79132 35932
rect 79190 35906 79790 35932
rect 77330 35864 77662 35906
rect 78046 35864 78378 35906
rect 78676 35864 79008 35906
rect 79348 35864 79680 35906
rect 77216 35838 77816 35864
rect 77874 35838 78474 35864
rect 78532 35838 79132 35864
rect 79190 35838 79790 35864
rect 80542 38676 81142 38702
rect 81200 38676 81800 38702
rect 81858 38676 82458 38702
rect 82516 38676 83116 38702
rect 80700 38634 81032 38676
rect 81346 38634 81678 38676
rect 82058 38634 82390 38676
rect 82648 38634 82980 38676
rect 80542 38608 81142 38634
rect 81200 38608 81800 38634
rect 81858 38608 82458 38634
rect 82516 38608 83116 38634
rect 80542 37982 81142 38008
rect 81200 37982 81800 38008
rect 81858 37982 82458 38008
rect 82516 37982 83116 38008
rect 80664 37940 80996 37982
rect 81370 37940 81702 37982
rect 82032 37940 82364 37982
rect 82610 37940 82942 37982
rect 80542 37914 81142 37940
rect 81200 37914 81800 37940
rect 81858 37914 82458 37940
rect 82516 37914 83116 37940
rect 80542 37288 81142 37314
rect 81200 37288 81800 37314
rect 81858 37288 82458 37314
rect 82516 37288 83116 37314
rect 80668 37246 81000 37288
rect 81372 37246 81704 37288
rect 82010 37246 82342 37288
rect 82654 37246 82986 37288
rect 80542 37220 81142 37246
rect 81200 37220 81800 37246
rect 81858 37220 82458 37246
rect 82516 37220 83116 37246
rect 80542 36594 81142 36620
rect 81200 36594 81800 36620
rect 81858 36594 82458 36620
rect 82516 36594 83116 36620
rect 80662 36552 80994 36594
rect 81342 36552 81674 36594
rect 82026 36552 82358 36594
rect 82660 36552 82992 36594
rect 80542 36526 81142 36552
rect 81200 36526 81800 36552
rect 81858 36526 82458 36552
rect 82516 36526 83116 36552
rect 80542 35900 81142 35926
rect 81200 35900 81800 35926
rect 81858 35900 82458 35926
rect 82516 35900 83116 35926
rect 80656 35858 80988 35900
rect 81372 35858 81704 35900
rect 82002 35858 82334 35900
rect 82674 35858 83006 35900
rect 80542 35832 81142 35858
rect 81200 35832 81800 35858
rect 81858 35832 82458 35858
rect 82516 35832 83116 35858
rect 77216 35212 77816 35238
rect 77874 35212 78474 35238
rect 78532 35212 79132 35238
rect 79190 35212 79790 35238
rect 83852 38676 84452 38702
rect 84510 38676 85110 38702
rect 85168 38676 85768 38702
rect 85826 38676 86426 38702
rect 84010 38634 84342 38676
rect 84656 38634 84988 38676
rect 85368 38634 85700 38676
rect 85958 38634 86290 38676
rect 83852 38608 84452 38634
rect 84510 38608 85110 38634
rect 85168 38608 85768 38634
rect 85826 38608 86426 38634
rect 83852 37982 84452 38008
rect 84510 37982 85110 38008
rect 85168 37982 85768 38008
rect 85826 37982 86426 38008
rect 83974 37940 84306 37982
rect 84680 37940 85012 37982
rect 85342 37940 85674 37982
rect 85920 37940 86252 37982
rect 83852 37914 84452 37940
rect 84510 37914 85110 37940
rect 85168 37914 85768 37940
rect 85826 37914 86426 37940
rect 83852 37288 84452 37314
rect 84510 37288 85110 37314
rect 85168 37288 85768 37314
rect 85826 37288 86426 37314
rect 83978 37246 84310 37288
rect 84682 37246 85014 37288
rect 85320 37246 85652 37288
rect 85964 37246 86296 37288
rect 83852 37220 84452 37246
rect 84510 37220 85110 37246
rect 85168 37220 85768 37246
rect 85826 37220 86426 37246
rect 83852 36594 84452 36620
rect 84510 36594 85110 36620
rect 85168 36594 85768 36620
rect 85826 36594 86426 36620
rect 83972 36552 84304 36594
rect 84652 36552 84984 36594
rect 85336 36552 85668 36594
rect 85970 36552 86302 36594
rect 83852 36526 84452 36552
rect 84510 36526 85110 36552
rect 85168 36526 85768 36552
rect 85826 36526 86426 36552
rect 83852 35900 84452 35926
rect 84510 35900 85110 35926
rect 85168 35900 85768 35926
rect 85826 35900 86426 35926
rect 83966 35858 84298 35900
rect 84682 35858 85014 35900
rect 85312 35858 85644 35900
rect 85984 35858 86316 35900
rect 83852 35832 84452 35858
rect 84510 35832 85110 35858
rect 85168 35832 85768 35858
rect 85826 35832 86426 35858
rect 80542 35206 81142 35232
rect 81200 35206 81800 35232
rect 81858 35206 82458 35232
rect 82516 35206 83116 35232
rect 83852 35206 84452 35232
rect 84510 35206 85110 35232
rect 85168 35206 85768 35232
rect 85826 35206 86426 35232
rect 54362 34392 54896 34434
rect 55416 34392 55950 34434
rect 56468 34392 57002 34434
rect 57576 34392 58110 34434
rect 58632 34392 59166 34434
rect 54138 34366 55138 34392
rect 55196 34366 56196 34392
rect 56254 34366 57254 34392
rect 57312 34366 58312 34392
rect 58370 34366 59370 34392
rect 2256 33240 2790 33282
rect 3354 33240 3888 33282
rect 4382 33240 4916 33282
rect 5346 33240 5880 33282
rect 6446 33240 6980 33282
rect 8770 33248 9304 33290
rect 9868 33248 10402 33290
rect 10896 33248 11430 33290
rect 11860 33248 12394 33290
rect 12960 33248 13494 33290
rect 15276 33256 15810 33298
rect 16374 33256 16908 33298
rect 17402 33256 17936 33298
rect 18366 33256 18900 33298
rect 19466 33256 20000 33298
rect 21514 33282 22514 33308
rect 22572 33282 23572 33308
rect 23630 33282 24630 33308
rect 24688 33282 25688 33308
rect 25746 33282 26746 33308
rect 28036 33298 29036 33324
rect 29094 33298 30094 33324
rect 30152 33298 31152 33324
rect 31210 33298 32210 33324
rect 32268 33298 33268 33324
rect 34546 33304 35546 33330
rect 35604 33304 36604 33330
rect 36662 33304 37662 33330
rect 37720 33304 38720 33330
rect 38778 33304 39778 33330
rect 41036 33304 42036 33330
rect 42094 33304 43094 33330
rect 43152 33304 44152 33330
rect 44210 33304 45210 33330
rect 45268 33304 46268 33330
rect 47624 33326 48624 33352
rect 48682 33326 49682 33352
rect 49740 33326 50740 33352
rect 50798 33326 51798 33352
rect 51856 33326 52856 33352
rect 54138 33340 55138 33366
rect 55196 33340 56196 33366
rect 56254 33340 57254 33366
rect 57312 33340 58312 33366
rect 58370 33340 59370 33366
rect 2004 33214 3004 33240
rect 3062 33214 4062 33240
rect 4120 33214 5120 33240
rect 5178 33214 6178 33240
rect 6236 33214 7236 33240
rect 8518 33222 9518 33248
rect 9576 33222 10576 33248
rect 10634 33222 11634 33248
rect 11692 33222 12692 33248
rect 12750 33222 13750 33248
rect 15024 33230 16024 33256
rect 16082 33230 17082 33256
rect 17140 33230 18140 33256
rect 18198 33230 19198 33256
rect 19256 33230 20256 33256
rect 21766 33240 22300 33282
rect 22864 33240 23398 33282
rect 23892 33240 24426 33282
rect 24856 33240 25390 33282
rect 25956 33240 26490 33282
rect 28288 33256 28822 33298
rect 29386 33256 29920 33298
rect 30414 33256 30948 33298
rect 31378 33256 31912 33298
rect 32478 33256 33012 33298
rect 34798 33262 35332 33304
rect 35896 33262 36430 33304
rect 36924 33262 37458 33304
rect 37888 33262 38422 33304
rect 38988 33262 39522 33304
rect 41288 33262 41822 33304
rect 42386 33262 42920 33304
rect 43414 33262 43948 33304
rect 44378 33262 44912 33304
rect 45478 33262 46012 33304
rect 47876 33284 48410 33326
rect 48974 33284 49508 33326
rect 50002 33284 50536 33326
rect 50966 33284 51500 33326
rect 52066 33284 52600 33326
rect 54390 33298 54924 33340
rect 55488 33298 56022 33340
rect 56516 33298 57050 33340
rect 57480 33298 58014 33340
rect 58580 33298 59114 33340
rect 21514 33214 22514 33240
rect 22572 33214 23572 33240
rect 23630 33214 24630 33240
rect 24688 33214 25688 33240
rect 25746 33214 26746 33240
rect 28036 33230 29036 33256
rect 29094 33230 30094 33256
rect 30152 33230 31152 33256
rect 31210 33230 32210 33256
rect 32268 33230 33268 33256
rect 34546 33236 35546 33262
rect 35604 33236 36604 33262
rect 36662 33236 37662 33262
rect 37720 33236 38720 33262
rect 38778 33236 39778 33262
rect 41036 33236 42036 33262
rect 42094 33236 43094 33262
rect 43152 33236 44152 33262
rect 44210 33236 45210 33262
rect 45268 33236 46268 33262
rect 47624 33258 48624 33284
rect 48682 33258 49682 33284
rect 49740 33258 50740 33284
rect 50798 33258 51798 33284
rect 51856 33258 52856 33284
rect 54138 33272 55138 33298
rect 55196 33272 56196 33298
rect 56254 33272 57254 33298
rect 57312 33272 58312 33298
rect 58370 33272 59370 33298
rect 2004 32188 3004 32214
rect 3062 32188 4062 32214
rect 4120 32188 5120 32214
rect 5178 32188 6178 32214
rect 6236 32188 7236 32214
rect 8518 32204 9518 32222
rect 9576 32204 10576 32222
rect 10634 32204 11634 32222
rect 11692 32204 12692 32222
rect 12750 32204 13750 32222
rect 15024 32210 16024 32230
rect 16082 32210 17082 32230
rect 17140 32210 18140 32230
rect 18198 32210 19198 32230
rect 19256 32210 20256 32230
rect 47624 32240 48624 32258
rect 48682 32240 49682 32258
rect 49740 32240 50740 32258
rect 50798 32240 51798 32258
rect 51856 32240 52856 32258
rect 54138 32254 55138 32272
rect 55196 32254 56196 32272
rect 56254 32254 57254 32272
rect 57312 32254 58312 32272
rect 58370 32254 59370 32272
rect 54138 32246 59370 32254
rect 15024 32204 20256 32210
rect 8518 32196 13750 32204
rect 2556 31824 2722 32188
rect 3390 31824 3556 32188
rect 4488 31824 4654 32188
rect 5488 31824 5654 32188
rect 6552 31824 6718 32188
rect 8948 32116 13560 32196
rect 11126 31832 11498 32116
rect 15460 32070 20002 32204
rect 21514 32196 22514 32214
rect 22572 32196 23572 32214
rect 23630 32196 24630 32214
rect 24688 32196 25688 32214
rect 25746 32196 26746 32214
rect 28036 32212 29036 32230
rect 29094 32212 30094 32230
rect 30152 32212 31152 32230
rect 31210 32212 32210 32230
rect 32268 32212 33268 32230
rect 28036 32204 33268 32212
rect 34546 32220 35546 32236
rect 35604 32220 36604 32236
rect 36662 32220 37662 32236
rect 37720 32220 38720 32236
rect 38778 32220 39778 32236
rect 34546 32210 39778 32220
rect 41036 32218 42036 32236
rect 42094 32218 43094 32236
rect 43152 32218 44152 32236
rect 44210 32218 45210 32236
rect 45268 32218 46268 32236
rect 47624 32232 52856 32240
rect 41036 32210 46268 32218
rect 21514 32188 26746 32196
rect 18756 31840 18920 32070
rect 21956 31988 26436 32188
rect 28512 32020 32992 32204
rect 35004 32034 39492 32210
rect 2454 31782 7080 31824
rect 8968 31790 13594 31832
rect 15474 31798 20100 31840
rect 23218 31824 23516 31988
rect 30016 31840 30314 32020
rect 36446 31846 36744 32034
rect 41490 32026 45974 32210
rect 48048 32050 52548 32232
rect 43084 31846 43382 32026
rect 50214 31868 50512 32050
rect 54598 32010 59064 32246
rect 55708 31882 55934 32010
rect 15024 31792 20256 31798
rect 8518 31784 13750 31790
rect 2004 31776 7236 31782
rect 2004 31756 3004 31776
rect 3062 31756 4062 31776
rect 4120 31756 5120 31776
rect 5178 31756 6178 31776
rect 6236 31756 7236 31776
rect 8518 31764 9518 31784
rect 9576 31764 10576 31784
rect 10634 31764 11634 31784
rect 11692 31764 12692 31784
rect 12750 31764 13750 31784
rect 15024 31772 16024 31792
rect 16082 31772 17082 31792
rect 17140 31772 18140 31792
rect 18198 31772 19198 31792
rect 19256 31772 20256 31792
rect 21964 31782 26590 31824
rect 28486 31798 33112 31840
rect 34996 31804 39622 31846
rect 41486 31804 46112 31846
rect 48074 31826 52700 31868
rect 54588 31840 59214 31882
rect 54138 31834 59370 31840
rect 47624 31820 52856 31826
rect 34546 31798 39778 31804
rect 28036 31792 33268 31798
rect 21514 31776 26746 31782
rect 21514 31756 22514 31776
rect 22572 31756 23572 31776
rect 23630 31756 24630 31776
rect 24688 31756 25688 31776
rect 25746 31756 26746 31776
rect 28036 31772 29036 31792
rect 29094 31772 30094 31792
rect 30152 31772 31152 31792
rect 31210 31772 32210 31792
rect 32268 31772 33268 31792
rect 34546 31778 35546 31798
rect 35604 31778 36604 31798
rect 36662 31778 37662 31798
rect 37720 31778 38720 31798
rect 38778 31778 39778 31798
rect 41036 31798 46268 31804
rect 47624 31800 48624 31820
rect 48682 31800 49682 31820
rect 49740 31800 50740 31820
rect 50798 31800 51798 31820
rect 51856 31800 52856 31820
rect 54138 31814 55138 31834
rect 55196 31814 56196 31834
rect 56254 31814 57254 31834
rect 57312 31814 58312 31834
rect 58370 31814 59370 31834
rect 41036 31778 42036 31798
rect 42094 31794 44152 31798
rect 42094 31778 43094 31794
rect 43152 31778 44152 31794
rect 44210 31778 45210 31798
rect 45268 31778 46268 31798
rect 2004 30730 3004 30756
rect 3062 30730 4062 30756
rect 4120 30730 5120 30756
rect 5178 30730 6178 30756
rect 6236 30730 7236 30756
rect 8518 30738 9518 30764
rect 9576 30738 10576 30764
rect 10634 30738 11634 30764
rect 11692 30738 12692 30764
rect 12750 30738 13750 30764
rect 15024 30746 16024 30772
rect 16082 30746 17082 30772
rect 17140 30746 18140 30772
rect 18198 30746 19198 30772
rect 19256 30746 20256 30772
rect 2256 30688 2790 30730
rect 3294 30688 3828 30730
rect 4412 30688 4946 30730
rect 5428 30688 5962 30730
rect 6494 30688 7028 30730
rect 8770 30696 9304 30738
rect 9808 30696 10342 30738
rect 10926 30696 11460 30738
rect 11942 30696 12476 30738
rect 13008 30696 13542 30738
rect 15276 30704 15810 30746
rect 16314 30704 16848 30746
rect 17432 30704 17966 30746
rect 18448 30704 18982 30746
rect 19514 30704 20048 30746
rect 21514 30730 22514 30756
rect 22572 30730 23572 30756
rect 23630 30730 24630 30756
rect 24688 30730 25688 30756
rect 25746 30730 26746 30756
rect 28036 30746 29036 30772
rect 29094 30746 30094 30772
rect 30152 30746 31152 30772
rect 31210 30746 32210 30772
rect 32268 30746 33268 30772
rect 34546 30752 35546 30778
rect 35604 30752 36604 30778
rect 36662 30752 37662 30778
rect 37720 30752 38720 30778
rect 38778 30752 39778 30778
rect 41036 30752 42036 30778
rect 42094 30752 43094 30778
rect 43152 30752 44152 30778
rect 44210 30752 45210 30778
rect 45268 30752 46268 30778
rect 47624 30774 48624 30800
rect 48682 30774 49682 30800
rect 49740 30774 50740 30800
rect 50798 30774 51798 30800
rect 51856 30774 52856 30800
rect 54138 30788 55138 30814
rect 55196 30788 56196 30814
rect 56254 30788 57254 30814
rect 57312 30788 58312 30814
rect 58370 30788 59370 30814
rect 2004 30662 3004 30688
rect 3062 30662 4062 30688
rect 4120 30662 5120 30688
rect 5178 30662 6178 30688
rect 6236 30662 7236 30688
rect 8518 30670 9518 30696
rect 9576 30670 10576 30696
rect 10634 30670 11634 30696
rect 11692 30670 12692 30696
rect 12750 30670 13750 30696
rect 15024 30678 16024 30704
rect 16082 30678 17082 30704
rect 17140 30678 18140 30704
rect 18198 30678 19198 30704
rect 19256 30678 20256 30704
rect 21766 30688 22300 30730
rect 22804 30688 23338 30730
rect 23922 30688 24456 30730
rect 24938 30688 25472 30730
rect 26004 30688 26538 30730
rect 28288 30704 28822 30746
rect 29326 30704 29860 30746
rect 30444 30704 30978 30746
rect 31460 30704 31994 30746
rect 32526 30704 33060 30746
rect 34798 30710 35332 30752
rect 35836 30710 36370 30752
rect 36954 30710 37488 30752
rect 37970 30710 38504 30752
rect 39036 30710 39570 30752
rect 41288 30710 41822 30752
rect 42326 30710 42860 30752
rect 43444 30710 43978 30752
rect 44460 30710 44994 30752
rect 45526 30710 46060 30752
rect 47876 30732 48410 30774
rect 48914 30732 49448 30774
rect 50032 30732 50566 30774
rect 51048 30732 51582 30774
rect 52114 30732 52648 30774
rect 54390 30746 54924 30788
rect 55428 30746 55962 30788
rect 56546 30746 57080 30788
rect 57562 30746 58096 30788
rect 58628 30746 59162 30788
rect 2004 29636 3004 29662
rect 3062 29636 4062 29662
rect 4120 29636 5120 29662
rect 5178 29636 6178 29662
rect 6236 29636 7236 29662
rect 2292 29594 2826 29636
rect 3248 29594 3782 29636
rect 4356 29594 4890 29636
rect 5462 29594 5996 29636
rect 6492 29594 7026 29636
rect 2004 29568 3004 29594
rect 3062 29568 4062 29594
rect 4120 29568 5120 29594
rect 5178 29568 6178 29594
rect 6236 29568 7236 29594
rect 8518 29644 9518 29670
rect 9576 29644 10576 29670
rect 10634 29644 11634 29670
rect 11692 29644 12692 29670
rect 12750 29644 13750 29670
rect 8806 29602 9340 29644
rect 9762 29602 10296 29644
rect 10870 29602 11404 29644
rect 11976 29602 12510 29644
rect 13006 29602 13540 29644
rect 8518 29576 9518 29602
rect 9576 29576 10576 29602
rect 10634 29576 11634 29602
rect 11692 29576 12692 29602
rect 12750 29576 13750 29602
rect 2004 28542 3004 28568
rect 3062 28542 4062 28568
rect 4120 28542 5120 28568
rect 5178 28542 6178 28568
rect 6236 28542 7236 28568
rect 2228 28500 2762 28542
rect 3282 28500 3816 28542
rect 4334 28500 4868 28542
rect 5442 28500 5976 28542
rect 6498 28500 7032 28542
rect 2004 28474 3004 28500
rect 3062 28474 4062 28500
rect 4120 28474 5120 28500
rect 5178 28474 6178 28500
rect 6236 28474 7236 28500
rect 21514 30662 22514 30688
rect 22572 30662 23572 30688
rect 23630 30662 24630 30688
rect 24688 30662 25688 30688
rect 25746 30662 26746 30688
rect 28036 30678 29036 30704
rect 29094 30678 30094 30704
rect 30152 30678 31152 30704
rect 31210 30678 32210 30704
rect 32268 30678 33268 30704
rect 34546 30684 35546 30710
rect 35604 30684 36604 30710
rect 36662 30684 37662 30710
rect 37720 30684 38720 30710
rect 38778 30684 39778 30710
rect 41036 30684 42036 30710
rect 42094 30684 43094 30710
rect 43152 30684 44152 30710
rect 44210 30684 45210 30710
rect 45268 30684 46268 30710
rect 47624 30706 48624 30732
rect 48682 30706 49682 30732
rect 49740 30706 50740 30732
rect 50798 30706 51798 30732
rect 51856 30706 52856 30732
rect 54138 30720 55138 30746
rect 55196 30720 56196 30746
rect 56254 30720 57254 30746
rect 57312 30720 58312 30746
rect 58370 30720 59370 30746
rect 15024 29652 16024 29678
rect 16082 29652 17082 29678
rect 17140 29652 18140 29678
rect 18198 29652 19198 29678
rect 19256 29652 20256 29678
rect 15312 29610 15846 29652
rect 16268 29610 16802 29652
rect 17376 29610 17910 29652
rect 18482 29610 19016 29652
rect 19512 29610 20046 29652
rect 15024 29584 16024 29610
rect 16082 29584 17082 29610
rect 17140 29584 18140 29610
rect 18198 29584 19198 29610
rect 19256 29584 20256 29610
rect 8518 28550 9518 28576
rect 9576 28550 10576 28576
rect 10634 28550 11634 28576
rect 11692 28550 12692 28576
rect 12750 28550 13750 28576
rect 8742 28508 9276 28550
rect 9796 28508 10330 28550
rect 10848 28508 11382 28550
rect 11956 28508 12490 28550
rect 13012 28508 13546 28550
rect 8518 28482 9518 28508
rect 9576 28482 10576 28508
rect 10634 28482 11634 28508
rect 11692 28482 12692 28508
rect 12750 28482 13750 28508
rect 21514 29636 22514 29662
rect 22572 29636 23572 29662
rect 23630 29636 24630 29662
rect 24688 29636 25688 29662
rect 25746 29636 26746 29662
rect 21802 29594 22336 29636
rect 22758 29594 23292 29636
rect 23866 29594 24400 29636
rect 24972 29594 25506 29636
rect 26002 29594 26536 29636
rect 21514 29568 22514 29594
rect 22572 29568 23572 29594
rect 23630 29568 24630 29594
rect 24688 29568 25688 29594
rect 25746 29568 26746 29594
rect 15024 28558 16024 28584
rect 16082 28558 17082 28584
rect 17140 28558 18140 28584
rect 18198 28558 19198 28584
rect 19256 28558 20256 28584
rect 15248 28516 15782 28558
rect 16302 28516 16836 28558
rect 17354 28516 17888 28558
rect 18462 28516 18996 28558
rect 19518 28516 20052 28558
rect 15024 28490 16024 28516
rect 16082 28490 17082 28516
rect 17140 28490 18140 28516
rect 18198 28490 19198 28516
rect 19256 28490 20256 28516
rect 28036 29652 29036 29678
rect 29094 29652 30094 29678
rect 30152 29652 31152 29678
rect 31210 29652 32210 29678
rect 32268 29652 33268 29678
rect 28324 29610 28858 29652
rect 29280 29610 29814 29652
rect 30388 29610 30922 29652
rect 31494 29610 32028 29652
rect 32524 29610 33058 29652
rect 28036 29584 29036 29610
rect 29094 29584 30094 29610
rect 30152 29584 31152 29610
rect 31210 29584 32210 29610
rect 32268 29584 33268 29610
rect 21514 28542 22514 28568
rect 22572 28542 23572 28568
rect 23630 28542 24630 28568
rect 24688 28542 25688 28568
rect 25746 28542 26746 28568
rect 21738 28500 22272 28542
rect 22792 28500 23326 28542
rect 23844 28500 24378 28542
rect 24952 28500 25486 28542
rect 26008 28500 26542 28542
rect 21514 28474 22514 28500
rect 22572 28474 23572 28500
rect 23630 28474 24630 28500
rect 24688 28474 25688 28500
rect 25746 28474 26746 28500
rect 2004 27448 3004 27474
rect 3062 27448 4062 27474
rect 4120 27448 5120 27474
rect 5178 27448 6178 27474
rect 6236 27448 7236 27474
rect 8518 27456 9518 27482
rect 9576 27456 10576 27482
rect 10634 27456 11634 27482
rect 11692 27456 12692 27482
rect 12750 27456 13750 27482
rect 15024 27464 16024 27490
rect 16082 27464 17082 27490
rect 17140 27464 18140 27490
rect 18198 27464 19198 27490
rect 19256 27464 20256 27490
rect 34546 29658 35546 29684
rect 35604 29658 36604 29684
rect 36662 29658 37662 29684
rect 37720 29658 38720 29684
rect 38778 29658 39778 29684
rect 34834 29616 35368 29658
rect 35790 29616 36324 29658
rect 36898 29616 37432 29658
rect 38004 29616 38538 29658
rect 39034 29616 39568 29658
rect 34546 29590 35546 29616
rect 35604 29590 36604 29616
rect 36662 29590 37662 29616
rect 37720 29590 38720 29616
rect 38778 29590 39778 29616
rect 28036 28558 29036 28584
rect 29094 28558 30094 28584
rect 30152 28558 31152 28584
rect 31210 28558 32210 28584
rect 32268 28558 33268 28584
rect 28260 28516 28794 28558
rect 29314 28516 29848 28558
rect 30366 28516 30900 28558
rect 31474 28516 32008 28558
rect 32530 28516 33064 28558
rect 28036 28490 29036 28516
rect 29094 28490 30094 28516
rect 30152 28490 31152 28516
rect 31210 28490 32210 28516
rect 32268 28490 33268 28516
rect 41036 29658 42036 29684
rect 42094 29658 43094 29684
rect 43152 29658 44152 29684
rect 44210 29658 45210 29684
rect 45268 29658 46268 29684
rect 41324 29616 41858 29658
rect 42280 29616 42814 29658
rect 43388 29616 43922 29658
rect 44494 29616 45028 29658
rect 45524 29616 46058 29658
rect 41036 29590 42036 29616
rect 42094 29590 43094 29616
rect 43152 29590 44152 29616
rect 44210 29590 45210 29616
rect 45268 29590 46268 29616
rect 34546 28564 35546 28590
rect 35604 28564 36604 28590
rect 36662 28564 37662 28590
rect 37720 28564 38720 28590
rect 38778 28564 39778 28590
rect 34770 28522 35304 28564
rect 35824 28522 36358 28564
rect 36876 28522 37410 28564
rect 37984 28522 38518 28564
rect 39040 28522 39574 28564
rect 34546 28496 35546 28522
rect 35604 28496 36604 28522
rect 36662 28496 37662 28522
rect 37720 28496 38720 28522
rect 38778 28496 39778 28522
rect 47624 29680 48624 29706
rect 48682 29680 49682 29706
rect 49740 29680 50740 29706
rect 50798 29680 51798 29706
rect 51856 29680 52856 29706
rect 47912 29638 48446 29680
rect 48868 29638 49402 29680
rect 49976 29638 50510 29680
rect 51082 29638 51616 29680
rect 52112 29638 52646 29680
rect 47624 29612 48624 29638
rect 48682 29612 49682 29638
rect 49740 29612 50740 29638
rect 50798 29612 51798 29638
rect 51856 29612 52856 29638
rect 41036 28564 42036 28590
rect 42094 28564 43094 28590
rect 43152 28564 44152 28590
rect 44210 28564 45210 28590
rect 45268 28564 46268 28590
rect 41260 28522 41794 28564
rect 42314 28522 42848 28564
rect 43366 28522 43900 28564
rect 44474 28522 45008 28564
rect 45530 28522 46064 28564
rect 41036 28496 42036 28522
rect 42094 28496 43094 28522
rect 43152 28496 44152 28522
rect 44210 28496 45210 28522
rect 45268 28496 46268 28522
rect 54138 29694 55138 29720
rect 55196 29694 56196 29720
rect 56254 29694 57254 29720
rect 57312 29694 58312 29720
rect 58370 29694 59370 29720
rect 54426 29652 54960 29694
rect 55382 29652 55916 29694
rect 56490 29652 57024 29694
rect 57596 29652 58130 29694
rect 58626 29652 59160 29694
rect 54138 29626 55138 29652
rect 55196 29626 56196 29652
rect 56254 29626 57254 29652
rect 57312 29626 58312 29652
rect 58370 29626 59370 29652
rect 47624 28586 48624 28612
rect 48682 28586 49682 28612
rect 49740 28586 50740 28612
rect 50798 28586 51798 28612
rect 51856 28586 52856 28612
rect 47848 28544 48382 28586
rect 48902 28544 49436 28586
rect 49954 28544 50488 28586
rect 51062 28544 51596 28586
rect 52118 28544 52652 28586
rect 47624 28518 48624 28544
rect 48682 28518 49682 28544
rect 49740 28518 50740 28544
rect 50798 28518 51798 28544
rect 51856 28518 52856 28544
rect 54138 28600 55138 28626
rect 55196 28600 56196 28626
rect 56254 28600 57254 28626
rect 57312 28600 58312 28626
rect 58370 28600 59370 28626
rect 54362 28558 54896 28600
rect 55416 28558 55950 28600
rect 56468 28558 57002 28600
rect 57576 28558 58110 28600
rect 58632 28558 59166 28600
rect 54138 28532 55138 28558
rect 55196 28532 56196 28558
rect 56254 28532 57254 28558
rect 57312 28532 58312 28558
rect 58370 28532 59370 28558
rect 2256 27406 2790 27448
rect 3354 27406 3888 27448
rect 4382 27406 4916 27448
rect 5346 27406 5880 27448
rect 6446 27406 6980 27448
rect 8770 27414 9304 27456
rect 9868 27414 10402 27456
rect 10896 27414 11430 27456
rect 11860 27414 12394 27456
rect 12960 27414 13494 27456
rect 15276 27422 15810 27464
rect 16374 27422 16908 27464
rect 17402 27422 17936 27464
rect 18366 27422 18900 27464
rect 19466 27422 20000 27464
rect 21514 27448 22514 27474
rect 22572 27448 23572 27474
rect 23630 27448 24630 27474
rect 24688 27448 25688 27474
rect 25746 27448 26746 27474
rect 28036 27464 29036 27490
rect 29094 27464 30094 27490
rect 30152 27464 31152 27490
rect 31210 27464 32210 27490
rect 32268 27464 33268 27490
rect 34546 27470 35546 27496
rect 35604 27470 36604 27496
rect 36662 27470 37662 27496
rect 37720 27470 38720 27496
rect 38778 27470 39778 27496
rect 41036 27470 42036 27496
rect 42094 27470 43094 27496
rect 43152 27470 44152 27496
rect 44210 27470 45210 27496
rect 45268 27470 46268 27496
rect 47624 27492 48624 27518
rect 48682 27492 49682 27518
rect 49740 27492 50740 27518
rect 50798 27492 51798 27518
rect 51856 27492 52856 27518
rect 54138 27506 55138 27532
rect 55196 27506 56196 27532
rect 56254 27506 57254 27532
rect 57312 27506 58312 27532
rect 58370 27506 59370 27532
rect 2004 27380 3004 27406
rect 3062 27380 4062 27406
rect 4120 27380 5120 27406
rect 5178 27380 6178 27406
rect 6236 27380 7236 27406
rect 8518 27388 9518 27414
rect 9576 27388 10576 27414
rect 10634 27388 11634 27414
rect 11692 27388 12692 27414
rect 12750 27388 13750 27414
rect 15024 27396 16024 27422
rect 16082 27396 17082 27422
rect 17140 27396 18140 27422
rect 18198 27396 19198 27422
rect 19256 27396 20256 27422
rect 21766 27406 22300 27448
rect 22864 27406 23398 27448
rect 23892 27406 24426 27448
rect 24856 27406 25390 27448
rect 25956 27406 26490 27448
rect 28288 27422 28822 27464
rect 29386 27422 29920 27464
rect 30414 27422 30948 27464
rect 31378 27422 31912 27464
rect 32478 27422 33012 27464
rect 34798 27428 35332 27470
rect 35896 27428 36430 27470
rect 36924 27428 37458 27470
rect 37888 27428 38422 27470
rect 38988 27428 39522 27470
rect 41288 27428 41822 27470
rect 42386 27428 42920 27470
rect 43414 27428 43948 27470
rect 44378 27428 44912 27470
rect 45478 27428 46012 27470
rect 47876 27450 48410 27492
rect 48974 27450 49508 27492
rect 50002 27450 50536 27492
rect 50966 27450 51500 27492
rect 52066 27450 52600 27492
rect 54390 27464 54924 27506
rect 55488 27464 56022 27506
rect 56516 27464 57050 27506
rect 57480 27464 58014 27506
rect 58580 27464 59114 27506
rect 21514 27380 22514 27406
rect 22572 27380 23572 27406
rect 23630 27380 24630 27406
rect 24688 27380 25688 27406
rect 25746 27380 26746 27406
rect 28036 27396 29036 27422
rect 29094 27396 30094 27422
rect 30152 27396 31152 27422
rect 31210 27396 32210 27422
rect 32268 27396 33268 27422
rect 34546 27402 35546 27428
rect 35604 27402 36604 27428
rect 36662 27402 37662 27428
rect 37720 27402 38720 27428
rect 38778 27402 39778 27428
rect 41036 27402 42036 27428
rect 42094 27402 43094 27428
rect 43152 27402 44152 27428
rect 44210 27402 45210 27428
rect 45268 27402 46268 27428
rect 47624 27424 48624 27450
rect 48682 27424 49682 27450
rect 49740 27424 50740 27450
rect 50798 27424 51798 27450
rect 51856 27424 52856 27450
rect 54138 27438 55138 27464
rect 55196 27438 56196 27464
rect 56254 27438 57254 27464
rect 57312 27438 58312 27464
rect 58370 27438 59370 27464
rect 2004 26354 3004 26380
rect 3062 26354 4062 26380
rect 4120 26354 5120 26380
rect 5178 26354 6178 26380
rect 6236 26354 7236 26380
rect 8518 26370 9518 26388
rect 9576 26370 10576 26388
rect 10634 26370 11634 26388
rect 11692 26370 12692 26388
rect 12750 26370 13750 26388
rect 15024 26376 16024 26396
rect 16082 26376 17082 26396
rect 17140 26376 18140 26396
rect 18198 26376 19198 26396
rect 19256 26376 20256 26396
rect 47624 26406 48624 26424
rect 48682 26406 49682 26424
rect 49740 26406 50740 26424
rect 50798 26406 51798 26424
rect 51856 26406 52856 26424
rect 54138 26420 55138 26438
rect 55196 26420 56196 26438
rect 56254 26420 57254 26438
rect 57312 26420 58312 26438
rect 58370 26420 59370 26438
rect 54138 26412 59370 26420
rect 28036 26380 29036 26396
rect 29094 26380 30094 26396
rect 30152 26380 31152 26396
rect 31210 26380 32210 26396
rect 32268 26380 33268 26396
rect 15024 26370 20256 26376
rect 8518 26362 13750 26370
rect 2556 25988 2722 26354
rect 3280 25988 3446 26354
rect 4326 25988 4492 26354
rect 5356 25988 5522 26354
rect 6500 25988 6666 26354
rect 8940 26296 13550 26362
rect 11400 25996 11474 26296
rect 15458 26216 19886 26370
rect 21514 26362 22514 26380
rect 22572 26362 23572 26380
rect 23630 26362 24630 26380
rect 24688 26362 25688 26380
rect 25746 26362 26746 26380
rect 28036 26370 33268 26380
rect 34546 26384 35546 26402
rect 35604 26384 36604 26402
rect 36662 26384 37662 26402
rect 37720 26384 38720 26402
rect 38778 26384 39778 26402
rect 34546 26376 39778 26384
rect 41036 26382 42036 26402
rect 42094 26382 43094 26402
rect 43152 26382 44152 26402
rect 44210 26382 45210 26402
rect 45268 26382 46268 26402
rect 47624 26398 52856 26406
rect 41036 26376 46268 26382
rect 21514 26354 26746 26362
rect 17938 26004 18160 26216
rect 22130 26142 26428 26354
rect 28514 26168 32994 26370
rect 35006 26178 39496 26376
rect 41486 26214 45990 26376
rect 48048 26216 52548 26398
rect 2454 25946 7080 25988
rect 8968 25954 13594 25996
rect 15474 25962 20100 26004
rect 23230 25988 23528 26142
rect 30290 26004 30588 26168
rect 36860 26010 37222 26178
rect 43368 26010 43594 26214
rect 49306 26032 49532 26216
rect 54642 26196 59116 26412
rect 55622 26046 55848 26196
rect 15024 25956 20256 25962
rect 8518 25948 13750 25954
rect 2004 25940 7236 25946
rect 2004 25920 3004 25940
rect 3062 25920 4062 25940
rect 4120 25920 5120 25940
rect 5178 25920 6178 25940
rect 6236 25920 7236 25940
rect 8518 25928 9518 25948
rect 9576 25928 10576 25948
rect 10634 25928 11634 25948
rect 11692 25928 12692 25948
rect 12750 25928 13750 25948
rect 15024 25936 16024 25956
rect 16082 25936 17082 25956
rect 17140 25936 18140 25956
rect 18198 25936 19198 25956
rect 19256 25936 20256 25956
rect 21964 25946 26590 25988
rect 28486 25962 33112 26004
rect 34996 25968 39622 26010
rect 41486 25968 46112 26010
rect 48074 25990 52700 26032
rect 54588 26004 59214 26046
rect 54138 25998 59370 26004
rect 47624 25984 52856 25990
rect 34546 25962 39778 25968
rect 28036 25956 33268 25962
rect 21514 25940 26746 25946
rect 21514 25920 22514 25940
rect 22572 25920 23572 25940
rect 23630 25920 24630 25940
rect 24688 25920 25688 25940
rect 25746 25920 26746 25940
rect 28036 25936 29036 25956
rect 29094 25936 30094 25956
rect 30152 25936 31152 25956
rect 31210 25936 32210 25956
rect 32268 25936 33268 25956
rect 34546 25942 35546 25962
rect 35604 25942 36604 25962
rect 36662 25942 37662 25962
rect 37720 25942 38720 25962
rect 38778 25942 39778 25962
rect 41036 25962 46268 25968
rect 47624 25964 48624 25984
rect 48682 25964 49682 25984
rect 49740 25964 50740 25984
rect 50798 25964 51798 25984
rect 51856 25964 52856 25984
rect 54138 25978 55138 25998
rect 55196 25978 56196 25998
rect 56254 25978 57254 25998
rect 57312 25978 58312 25998
rect 58370 25978 59370 25998
rect 41036 25942 42036 25962
rect 42094 25942 43094 25962
rect 43152 25942 44152 25962
rect 44210 25942 45210 25962
rect 45268 25942 46268 25962
rect 2004 24894 3004 24920
rect 3062 24894 4062 24920
rect 4120 24894 5120 24920
rect 5178 24894 6178 24920
rect 6236 24894 7236 24920
rect 8518 24902 9518 24928
rect 9576 24902 10576 24928
rect 10634 24902 11634 24928
rect 11692 24902 12692 24928
rect 12750 24902 13750 24928
rect 15024 24910 16024 24936
rect 16082 24910 17082 24936
rect 17140 24910 18140 24936
rect 18198 24910 19198 24936
rect 19256 24910 20256 24936
rect 2256 24852 2790 24894
rect 3294 24852 3828 24894
rect 4412 24852 4946 24894
rect 5428 24852 5962 24894
rect 6494 24852 7028 24894
rect 8770 24860 9304 24902
rect 9808 24860 10342 24902
rect 10926 24860 11460 24902
rect 11942 24860 12476 24902
rect 13008 24860 13542 24902
rect 15276 24868 15810 24910
rect 16314 24868 16848 24910
rect 17432 24868 17966 24910
rect 18448 24868 18982 24910
rect 19514 24868 20048 24910
rect 21514 24894 22514 24920
rect 22572 24894 23572 24920
rect 23630 24894 24630 24920
rect 24688 24894 25688 24920
rect 25746 24894 26746 24920
rect 28036 24910 29036 24936
rect 29094 24910 30094 24936
rect 30152 24910 31152 24936
rect 31210 24910 32210 24936
rect 32268 24910 33268 24936
rect 34546 24916 35546 24942
rect 35604 24916 36604 24942
rect 36662 24916 37662 24942
rect 37720 24916 38720 24942
rect 38778 24916 39778 24942
rect 41036 24916 42036 24942
rect 42094 24916 43094 24942
rect 43152 24916 44152 24942
rect 44210 24916 45210 24942
rect 45268 24916 46268 24942
rect 47624 24938 48624 24964
rect 48682 24938 49682 24964
rect 49740 24938 50740 24964
rect 50798 24938 51798 24964
rect 51856 24938 52856 24964
rect 54138 24952 55138 24978
rect 55196 24952 56196 24978
rect 56254 24952 57254 24978
rect 57312 24952 58312 24978
rect 58370 24952 59370 24978
rect 2004 24826 3004 24852
rect 3062 24826 4062 24852
rect 4120 24826 5120 24852
rect 5178 24826 6178 24852
rect 6236 24826 7236 24852
rect 8518 24834 9518 24860
rect 9576 24834 10576 24860
rect 10634 24834 11634 24860
rect 11692 24834 12692 24860
rect 12750 24834 13750 24860
rect 15024 24842 16024 24868
rect 16082 24842 17082 24868
rect 17140 24842 18140 24868
rect 18198 24842 19198 24868
rect 19256 24842 20256 24868
rect 21766 24852 22300 24894
rect 22804 24852 23338 24894
rect 23922 24852 24456 24894
rect 24938 24852 25472 24894
rect 26004 24852 26538 24894
rect 28288 24868 28822 24910
rect 29326 24868 29860 24910
rect 30444 24868 30978 24910
rect 31460 24868 31994 24910
rect 32526 24868 33060 24910
rect 34798 24874 35332 24916
rect 35836 24874 36370 24916
rect 36954 24874 37488 24916
rect 37970 24874 38504 24916
rect 39036 24874 39570 24916
rect 41288 24874 41822 24916
rect 42326 24874 42860 24916
rect 43444 24874 43978 24916
rect 44460 24874 44994 24916
rect 45526 24874 46060 24916
rect 47876 24896 48410 24938
rect 48914 24896 49448 24938
rect 50032 24896 50566 24938
rect 51048 24896 51582 24938
rect 52114 24896 52648 24938
rect 54390 24910 54924 24952
rect 55428 24910 55962 24952
rect 56546 24910 57080 24952
rect 57562 24910 58096 24952
rect 58628 24910 59162 24952
rect 2004 23800 3004 23826
rect 3062 23800 4062 23826
rect 4120 23800 5120 23826
rect 5178 23800 6178 23826
rect 6236 23800 7236 23826
rect 2292 23758 2826 23800
rect 3248 23758 3782 23800
rect 4356 23758 4890 23800
rect 5462 23758 5996 23800
rect 6492 23758 7026 23800
rect 2004 23732 3004 23758
rect 3062 23732 4062 23758
rect 4120 23732 5120 23758
rect 5178 23732 6178 23758
rect 6236 23732 7236 23758
rect 8518 23808 9518 23834
rect 9576 23808 10576 23834
rect 10634 23808 11634 23834
rect 11692 23808 12692 23834
rect 12750 23808 13750 23834
rect 8806 23766 9340 23808
rect 9762 23766 10296 23808
rect 10870 23766 11404 23808
rect 11976 23766 12510 23808
rect 13006 23766 13540 23808
rect 8518 23740 9518 23766
rect 9576 23740 10576 23766
rect 10634 23740 11634 23766
rect 11692 23740 12692 23766
rect 12750 23740 13750 23766
rect 2004 22706 3004 22732
rect 3062 22706 4062 22732
rect 4120 22706 5120 22732
rect 5178 22706 6178 22732
rect 6236 22706 7236 22732
rect 2228 22664 2762 22706
rect 3282 22664 3816 22706
rect 4334 22664 4868 22706
rect 5442 22664 5976 22706
rect 6498 22664 7032 22706
rect 2004 22638 3004 22664
rect 3062 22638 4062 22664
rect 4120 22638 5120 22664
rect 5178 22638 6178 22664
rect 6236 22638 7236 22664
rect 21514 24826 22514 24852
rect 22572 24826 23572 24852
rect 23630 24826 24630 24852
rect 24688 24826 25688 24852
rect 25746 24826 26746 24852
rect 28036 24842 29036 24868
rect 29094 24842 30094 24868
rect 30152 24842 31152 24868
rect 31210 24842 32210 24868
rect 32268 24842 33268 24868
rect 34546 24848 35546 24874
rect 35604 24848 36604 24874
rect 36662 24848 37662 24874
rect 37720 24848 38720 24874
rect 38778 24848 39778 24874
rect 41036 24848 42036 24874
rect 42094 24848 43094 24874
rect 43152 24848 44152 24874
rect 44210 24848 45210 24874
rect 45268 24848 46268 24874
rect 47624 24870 48624 24896
rect 48682 24870 49682 24896
rect 49740 24870 50740 24896
rect 50798 24870 51798 24896
rect 51856 24870 52856 24896
rect 54138 24884 55138 24910
rect 55196 24884 56196 24910
rect 56254 24884 57254 24910
rect 57312 24884 58312 24910
rect 58370 24884 59370 24910
rect 15024 23816 16024 23842
rect 16082 23816 17082 23842
rect 17140 23816 18140 23842
rect 18198 23816 19198 23842
rect 19256 23816 20256 23842
rect 15312 23774 15846 23816
rect 16268 23774 16802 23816
rect 17376 23774 17910 23816
rect 18482 23774 19016 23816
rect 19512 23774 20046 23816
rect 15024 23748 16024 23774
rect 16082 23748 17082 23774
rect 17140 23748 18140 23774
rect 18198 23748 19198 23774
rect 19256 23748 20256 23774
rect 8518 22714 9518 22740
rect 9576 22714 10576 22740
rect 10634 22714 11634 22740
rect 11692 22714 12692 22740
rect 12750 22714 13750 22740
rect 8742 22672 9276 22714
rect 9796 22672 10330 22714
rect 10848 22672 11382 22714
rect 11956 22672 12490 22714
rect 13012 22672 13546 22714
rect 8518 22646 9518 22672
rect 9576 22646 10576 22672
rect 10634 22646 11634 22672
rect 11692 22646 12692 22672
rect 12750 22646 13750 22672
rect 21514 23800 22514 23826
rect 22572 23800 23572 23826
rect 23630 23800 24630 23826
rect 24688 23800 25688 23826
rect 25746 23800 26746 23826
rect 21802 23758 22336 23800
rect 22758 23758 23292 23800
rect 23866 23758 24400 23800
rect 24972 23758 25506 23800
rect 26002 23758 26536 23800
rect 21514 23732 22514 23758
rect 22572 23732 23572 23758
rect 23630 23732 24630 23758
rect 24688 23732 25688 23758
rect 25746 23732 26746 23758
rect 15024 22722 16024 22748
rect 16082 22722 17082 22748
rect 17140 22722 18140 22748
rect 18198 22722 19198 22748
rect 19256 22722 20256 22748
rect 15248 22680 15782 22722
rect 16302 22680 16836 22722
rect 17354 22680 17888 22722
rect 18462 22680 18996 22722
rect 19518 22680 20052 22722
rect 15024 22654 16024 22680
rect 16082 22654 17082 22680
rect 17140 22654 18140 22680
rect 18198 22654 19198 22680
rect 19256 22654 20256 22680
rect 28036 23816 29036 23842
rect 29094 23816 30094 23842
rect 30152 23816 31152 23842
rect 31210 23816 32210 23842
rect 32268 23816 33268 23842
rect 28324 23774 28858 23816
rect 29280 23774 29814 23816
rect 30388 23774 30922 23816
rect 31494 23774 32028 23816
rect 32524 23774 33058 23816
rect 28036 23748 29036 23774
rect 29094 23748 30094 23774
rect 30152 23748 31152 23774
rect 31210 23748 32210 23774
rect 32268 23748 33268 23774
rect 21514 22706 22514 22732
rect 22572 22706 23572 22732
rect 23630 22706 24630 22732
rect 24688 22706 25688 22732
rect 25746 22706 26746 22732
rect 21738 22664 22272 22706
rect 22792 22664 23326 22706
rect 23844 22664 24378 22706
rect 24952 22664 25486 22706
rect 26008 22664 26542 22706
rect 21514 22638 22514 22664
rect 22572 22638 23572 22664
rect 23630 22638 24630 22664
rect 24688 22638 25688 22664
rect 25746 22638 26746 22664
rect 2004 21612 3004 21638
rect 3062 21612 4062 21638
rect 4120 21612 5120 21638
rect 5178 21612 6178 21638
rect 6236 21612 7236 21638
rect 8518 21620 9518 21646
rect 9576 21620 10576 21646
rect 10634 21620 11634 21646
rect 11692 21620 12692 21646
rect 12750 21620 13750 21646
rect 15024 21628 16024 21654
rect 16082 21628 17082 21654
rect 17140 21628 18140 21654
rect 18198 21628 19198 21654
rect 19256 21628 20256 21654
rect 34546 23822 35546 23848
rect 35604 23822 36604 23848
rect 36662 23822 37662 23848
rect 37720 23822 38720 23848
rect 38778 23822 39778 23848
rect 34834 23780 35368 23822
rect 35790 23780 36324 23822
rect 36898 23780 37432 23822
rect 38004 23780 38538 23822
rect 39034 23780 39568 23822
rect 34546 23754 35546 23780
rect 35604 23754 36604 23780
rect 36662 23754 37662 23780
rect 37720 23754 38720 23780
rect 38778 23754 39778 23780
rect 28036 22722 29036 22748
rect 29094 22722 30094 22748
rect 30152 22722 31152 22748
rect 31210 22722 32210 22748
rect 32268 22722 33268 22748
rect 28260 22680 28794 22722
rect 29314 22680 29848 22722
rect 30366 22680 30900 22722
rect 31474 22680 32008 22722
rect 32530 22680 33064 22722
rect 28036 22654 29036 22680
rect 29094 22654 30094 22680
rect 30152 22654 31152 22680
rect 31210 22654 32210 22680
rect 32268 22654 33268 22680
rect 41036 23822 42036 23848
rect 42094 23822 43094 23848
rect 43152 23822 44152 23848
rect 44210 23822 45210 23848
rect 45268 23822 46268 23848
rect 41324 23780 41858 23822
rect 42280 23780 42814 23822
rect 43388 23780 43922 23822
rect 44494 23780 45028 23822
rect 45524 23780 46058 23822
rect 41036 23754 42036 23780
rect 42094 23754 43094 23780
rect 43152 23754 44152 23780
rect 44210 23754 45210 23780
rect 45268 23754 46268 23780
rect 34546 22728 35546 22754
rect 35604 22728 36604 22754
rect 36662 22728 37662 22754
rect 37720 22728 38720 22754
rect 38778 22728 39778 22754
rect 34770 22686 35304 22728
rect 35824 22686 36358 22728
rect 36876 22686 37410 22728
rect 37984 22686 38518 22728
rect 39040 22686 39574 22728
rect 34546 22660 35546 22686
rect 35604 22660 36604 22686
rect 36662 22660 37662 22686
rect 37720 22660 38720 22686
rect 38778 22660 39778 22686
rect 47624 23844 48624 23870
rect 48682 23844 49682 23870
rect 49740 23844 50740 23870
rect 50798 23844 51798 23870
rect 51856 23844 52856 23870
rect 47912 23802 48446 23844
rect 48868 23802 49402 23844
rect 49976 23802 50510 23844
rect 51082 23802 51616 23844
rect 52112 23802 52646 23844
rect 47624 23776 48624 23802
rect 48682 23776 49682 23802
rect 49740 23776 50740 23802
rect 50798 23776 51798 23802
rect 51856 23776 52856 23802
rect 41036 22728 42036 22754
rect 42094 22728 43094 22754
rect 43152 22728 44152 22754
rect 44210 22728 45210 22754
rect 45268 22728 46268 22754
rect 41260 22686 41794 22728
rect 42314 22686 42848 22728
rect 43366 22686 43900 22728
rect 44474 22686 45008 22728
rect 45530 22686 46064 22728
rect 41036 22660 42036 22686
rect 42094 22660 43094 22686
rect 43152 22660 44152 22686
rect 44210 22660 45210 22686
rect 45268 22660 46268 22686
rect 54138 23858 55138 23884
rect 55196 23858 56196 23884
rect 56254 23858 57254 23884
rect 57312 23858 58312 23884
rect 58370 23858 59370 23884
rect 54426 23816 54960 23858
rect 55382 23816 55916 23858
rect 56490 23816 57024 23858
rect 57596 23816 58130 23858
rect 58626 23816 59160 23858
rect 54138 23790 55138 23816
rect 55196 23790 56196 23816
rect 56254 23790 57254 23816
rect 57312 23790 58312 23816
rect 58370 23790 59370 23816
rect 47624 22750 48624 22776
rect 48682 22750 49682 22776
rect 49740 22750 50740 22776
rect 50798 22750 51798 22776
rect 51856 22750 52856 22776
rect 47848 22708 48382 22750
rect 48902 22708 49436 22750
rect 49954 22708 50488 22750
rect 51062 22708 51596 22750
rect 52118 22708 52652 22750
rect 47624 22682 48624 22708
rect 48682 22682 49682 22708
rect 49740 22682 50740 22708
rect 50798 22682 51798 22708
rect 51856 22682 52856 22708
rect 54138 22764 55138 22790
rect 55196 22764 56196 22790
rect 56254 22764 57254 22790
rect 57312 22764 58312 22790
rect 58370 22764 59370 22790
rect 54362 22722 54896 22764
rect 55416 22722 55950 22764
rect 56468 22722 57002 22764
rect 57576 22722 58110 22764
rect 58632 22722 59166 22764
rect 54138 22696 55138 22722
rect 55196 22696 56196 22722
rect 56254 22696 57254 22722
rect 57312 22696 58312 22722
rect 58370 22696 59370 22722
rect 2256 21570 2790 21612
rect 3354 21570 3888 21612
rect 4382 21570 4916 21612
rect 5346 21570 5880 21612
rect 6446 21570 6980 21612
rect 8770 21578 9304 21620
rect 9868 21578 10402 21620
rect 10896 21578 11430 21620
rect 11860 21578 12394 21620
rect 12960 21578 13494 21620
rect 15276 21586 15810 21628
rect 16374 21586 16908 21628
rect 17402 21586 17936 21628
rect 18366 21586 18900 21628
rect 19466 21586 20000 21628
rect 21514 21612 22514 21638
rect 22572 21612 23572 21638
rect 23630 21612 24630 21638
rect 24688 21612 25688 21638
rect 25746 21612 26746 21638
rect 28036 21628 29036 21654
rect 29094 21628 30094 21654
rect 30152 21628 31152 21654
rect 31210 21628 32210 21654
rect 32268 21628 33268 21654
rect 34546 21634 35546 21660
rect 35604 21634 36604 21660
rect 36662 21634 37662 21660
rect 37720 21634 38720 21660
rect 38778 21634 39778 21660
rect 41036 21634 42036 21660
rect 42094 21634 43094 21660
rect 43152 21634 44152 21660
rect 44210 21634 45210 21660
rect 45268 21634 46268 21660
rect 47624 21656 48624 21682
rect 48682 21656 49682 21682
rect 49740 21656 50740 21682
rect 50798 21656 51798 21682
rect 51856 21656 52856 21682
rect 54138 21670 55138 21696
rect 55196 21670 56196 21696
rect 56254 21670 57254 21696
rect 57312 21670 58312 21696
rect 58370 21670 59370 21696
rect 2004 21544 3004 21570
rect 3062 21544 4062 21570
rect 4120 21544 5120 21570
rect 5178 21544 6178 21570
rect 6236 21544 7236 21570
rect 8518 21552 9518 21578
rect 9576 21552 10576 21578
rect 10634 21552 11634 21578
rect 11692 21552 12692 21578
rect 12750 21552 13750 21578
rect 15024 21560 16024 21586
rect 16082 21560 17082 21586
rect 17140 21560 18140 21586
rect 18198 21560 19198 21586
rect 19256 21560 20256 21586
rect 21766 21570 22300 21612
rect 22864 21570 23398 21612
rect 23892 21570 24426 21612
rect 24856 21570 25390 21612
rect 25956 21570 26490 21612
rect 28288 21586 28822 21628
rect 29386 21586 29920 21628
rect 30414 21586 30948 21628
rect 31378 21586 31912 21628
rect 32478 21586 33012 21628
rect 34798 21592 35332 21634
rect 35896 21592 36430 21634
rect 36924 21592 37458 21634
rect 37888 21592 38422 21634
rect 38988 21592 39522 21634
rect 41288 21592 41822 21634
rect 42386 21592 42920 21634
rect 43414 21592 43948 21634
rect 44378 21592 44912 21634
rect 45478 21592 46012 21634
rect 47876 21614 48410 21656
rect 48974 21614 49508 21656
rect 50002 21614 50536 21656
rect 50966 21614 51500 21656
rect 52066 21614 52600 21656
rect 54390 21628 54924 21670
rect 55488 21628 56022 21670
rect 56516 21628 57050 21670
rect 57480 21628 58014 21670
rect 58580 21628 59114 21670
rect 21514 21544 22514 21570
rect 22572 21544 23572 21570
rect 23630 21544 24630 21570
rect 24688 21544 25688 21570
rect 25746 21544 26746 21570
rect 28036 21560 29036 21586
rect 29094 21560 30094 21586
rect 30152 21560 31152 21586
rect 31210 21560 32210 21586
rect 32268 21560 33268 21586
rect 34546 21566 35546 21592
rect 35604 21566 36604 21592
rect 36662 21566 37662 21592
rect 37720 21566 38720 21592
rect 38778 21566 39778 21592
rect 41036 21566 42036 21592
rect 42094 21566 43094 21592
rect 43152 21566 44152 21592
rect 44210 21566 45210 21592
rect 45268 21566 46268 21592
rect 47624 21588 48624 21614
rect 48682 21588 49682 21614
rect 49740 21588 50740 21614
rect 50798 21588 51798 21614
rect 51856 21588 52856 21614
rect 54138 21602 55138 21628
rect 55196 21602 56196 21628
rect 56254 21602 57254 21628
rect 57312 21602 58312 21628
rect 58370 21602 59370 21628
rect 2004 20518 3004 20544
rect 3062 20518 4062 20544
rect 4120 20518 5120 20544
rect 5178 20518 6178 20544
rect 6236 20518 7236 20544
rect 8518 20534 9518 20552
rect 9576 20534 10576 20552
rect 10634 20534 11634 20552
rect 11692 20534 12692 20552
rect 12750 20534 13750 20552
rect 15024 20542 16024 20560
rect 16082 20542 17082 20560
rect 17140 20542 18140 20560
rect 18198 20542 19198 20560
rect 19256 20542 20256 20560
rect 47624 20572 48624 20588
rect 48682 20572 49682 20588
rect 49740 20572 50740 20588
rect 50798 20572 51798 20588
rect 51856 20572 52856 20588
rect 54138 20582 55138 20602
rect 55196 20582 56196 20602
rect 56254 20582 57254 20602
rect 57312 20582 58312 20602
rect 58370 20582 59370 20602
rect 54138 20576 59370 20582
rect 15024 20534 20256 20542
rect 8518 20526 13750 20534
rect 2598 20124 2814 20518
rect 3366 20124 3582 20518
rect 4412 20124 4628 20518
rect 5450 20124 5666 20518
rect 6390 20124 6606 20518
rect 8948 20486 13634 20526
rect 11048 20132 11228 20486
rect 15464 20322 19726 20534
rect 21514 20528 22514 20544
rect 22572 20528 23572 20544
rect 23630 20528 24630 20544
rect 24688 20528 25688 20544
rect 25746 20528 26746 20544
rect 28036 20538 29036 20560
rect 29094 20538 30094 20560
rect 30152 20538 31152 20560
rect 31210 20538 32210 20560
rect 32268 20538 33268 20560
rect 34546 20546 35546 20566
rect 35604 20546 36604 20566
rect 36662 20546 37662 20566
rect 37720 20546 38720 20566
rect 38778 20546 39778 20566
rect 34546 20540 39778 20546
rect 41036 20550 42036 20566
rect 42094 20550 43094 20566
rect 43152 20550 44152 20566
rect 44210 20550 45210 20566
rect 45268 20550 46268 20566
rect 47624 20562 52856 20572
rect 41036 20540 46268 20550
rect 28036 20534 33268 20538
rect 21514 20518 26746 20528
rect 17880 20140 18024 20322
rect 21998 20302 26298 20518
rect 28398 20338 32876 20534
rect 34948 20340 39438 20540
rect 41482 20354 45982 20540
rect 47950 20382 52450 20562
rect 2454 20082 7080 20124
rect 8968 20090 13594 20132
rect 15474 20098 20100 20140
rect 23112 20124 23318 20302
rect 30426 20140 30632 20338
rect 36984 20146 37190 20340
rect 43400 20146 43626 20354
rect 49328 20168 49554 20382
rect 54558 20358 59032 20576
rect 55654 20182 55880 20358
rect 15024 20092 20256 20098
rect 8518 20084 13750 20090
rect 2004 20076 7236 20082
rect 2004 20056 3004 20076
rect 3062 20056 4062 20076
rect 4120 20056 5120 20076
rect 5178 20056 6178 20076
rect 6236 20056 7236 20076
rect 8518 20064 9518 20084
rect 9576 20064 10576 20084
rect 10634 20064 11634 20084
rect 11692 20064 12692 20084
rect 12750 20064 13750 20084
rect 15024 20072 16024 20092
rect 16082 20072 17082 20092
rect 17140 20072 18140 20092
rect 18198 20072 19198 20092
rect 19256 20072 20256 20092
rect 21964 20082 26590 20124
rect 28486 20098 33112 20140
rect 34996 20104 39622 20146
rect 41486 20104 46112 20146
rect 48074 20126 52700 20168
rect 54588 20140 59214 20182
rect 54138 20134 59370 20140
rect 47624 20120 52856 20126
rect 34546 20098 39778 20104
rect 28036 20092 33268 20098
rect 21514 20076 26746 20082
rect 21514 20056 22514 20076
rect 22572 20056 23572 20076
rect 23630 20056 24630 20076
rect 24688 20056 25688 20076
rect 25746 20056 26746 20076
rect 28036 20072 29036 20092
rect 29094 20072 30094 20092
rect 30152 20072 31152 20092
rect 31210 20072 32210 20092
rect 32268 20072 33268 20092
rect 34546 20078 35546 20098
rect 35604 20078 36604 20098
rect 36662 20078 37662 20098
rect 37720 20078 38720 20098
rect 38778 20078 39778 20098
rect 41036 20098 46268 20104
rect 47624 20100 48624 20120
rect 48682 20100 49682 20120
rect 49740 20100 50740 20120
rect 50798 20100 51798 20120
rect 51856 20100 52856 20120
rect 54138 20114 55138 20134
rect 55196 20114 56196 20134
rect 56254 20114 57254 20134
rect 57312 20114 58312 20134
rect 58370 20114 59370 20134
rect 41036 20078 42036 20098
rect 42094 20078 43094 20098
rect 43152 20078 44152 20098
rect 44210 20078 45210 20098
rect 45268 20078 46268 20098
rect 2004 19030 3004 19056
rect 3062 19030 4062 19056
rect 4120 19030 5120 19056
rect 5178 19030 6178 19056
rect 6236 19030 7236 19056
rect 8518 19038 9518 19064
rect 9576 19038 10576 19064
rect 10634 19038 11634 19064
rect 11692 19038 12692 19064
rect 12750 19038 13750 19064
rect 15024 19046 16024 19072
rect 16082 19046 17082 19072
rect 17140 19046 18140 19072
rect 18198 19046 19198 19072
rect 19256 19046 20256 19072
rect 2256 18988 2790 19030
rect 3294 18988 3828 19030
rect 4412 18988 4946 19030
rect 5428 18988 5962 19030
rect 6494 18988 7028 19030
rect 8770 18996 9304 19038
rect 9808 18996 10342 19038
rect 10926 18996 11460 19038
rect 11942 18996 12476 19038
rect 13008 18996 13542 19038
rect 15276 19004 15810 19046
rect 16314 19004 16848 19046
rect 17432 19004 17966 19046
rect 18448 19004 18982 19046
rect 19514 19004 20048 19046
rect 21514 19030 22514 19056
rect 22572 19030 23572 19056
rect 23630 19030 24630 19056
rect 24688 19030 25688 19056
rect 25746 19030 26746 19056
rect 28036 19046 29036 19072
rect 29094 19046 30094 19072
rect 30152 19046 31152 19072
rect 31210 19046 32210 19072
rect 32268 19046 33268 19072
rect 34546 19052 35546 19078
rect 35604 19052 36604 19078
rect 36662 19052 37662 19078
rect 37720 19052 38720 19078
rect 38778 19052 39778 19078
rect 41036 19052 42036 19078
rect 42094 19052 43094 19078
rect 43152 19052 44152 19078
rect 44210 19052 45210 19078
rect 45268 19052 46268 19078
rect 47624 19074 48624 19100
rect 48682 19074 49682 19100
rect 49740 19074 50740 19100
rect 50798 19074 51798 19100
rect 51856 19074 52856 19100
rect 54138 19088 55138 19114
rect 55196 19088 56196 19114
rect 56254 19088 57254 19114
rect 57312 19088 58312 19114
rect 58370 19088 59370 19114
rect 2004 18962 3004 18988
rect 3062 18962 4062 18988
rect 4120 18962 5120 18988
rect 5178 18962 6178 18988
rect 6236 18962 7236 18988
rect 8518 18970 9518 18996
rect 9576 18970 10576 18996
rect 10634 18970 11634 18996
rect 11692 18970 12692 18996
rect 12750 18970 13750 18996
rect 15024 18978 16024 19004
rect 16082 18978 17082 19004
rect 17140 18978 18140 19004
rect 18198 18978 19198 19004
rect 19256 18978 20256 19004
rect 21766 18988 22300 19030
rect 22804 18988 23338 19030
rect 23922 18988 24456 19030
rect 24938 18988 25472 19030
rect 26004 18988 26538 19030
rect 28288 19004 28822 19046
rect 29326 19004 29860 19046
rect 30444 19004 30978 19046
rect 31460 19004 31994 19046
rect 32526 19004 33060 19046
rect 34798 19010 35332 19052
rect 35836 19010 36370 19052
rect 36954 19010 37488 19052
rect 37970 19010 38504 19052
rect 39036 19010 39570 19052
rect 41288 19010 41822 19052
rect 42326 19010 42860 19052
rect 43444 19010 43978 19052
rect 44460 19010 44994 19052
rect 45526 19010 46060 19052
rect 47876 19032 48410 19074
rect 48914 19032 49448 19074
rect 50032 19032 50566 19074
rect 51048 19032 51582 19074
rect 52114 19032 52648 19074
rect 54390 19046 54924 19088
rect 55428 19046 55962 19088
rect 56546 19046 57080 19088
rect 57562 19046 58096 19088
rect 58628 19046 59162 19088
rect 2004 17936 3004 17962
rect 3062 17936 4062 17962
rect 4120 17936 5120 17962
rect 5178 17936 6178 17962
rect 6236 17936 7236 17962
rect 2292 17894 2826 17936
rect 3248 17894 3782 17936
rect 4356 17894 4890 17936
rect 5462 17894 5996 17936
rect 6492 17894 7026 17936
rect 2004 17868 3004 17894
rect 3062 17868 4062 17894
rect 4120 17868 5120 17894
rect 5178 17868 6178 17894
rect 6236 17868 7236 17894
rect 8518 17944 9518 17970
rect 9576 17944 10576 17970
rect 10634 17944 11634 17970
rect 11692 17944 12692 17970
rect 12750 17944 13750 17970
rect 8806 17902 9340 17944
rect 9762 17902 10296 17944
rect 10870 17902 11404 17944
rect 11976 17902 12510 17944
rect 13006 17902 13540 17944
rect 8518 17876 9518 17902
rect 9576 17876 10576 17902
rect 10634 17876 11634 17902
rect 11692 17876 12692 17902
rect 12750 17876 13750 17902
rect 2004 16842 3004 16868
rect 3062 16842 4062 16868
rect 4120 16842 5120 16868
rect 5178 16842 6178 16868
rect 6236 16842 7236 16868
rect 2228 16800 2762 16842
rect 3282 16800 3816 16842
rect 4334 16800 4868 16842
rect 5442 16800 5976 16842
rect 6498 16800 7032 16842
rect 2004 16774 3004 16800
rect 3062 16774 4062 16800
rect 4120 16774 5120 16800
rect 5178 16774 6178 16800
rect 6236 16774 7236 16800
rect 21514 18962 22514 18988
rect 22572 18962 23572 18988
rect 23630 18962 24630 18988
rect 24688 18962 25688 18988
rect 25746 18962 26746 18988
rect 28036 18978 29036 19004
rect 29094 18978 30094 19004
rect 30152 18978 31152 19004
rect 31210 18978 32210 19004
rect 32268 18978 33268 19004
rect 34546 18984 35546 19010
rect 35604 18984 36604 19010
rect 36662 18984 37662 19010
rect 37720 18984 38720 19010
rect 38778 18984 39778 19010
rect 41036 18984 42036 19010
rect 42094 18984 43094 19010
rect 43152 18984 44152 19010
rect 44210 18984 45210 19010
rect 45268 18984 46268 19010
rect 47624 19006 48624 19032
rect 48682 19006 49682 19032
rect 49740 19006 50740 19032
rect 50798 19006 51798 19032
rect 51856 19006 52856 19032
rect 54138 19020 55138 19046
rect 55196 19020 56196 19046
rect 56254 19020 57254 19046
rect 57312 19020 58312 19046
rect 58370 19020 59370 19046
rect 15024 17952 16024 17978
rect 16082 17952 17082 17978
rect 17140 17952 18140 17978
rect 18198 17952 19198 17978
rect 19256 17952 20256 17978
rect 15312 17910 15846 17952
rect 16268 17910 16802 17952
rect 17376 17910 17910 17952
rect 18482 17910 19016 17952
rect 19512 17910 20046 17952
rect 15024 17884 16024 17910
rect 16082 17884 17082 17910
rect 17140 17884 18140 17910
rect 18198 17884 19198 17910
rect 19256 17884 20256 17910
rect 8518 16850 9518 16876
rect 9576 16850 10576 16876
rect 10634 16850 11634 16876
rect 11692 16850 12692 16876
rect 12750 16850 13750 16876
rect 8742 16808 9276 16850
rect 9796 16808 10330 16850
rect 10848 16808 11382 16850
rect 11956 16808 12490 16850
rect 13012 16808 13546 16850
rect 8518 16782 9518 16808
rect 9576 16782 10576 16808
rect 10634 16782 11634 16808
rect 11692 16782 12692 16808
rect 12750 16782 13750 16808
rect 21514 17936 22514 17962
rect 22572 17936 23572 17962
rect 23630 17936 24630 17962
rect 24688 17936 25688 17962
rect 25746 17936 26746 17962
rect 21802 17894 22336 17936
rect 22758 17894 23292 17936
rect 23866 17894 24400 17936
rect 24972 17894 25506 17936
rect 26002 17894 26536 17936
rect 21514 17868 22514 17894
rect 22572 17868 23572 17894
rect 23630 17868 24630 17894
rect 24688 17868 25688 17894
rect 25746 17868 26746 17894
rect 15024 16858 16024 16884
rect 16082 16858 17082 16884
rect 17140 16858 18140 16884
rect 18198 16858 19198 16884
rect 19256 16858 20256 16884
rect 15248 16816 15782 16858
rect 16302 16816 16836 16858
rect 17354 16816 17888 16858
rect 18462 16816 18996 16858
rect 19518 16816 20052 16858
rect 15024 16790 16024 16816
rect 16082 16790 17082 16816
rect 17140 16790 18140 16816
rect 18198 16790 19198 16816
rect 19256 16790 20256 16816
rect 28036 17952 29036 17978
rect 29094 17952 30094 17978
rect 30152 17952 31152 17978
rect 31210 17952 32210 17978
rect 32268 17952 33268 17978
rect 28324 17910 28858 17952
rect 29280 17910 29814 17952
rect 30388 17910 30922 17952
rect 31494 17910 32028 17952
rect 32524 17910 33058 17952
rect 28036 17884 29036 17910
rect 29094 17884 30094 17910
rect 30152 17884 31152 17910
rect 31210 17884 32210 17910
rect 32268 17884 33268 17910
rect 21514 16842 22514 16868
rect 22572 16842 23572 16868
rect 23630 16842 24630 16868
rect 24688 16842 25688 16868
rect 25746 16842 26746 16868
rect 21738 16800 22272 16842
rect 22792 16800 23326 16842
rect 23844 16800 24378 16842
rect 24952 16800 25486 16842
rect 26008 16800 26542 16842
rect 21514 16774 22514 16800
rect 22572 16774 23572 16800
rect 23630 16774 24630 16800
rect 24688 16774 25688 16800
rect 25746 16774 26746 16800
rect 2004 15748 3004 15774
rect 3062 15748 4062 15774
rect 4120 15748 5120 15774
rect 5178 15748 6178 15774
rect 6236 15748 7236 15774
rect 8518 15756 9518 15782
rect 9576 15756 10576 15782
rect 10634 15756 11634 15782
rect 11692 15756 12692 15782
rect 12750 15756 13750 15782
rect 15024 15764 16024 15790
rect 16082 15764 17082 15790
rect 17140 15764 18140 15790
rect 18198 15764 19198 15790
rect 19256 15764 20256 15790
rect 34546 17958 35546 17984
rect 35604 17958 36604 17984
rect 36662 17958 37662 17984
rect 37720 17958 38720 17984
rect 38778 17958 39778 17984
rect 34834 17916 35368 17958
rect 35790 17916 36324 17958
rect 36898 17916 37432 17958
rect 38004 17916 38538 17958
rect 39034 17916 39568 17958
rect 34546 17890 35546 17916
rect 35604 17890 36604 17916
rect 36662 17890 37662 17916
rect 37720 17890 38720 17916
rect 38778 17890 39778 17916
rect 28036 16858 29036 16884
rect 29094 16858 30094 16884
rect 30152 16858 31152 16884
rect 31210 16858 32210 16884
rect 32268 16858 33268 16884
rect 28260 16816 28794 16858
rect 29314 16816 29848 16858
rect 30366 16816 30900 16858
rect 31474 16816 32008 16858
rect 32530 16816 33064 16858
rect 28036 16790 29036 16816
rect 29094 16790 30094 16816
rect 30152 16790 31152 16816
rect 31210 16790 32210 16816
rect 32268 16790 33268 16816
rect 41036 17958 42036 17984
rect 42094 17958 43094 17984
rect 43152 17958 44152 17984
rect 44210 17958 45210 17984
rect 45268 17958 46268 17984
rect 41324 17916 41858 17958
rect 42280 17916 42814 17958
rect 43388 17916 43922 17958
rect 44494 17916 45028 17958
rect 45524 17916 46058 17958
rect 41036 17890 42036 17916
rect 42094 17890 43094 17916
rect 43152 17890 44152 17916
rect 44210 17890 45210 17916
rect 45268 17890 46268 17916
rect 34546 16864 35546 16890
rect 35604 16864 36604 16890
rect 36662 16864 37662 16890
rect 37720 16864 38720 16890
rect 38778 16864 39778 16890
rect 34770 16822 35304 16864
rect 35824 16822 36358 16864
rect 36876 16822 37410 16864
rect 37984 16822 38518 16864
rect 39040 16822 39574 16864
rect 34546 16796 35546 16822
rect 35604 16796 36604 16822
rect 36662 16796 37662 16822
rect 37720 16796 38720 16822
rect 38778 16796 39778 16822
rect 47624 17980 48624 18006
rect 48682 17980 49682 18006
rect 49740 17980 50740 18006
rect 50798 17980 51798 18006
rect 51856 17980 52856 18006
rect 47912 17938 48446 17980
rect 48868 17938 49402 17980
rect 49976 17938 50510 17980
rect 51082 17938 51616 17980
rect 52112 17938 52646 17980
rect 47624 17912 48624 17938
rect 48682 17912 49682 17938
rect 49740 17912 50740 17938
rect 50798 17912 51798 17938
rect 51856 17912 52856 17938
rect 41036 16864 42036 16890
rect 42094 16864 43094 16890
rect 43152 16864 44152 16890
rect 44210 16864 45210 16890
rect 45268 16864 46268 16890
rect 41260 16822 41794 16864
rect 42314 16822 42848 16864
rect 43366 16822 43900 16864
rect 44474 16822 45008 16864
rect 45530 16822 46064 16864
rect 41036 16796 42036 16822
rect 42094 16796 43094 16822
rect 43152 16796 44152 16822
rect 44210 16796 45210 16822
rect 45268 16796 46268 16822
rect 54138 17994 55138 18020
rect 55196 17994 56196 18020
rect 56254 17994 57254 18020
rect 57312 17994 58312 18020
rect 58370 17994 59370 18020
rect 54426 17952 54960 17994
rect 55382 17952 55916 17994
rect 56490 17952 57024 17994
rect 57596 17952 58130 17994
rect 58626 17952 59160 17994
rect 54138 17926 55138 17952
rect 55196 17926 56196 17952
rect 56254 17926 57254 17952
rect 57312 17926 58312 17952
rect 58370 17926 59370 17952
rect 47624 16886 48624 16912
rect 48682 16886 49682 16912
rect 49740 16886 50740 16912
rect 50798 16886 51798 16912
rect 51856 16886 52856 16912
rect 47848 16844 48382 16886
rect 48902 16844 49436 16886
rect 49954 16844 50488 16886
rect 51062 16844 51596 16886
rect 52118 16844 52652 16886
rect 47624 16818 48624 16844
rect 48682 16818 49682 16844
rect 49740 16818 50740 16844
rect 50798 16818 51798 16844
rect 51856 16818 52856 16844
rect 54138 16900 55138 16926
rect 55196 16900 56196 16926
rect 56254 16900 57254 16926
rect 57312 16900 58312 16926
rect 58370 16900 59370 16926
rect 54362 16858 54896 16900
rect 55416 16858 55950 16900
rect 56468 16858 57002 16900
rect 57576 16858 58110 16900
rect 58632 16858 59166 16900
rect 54138 16832 55138 16858
rect 55196 16832 56196 16858
rect 56254 16832 57254 16858
rect 57312 16832 58312 16858
rect 58370 16832 59370 16858
rect 2256 15706 2790 15748
rect 3354 15706 3888 15748
rect 4382 15706 4916 15748
rect 5346 15706 5880 15748
rect 6446 15706 6980 15748
rect 8770 15714 9304 15756
rect 9868 15714 10402 15756
rect 10896 15714 11430 15756
rect 11860 15714 12394 15756
rect 12960 15714 13494 15756
rect 15276 15722 15810 15764
rect 16374 15722 16908 15764
rect 17402 15722 17936 15764
rect 18366 15722 18900 15764
rect 19466 15722 20000 15764
rect 21514 15748 22514 15774
rect 22572 15748 23572 15774
rect 23630 15748 24630 15774
rect 24688 15748 25688 15774
rect 25746 15748 26746 15774
rect 28036 15764 29036 15790
rect 29094 15764 30094 15790
rect 30152 15764 31152 15790
rect 31210 15764 32210 15790
rect 32268 15764 33268 15790
rect 34546 15770 35546 15796
rect 35604 15770 36604 15796
rect 36662 15770 37662 15796
rect 37720 15770 38720 15796
rect 38778 15770 39778 15796
rect 41036 15770 42036 15796
rect 42094 15770 43094 15796
rect 43152 15770 44152 15796
rect 44210 15770 45210 15796
rect 45268 15770 46268 15796
rect 47624 15792 48624 15818
rect 48682 15792 49682 15818
rect 49740 15792 50740 15818
rect 50798 15792 51798 15818
rect 51856 15792 52856 15818
rect 54138 15806 55138 15832
rect 55196 15806 56196 15832
rect 56254 15806 57254 15832
rect 57312 15806 58312 15832
rect 58370 15806 59370 15832
rect 2004 15680 3004 15706
rect 3062 15680 4062 15706
rect 4120 15680 5120 15706
rect 5178 15680 6178 15706
rect 6236 15680 7236 15706
rect 8518 15688 9518 15714
rect 9576 15688 10576 15714
rect 10634 15688 11634 15714
rect 11692 15688 12692 15714
rect 12750 15688 13750 15714
rect 15024 15696 16024 15722
rect 16082 15696 17082 15722
rect 17140 15696 18140 15722
rect 18198 15696 19198 15722
rect 19256 15696 20256 15722
rect 21766 15706 22300 15748
rect 22864 15706 23398 15748
rect 23892 15706 24426 15748
rect 24856 15706 25390 15748
rect 25956 15706 26490 15748
rect 28288 15722 28822 15764
rect 29386 15722 29920 15764
rect 30414 15722 30948 15764
rect 31378 15722 31912 15764
rect 32478 15722 33012 15764
rect 34798 15728 35332 15770
rect 35896 15728 36430 15770
rect 36924 15728 37458 15770
rect 37888 15728 38422 15770
rect 38988 15728 39522 15770
rect 41288 15728 41822 15770
rect 42386 15728 42920 15770
rect 43414 15728 43948 15770
rect 44378 15728 44912 15770
rect 45478 15728 46012 15770
rect 47876 15750 48410 15792
rect 48974 15750 49508 15792
rect 50002 15750 50536 15792
rect 50966 15750 51500 15792
rect 52066 15750 52600 15792
rect 54390 15764 54924 15806
rect 55488 15764 56022 15806
rect 56516 15764 57050 15806
rect 57480 15764 58014 15806
rect 58580 15764 59114 15806
rect 21514 15680 22514 15706
rect 22572 15680 23572 15706
rect 23630 15680 24630 15706
rect 24688 15680 25688 15706
rect 25746 15680 26746 15706
rect 28036 15696 29036 15722
rect 29094 15696 30094 15722
rect 30152 15696 31152 15722
rect 31210 15696 32210 15722
rect 32268 15696 33268 15722
rect 34546 15702 35546 15728
rect 35604 15702 36604 15728
rect 36662 15702 37662 15728
rect 37720 15702 38720 15728
rect 38778 15702 39778 15728
rect 41036 15702 42036 15728
rect 42094 15702 43094 15728
rect 43152 15702 44152 15728
rect 44210 15702 45210 15728
rect 45268 15702 46268 15728
rect 47624 15724 48624 15750
rect 48682 15724 49682 15750
rect 49740 15724 50740 15750
rect 50798 15724 51798 15750
rect 51856 15724 52856 15750
rect 54138 15738 55138 15764
rect 55196 15738 56196 15764
rect 56254 15738 57254 15764
rect 57312 15738 58312 15764
rect 58370 15738 59370 15764
rect 2004 14654 3004 14680
rect 3062 14654 4062 14680
rect 4120 14654 5120 14680
rect 5178 14654 6178 14680
rect 6236 14654 7236 14680
rect 8518 14670 9518 14688
rect 9576 14670 10576 14688
rect 10634 14670 11634 14688
rect 11692 14670 12692 14688
rect 12750 14670 13750 14688
rect 15024 14680 16024 14696
rect 16082 14680 17082 14696
rect 17140 14680 18140 14696
rect 18198 14680 19198 14696
rect 19256 14680 20256 14696
rect 47624 14706 48624 14724
rect 48682 14706 49682 14724
rect 49740 14706 50740 14724
rect 50798 14706 51798 14724
rect 51856 14706 52856 14724
rect 54138 14722 55138 14738
rect 55196 14722 56196 14738
rect 56254 14722 57254 14738
rect 57312 14722 58312 14738
rect 58370 14722 59370 14738
rect 54138 14712 59370 14722
rect 28036 14680 29036 14696
rect 29094 14680 30094 14696
rect 30152 14680 31152 14696
rect 31210 14680 32210 14696
rect 32268 14680 33268 14696
rect 15024 14670 20256 14680
rect 8518 14662 13750 14670
rect 2568 14268 2784 14654
rect 3336 14268 3552 14654
rect 4378 14268 4594 14654
rect 5428 14268 5644 14654
rect 6548 14268 6764 14654
rect 8958 14576 13514 14662
rect 11074 14276 11254 14576
rect 15500 14514 19968 14670
rect 21514 14662 22514 14680
rect 22572 14662 23572 14680
rect 23630 14662 24630 14680
rect 24688 14662 25688 14680
rect 25746 14662 26746 14680
rect 28036 14670 33268 14680
rect 34546 14682 35546 14702
rect 35604 14682 36604 14702
rect 36662 14682 37662 14702
rect 37720 14682 38720 14702
rect 38778 14682 39778 14702
rect 34546 14676 39778 14682
rect 41036 14684 42036 14702
rect 42094 14684 43094 14702
rect 43152 14684 44152 14702
rect 44210 14684 45210 14702
rect 45268 14684 46268 14702
rect 47624 14698 52856 14706
rect 41036 14676 46268 14684
rect 21514 14654 26746 14662
rect 17714 14284 17882 14514
rect 21952 14436 26252 14654
rect 28578 14464 32868 14670
rect 35006 14472 39498 14676
rect 2464 14226 7090 14268
rect 8978 14234 13604 14276
rect 15484 14242 20110 14284
rect 23042 14268 23248 14436
rect 30500 14284 30706 14464
rect 36942 14290 37148 14472
rect 41474 14468 45972 14676
rect 48102 14510 52578 14698
rect 43410 14290 43636 14468
rect 49994 14312 50220 14510
rect 54586 14498 59060 14712
rect 55612 14326 55838 14498
rect 15034 14236 20266 14242
rect 8528 14228 13760 14234
rect 2014 14220 7246 14226
rect 2014 14200 3014 14220
rect 3072 14200 4072 14220
rect 4130 14200 5130 14220
rect 5188 14200 6188 14220
rect 6246 14200 7246 14220
rect 8528 14208 9528 14228
rect 9586 14208 10586 14228
rect 10644 14208 11644 14228
rect 11702 14208 12702 14228
rect 12760 14208 13760 14228
rect 15034 14216 16034 14236
rect 16092 14216 17092 14236
rect 17150 14216 18150 14236
rect 18208 14216 19208 14236
rect 19266 14216 20266 14236
rect 21974 14226 26600 14268
rect 28496 14242 33122 14284
rect 35006 14248 39632 14290
rect 41496 14248 46122 14290
rect 48084 14270 52710 14312
rect 54598 14284 59224 14326
rect 54148 14278 59380 14284
rect 47634 14264 52866 14270
rect 34556 14242 39788 14248
rect 28046 14236 33278 14242
rect 21524 14220 26756 14226
rect 21524 14200 22524 14220
rect 22582 14200 23582 14220
rect 23640 14200 24640 14220
rect 24698 14200 25698 14220
rect 25756 14200 26756 14220
rect 28046 14216 29046 14236
rect 29104 14216 30104 14236
rect 30162 14216 31162 14236
rect 31220 14216 32220 14236
rect 32278 14216 33278 14236
rect 34556 14222 35556 14242
rect 35614 14222 36614 14242
rect 36672 14222 37672 14242
rect 37730 14222 38730 14242
rect 38788 14222 39788 14242
rect 41046 14242 46278 14248
rect 47634 14244 48634 14264
rect 48692 14244 49692 14264
rect 49750 14244 50750 14264
rect 50808 14244 51808 14264
rect 51866 14244 52866 14264
rect 54148 14258 55148 14278
rect 55206 14258 56206 14278
rect 56264 14258 57264 14278
rect 57322 14258 58322 14278
rect 58380 14258 59380 14278
rect 41046 14222 42046 14242
rect 42104 14222 43104 14242
rect 43162 14222 44162 14242
rect 44220 14222 45220 14242
rect 45278 14222 46278 14242
rect 2014 13174 3014 13200
rect 3072 13174 4072 13200
rect 4130 13174 5130 13200
rect 5188 13174 6188 13200
rect 6246 13174 7246 13200
rect 8528 13182 9528 13208
rect 9586 13182 10586 13208
rect 10644 13182 11644 13208
rect 11702 13182 12702 13208
rect 12760 13182 13760 13208
rect 15034 13190 16034 13216
rect 16092 13190 17092 13216
rect 17150 13190 18150 13216
rect 18208 13190 19208 13216
rect 19266 13190 20266 13216
rect 2266 13132 2800 13174
rect 3304 13132 3838 13174
rect 4422 13132 4956 13174
rect 5438 13132 5972 13174
rect 6504 13132 7038 13174
rect 8780 13140 9314 13182
rect 9818 13140 10352 13182
rect 10936 13140 11470 13182
rect 11952 13140 12486 13182
rect 13018 13140 13552 13182
rect 15286 13148 15820 13190
rect 16324 13148 16858 13190
rect 17442 13148 17976 13190
rect 18458 13148 18992 13190
rect 19524 13148 20058 13190
rect 21524 13174 22524 13200
rect 22582 13174 23582 13200
rect 23640 13174 24640 13200
rect 24698 13174 25698 13200
rect 25756 13174 26756 13200
rect 28046 13190 29046 13216
rect 29104 13190 30104 13216
rect 30162 13190 31162 13216
rect 31220 13190 32220 13216
rect 32278 13190 33278 13216
rect 34556 13196 35556 13222
rect 35614 13196 36614 13222
rect 36672 13196 37672 13222
rect 37730 13196 38730 13222
rect 38788 13196 39788 13222
rect 41046 13196 42046 13222
rect 42104 13196 43104 13222
rect 43162 13196 44162 13222
rect 44220 13196 45220 13222
rect 45278 13196 46278 13222
rect 47634 13218 48634 13244
rect 48692 13218 49692 13244
rect 49750 13218 50750 13244
rect 50808 13218 51808 13244
rect 51866 13218 52866 13244
rect 54148 13232 55148 13258
rect 55206 13232 56206 13258
rect 56264 13232 57264 13258
rect 57322 13232 58322 13258
rect 58380 13232 59380 13258
rect 2014 13106 3014 13132
rect 3072 13106 4072 13132
rect 4130 13106 5130 13132
rect 5188 13106 6188 13132
rect 6246 13106 7246 13132
rect 8528 13114 9528 13140
rect 9586 13114 10586 13140
rect 10644 13114 11644 13140
rect 11702 13114 12702 13140
rect 12760 13114 13760 13140
rect 15034 13122 16034 13148
rect 16092 13122 17092 13148
rect 17150 13122 18150 13148
rect 18208 13122 19208 13148
rect 19266 13122 20266 13148
rect 21776 13132 22310 13174
rect 22814 13132 23348 13174
rect 23932 13132 24466 13174
rect 24948 13132 25482 13174
rect 26014 13132 26548 13174
rect 28298 13148 28832 13190
rect 29336 13148 29870 13190
rect 30454 13148 30988 13190
rect 31470 13148 32004 13190
rect 32536 13148 33070 13190
rect 34808 13154 35342 13196
rect 35846 13154 36380 13196
rect 36964 13154 37498 13196
rect 37980 13154 38514 13196
rect 39046 13154 39580 13196
rect 41298 13154 41832 13196
rect 42336 13154 42870 13196
rect 43454 13154 43988 13196
rect 44470 13154 45004 13196
rect 45536 13154 46070 13196
rect 47886 13176 48420 13218
rect 48924 13176 49458 13218
rect 50042 13176 50576 13218
rect 51058 13176 51592 13218
rect 52124 13176 52658 13218
rect 54400 13190 54934 13232
rect 55438 13190 55972 13232
rect 56556 13190 57090 13232
rect 57572 13190 58106 13232
rect 58638 13190 59172 13232
rect 2014 12080 3014 12106
rect 3072 12080 4072 12106
rect 4130 12080 5130 12106
rect 5188 12080 6188 12106
rect 6246 12080 7246 12106
rect 2302 12038 2836 12080
rect 3258 12038 3792 12080
rect 4366 12038 4900 12080
rect 5472 12038 6006 12080
rect 6502 12038 7036 12080
rect 2014 12012 3014 12038
rect 3072 12012 4072 12038
rect 4130 12012 5130 12038
rect 5188 12012 6188 12038
rect 6246 12012 7246 12038
rect 8528 12088 9528 12114
rect 9586 12088 10586 12114
rect 10644 12088 11644 12114
rect 11702 12088 12702 12114
rect 12760 12088 13760 12114
rect 8816 12046 9350 12088
rect 9772 12046 10306 12088
rect 10880 12046 11414 12088
rect 11986 12046 12520 12088
rect 13016 12046 13550 12088
rect 8528 12020 9528 12046
rect 9586 12020 10586 12046
rect 10644 12020 11644 12046
rect 11702 12020 12702 12046
rect 12760 12020 13760 12046
rect 2014 10986 3014 11012
rect 3072 10986 4072 11012
rect 4130 10986 5130 11012
rect 5188 10986 6188 11012
rect 6246 10986 7246 11012
rect 2238 10944 2772 10986
rect 3292 10944 3826 10986
rect 4344 10944 4878 10986
rect 5452 10944 5986 10986
rect 6508 10944 7042 10986
rect 2014 10918 3014 10944
rect 3072 10918 4072 10944
rect 4130 10918 5130 10944
rect 5188 10918 6188 10944
rect 6246 10918 7246 10944
rect 21524 13106 22524 13132
rect 22582 13106 23582 13132
rect 23640 13106 24640 13132
rect 24698 13106 25698 13132
rect 25756 13106 26756 13132
rect 28046 13122 29046 13148
rect 29104 13122 30104 13148
rect 30162 13122 31162 13148
rect 31220 13122 32220 13148
rect 32278 13122 33278 13148
rect 34556 13128 35556 13154
rect 35614 13128 36614 13154
rect 36672 13128 37672 13154
rect 37730 13128 38730 13154
rect 38788 13128 39788 13154
rect 41046 13128 42046 13154
rect 42104 13128 43104 13154
rect 43162 13128 44162 13154
rect 44220 13128 45220 13154
rect 45278 13128 46278 13154
rect 47634 13150 48634 13176
rect 48692 13150 49692 13176
rect 49750 13150 50750 13176
rect 50808 13150 51808 13176
rect 51866 13150 52866 13176
rect 54148 13164 55148 13190
rect 55206 13164 56206 13190
rect 56264 13164 57264 13190
rect 57322 13164 58322 13190
rect 58380 13164 59380 13190
rect 15034 12096 16034 12122
rect 16092 12096 17092 12122
rect 17150 12096 18150 12122
rect 18208 12096 19208 12122
rect 19266 12096 20266 12122
rect 15322 12054 15856 12096
rect 16278 12054 16812 12096
rect 17386 12054 17920 12096
rect 18492 12054 19026 12096
rect 19522 12054 20056 12096
rect 15034 12028 16034 12054
rect 16092 12028 17092 12054
rect 17150 12028 18150 12054
rect 18208 12028 19208 12054
rect 19266 12028 20266 12054
rect 8528 10994 9528 11020
rect 9586 10994 10586 11020
rect 10644 10994 11644 11020
rect 11702 10994 12702 11020
rect 12760 10994 13760 11020
rect 8752 10952 9286 10994
rect 9806 10952 10340 10994
rect 10858 10952 11392 10994
rect 11966 10952 12500 10994
rect 13022 10952 13556 10994
rect 8528 10926 9528 10952
rect 9586 10926 10586 10952
rect 10644 10926 11644 10952
rect 11702 10926 12702 10952
rect 12760 10926 13760 10952
rect 21524 12080 22524 12106
rect 22582 12080 23582 12106
rect 23640 12080 24640 12106
rect 24698 12080 25698 12106
rect 25756 12080 26756 12106
rect 21812 12038 22346 12080
rect 22768 12038 23302 12080
rect 23876 12038 24410 12080
rect 24982 12038 25516 12080
rect 26012 12038 26546 12080
rect 21524 12012 22524 12038
rect 22582 12012 23582 12038
rect 23640 12012 24640 12038
rect 24698 12012 25698 12038
rect 25756 12012 26756 12038
rect 15034 11002 16034 11028
rect 16092 11002 17092 11028
rect 17150 11002 18150 11028
rect 18208 11002 19208 11028
rect 19266 11002 20266 11028
rect 15258 10960 15792 11002
rect 16312 10960 16846 11002
rect 17364 10960 17898 11002
rect 18472 10960 19006 11002
rect 19528 10960 20062 11002
rect 15034 10934 16034 10960
rect 16092 10934 17092 10960
rect 17150 10934 18150 10960
rect 18208 10934 19208 10960
rect 19266 10934 20266 10960
rect 28046 12096 29046 12122
rect 29104 12096 30104 12122
rect 30162 12096 31162 12122
rect 31220 12096 32220 12122
rect 32278 12096 33278 12122
rect 28334 12054 28868 12096
rect 29290 12054 29824 12096
rect 30398 12054 30932 12096
rect 31504 12054 32038 12096
rect 32534 12054 33068 12096
rect 28046 12028 29046 12054
rect 29104 12028 30104 12054
rect 30162 12028 31162 12054
rect 31220 12028 32220 12054
rect 32278 12028 33278 12054
rect 21524 10986 22524 11012
rect 22582 10986 23582 11012
rect 23640 10986 24640 11012
rect 24698 10986 25698 11012
rect 25756 10986 26756 11012
rect 21748 10944 22282 10986
rect 22802 10944 23336 10986
rect 23854 10944 24388 10986
rect 24962 10944 25496 10986
rect 26018 10944 26552 10986
rect 21524 10918 22524 10944
rect 22582 10918 23582 10944
rect 23640 10918 24640 10944
rect 24698 10918 25698 10944
rect 25756 10918 26756 10944
rect 2014 9892 3014 9918
rect 3072 9892 4072 9918
rect 4130 9892 5130 9918
rect 5188 9892 6188 9918
rect 6246 9892 7246 9918
rect 8528 9900 9528 9926
rect 9586 9900 10586 9926
rect 10644 9900 11644 9926
rect 11702 9900 12702 9926
rect 12760 9900 13760 9926
rect 15034 9908 16034 9934
rect 16092 9908 17092 9934
rect 17150 9908 18150 9934
rect 18208 9908 19208 9934
rect 19266 9908 20266 9934
rect 34556 12102 35556 12128
rect 35614 12102 36614 12128
rect 36672 12102 37672 12128
rect 37730 12102 38730 12128
rect 38788 12102 39788 12128
rect 34844 12060 35378 12102
rect 35800 12060 36334 12102
rect 36908 12060 37442 12102
rect 38014 12060 38548 12102
rect 39044 12060 39578 12102
rect 34556 12034 35556 12060
rect 35614 12034 36614 12060
rect 36672 12034 37672 12060
rect 37730 12034 38730 12060
rect 38788 12034 39788 12060
rect 28046 11002 29046 11028
rect 29104 11002 30104 11028
rect 30162 11002 31162 11028
rect 31220 11002 32220 11028
rect 32278 11002 33278 11028
rect 28270 10960 28804 11002
rect 29324 10960 29858 11002
rect 30376 10960 30910 11002
rect 31484 10960 32018 11002
rect 32540 10960 33074 11002
rect 28046 10934 29046 10960
rect 29104 10934 30104 10960
rect 30162 10934 31162 10960
rect 31220 10934 32220 10960
rect 32278 10934 33278 10960
rect 41046 12102 42046 12128
rect 42104 12102 43104 12128
rect 43162 12102 44162 12128
rect 44220 12102 45220 12128
rect 45278 12102 46278 12128
rect 41334 12060 41868 12102
rect 42290 12060 42824 12102
rect 43398 12060 43932 12102
rect 44504 12060 45038 12102
rect 45534 12060 46068 12102
rect 41046 12034 42046 12060
rect 42104 12034 43104 12060
rect 43162 12034 44162 12060
rect 44220 12034 45220 12060
rect 45278 12034 46278 12060
rect 34556 11008 35556 11034
rect 35614 11008 36614 11034
rect 36672 11008 37672 11034
rect 37730 11008 38730 11034
rect 38788 11008 39788 11034
rect 34780 10966 35314 11008
rect 35834 10966 36368 11008
rect 36886 10966 37420 11008
rect 37994 10966 38528 11008
rect 39050 10966 39584 11008
rect 34556 10940 35556 10966
rect 35614 10940 36614 10966
rect 36672 10940 37672 10966
rect 37730 10940 38730 10966
rect 38788 10940 39788 10966
rect 47634 12124 48634 12150
rect 48692 12124 49692 12150
rect 49750 12124 50750 12150
rect 50808 12124 51808 12150
rect 51866 12124 52866 12150
rect 47922 12082 48456 12124
rect 48878 12082 49412 12124
rect 49986 12082 50520 12124
rect 51092 12082 51626 12124
rect 52122 12082 52656 12124
rect 47634 12056 48634 12082
rect 48692 12056 49692 12082
rect 49750 12056 50750 12082
rect 50808 12056 51808 12082
rect 51866 12056 52866 12082
rect 41046 11008 42046 11034
rect 42104 11008 43104 11034
rect 43162 11008 44162 11034
rect 44220 11008 45220 11034
rect 45278 11008 46278 11034
rect 41270 10966 41804 11008
rect 42324 10966 42858 11008
rect 43376 10966 43910 11008
rect 44484 10966 45018 11008
rect 45540 10966 46074 11008
rect 41046 10940 42046 10966
rect 42104 10940 43104 10966
rect 43162 10940 44162 10966
rect 44220 10940 45220 10966
rect 45278 10940 46278 10966
rect 54148 12138 55148 12164
rect 55206 12138 56206 12164
rect 56264 12138 57264 12164
rect 57322 12138 58322 12164
rect 58380 12138 59380 12164
rect 54436 12096 54970 12138
rect 55392 12096 55926 12138
rect 56500 12096 57034 12138
rect 57606 12096 58140 12138
rect 58636 12096 59170 12138
rect 54148 12070 55148 12096
rect 55206 12070 56206 12096
rect 56264 12070 57264 12096
rect 57322 12070 58322 12096
rect 58380 12070 59380 12096
rect 47634 11030 48634 11056
rect 48692 11030 49692 11056
rect 49750 11030 50750 11056
rect 50808 11030 51808 11056
rect 51866 11030 52866 11056
rect 47858 10988 48392 11030
rect 48912 10988 49446 11030
rect 49964 10988 50498 11030
rect 51072 10988 51606 11030
rect 52128 10988 52662 11030
rect 47634 10962 48634 10988
rect 48692 10962 49692 10988
rect 49750 10962 50750 10988
rect 50808 10962 51808 10988
rect 51866 10962 52866 10988
rect 54148 11044 55148 11070
rect 55206 11044 56206 11070
rect 56264 11044 57264 11070
rect 57322 11044 58322 11070
rect 58380 11044 59380 11070
rect 54372 11002 54906 11044
rect 55426 11002 55960 11044
rect 56478 11002 57012 11044
rect 57586 11002 58120 11044
rect 58642 11002 59176 11044
rect 54148 10976 55148 11002
rect 55206 10976 56206 11002
rect 56264 10976 57264 11002
rect 57322 10976 58322 11002
rect 58380 10976 59380 11002
rect 2266 9850 2800 9892
rect 3364 9850 3898 9892
rect 4392 9850 4926 9892
rect 5356 9850 5890 9892
rect 6456 9850 6990 9892
rect 8780 9858 9314 9900
rect 9878 9858 10412 9900
rect 10906 9858 11440 9900
rect 11870 9858 12404 9900
rect 12970 9858 13504 9900
rect 15286 9866 15820 9908
rect 16384 9866 16918 9908
rect 17412 9866 17946 9908
rect 18376 9866 18910 9908
rect 19476 9866 20010 9908
rect 21524 9892 22524 9918
rect 22582 9892 23582 9918
rect 23640 9892 24640 9918
rect 24698 9892 25698 9918
rect 25756 9892 26756 9918
rect 28046 9908 29046 9934
rect 29104 9908 30104 9934
rect 30162 9908 31162 9934
rect 31220 9908 32220 9934
rect 32278 9908 33278 9934
rect 34556 9914 35556 9940
rect 35614 9914 36614 9940
rect 36672 9914 37672 9940
rect 37730 9914 38730 9940
rect 38788 9914 39788 9940
rect 41046 9914 42046 9940
rect 42104 9914 43104 9940
rect 43162 9914 44162 9940
rect 44220 9914 45220 9940
rect 45278 9914 46278 9940
rect 47634 9936 48634 9962
rect 48692 9936 49692 9962
rect 49750 9936 50750 9962
rect 50808 9936 51808 9962
rect 51866 9936 52866 9962
rect 54148 9950 55148 9976
rect 55206 9950 56206 9976
rect 56264 9950 57264 9976
rect 57322 9950 58322 9976
rect 58380 9950 59380 9976
rect 2014 9824 3014 9850
rect 3072 9824 4072 9850
rect 4130 9824 5130 9850
rect 5188 9824 6188 9850
rect 6246 9824 7246 9850
rect 8528 9832 9528 9858
rect 9586 9832 10586 9858
rect 10644 9832 11644 9858
rect 11702 9832 12702 9858
rect 12760 9832 13760 9858
rect 15034 9840 16034 9866
rect 16092 9840 17092 9866
rect 17150 9840 18150 9866
rect 18208 9840 19208 9866
rect 19266 9840 20266 9866
rect 21776 9850 22310 9892
rect 22874 9850 23408 9892
rect 23902 9850 24436 9892
rect 24866 9850 25400 9892
rect 25966 9850 26500 9892
rect 28298 9866 28832 9908
rect 29396 9866 29930 9908
rect 30424 9866 30958 9908
rect 31388 9866 31922 9908
rect 32488 9866 33022 9908
rect 34808 9872 35342 9914
rect 35906 9872 36440 9914
rect 36934 9872 37468 9914
rect 37898 9872 38432 9914
rect 38998 9872 39532 9914
rect 41298 9872 41832 9914
rect 42396 9872 42930 9914
rect 43424 9872 43958 9914
rect 44388 9872 44922 9914
rect 45488 9872 46022 9914
rect 47886 9894 48420 9936
rect 48984 9894 49518 9936
rect 50012 9894 50546 9936
rect 50976 9894 51510 9936
rect 52076 9894 52610 9936
rect 54400 9908 54934 9950
rect 55498 9908 56032 9950
rect 56526 9908 57060 9950
rect 57490 9908 58024 9950
rect 58590 9908 59124 9950
rect 21524 9824 22524 9850
rect 22582 9824 23582 9850
rect 23640 9824 24640 9850
rect 24698 9824 25698 9850
rect 25756 9824 26756 9850
rect 28046 9840 29046 9866
rect 29104 9840 30104 9866
rect 30162 9840 31162 9866
rect 31220 9840 32220 9866
rect 32278 9840 33278 9866
rect 34556 9846 35556 9872
rect 35614 9846 36614 9872
rect 36672 9846 37672 9872
rect 37730 9846 38730 9872
rect 38788 9846 39788 9872
rect 41046 9846 42046 9872
rect 42104 9846 43104 9872
rect 43162 9846 44162 9872
rect 44220 9846 45220 9872
rect 45278 9846 46278 9872
rect 47634 9868 48634 9894
rect 48692 9868 49692 9894
rect 49750 9868 50750 9894
rect 50808 9868 51808 9894
rect 51866 9868 52866 9894
rect 54148 9882 55148 9908
rect 55206 9882 56206 9908
rect 56264 9882 57264 9908
rect 57322 9882 58322 9908
rect 58380 9882 59380 9908
rect 2014 8798 3014 8824
rect 3072 8798 4072 8824
rect 4130 8798 5130 8824
rect 5188 8798 6188 8824
rect 6246 8798 7246 8824
rect 8528 8814 9528 8832
rect 9586 8814 10586 8832
rect 10644 8814 11644 8832
rect 11702 8814 12702 8832
rect 12760 8814 13760 8832
rect 15034 8822 16034 8840
rect 16092 8822 17092 8840
rect 17150 8822 18150 8840
rect 18208 8822 19208 8840
rect 19266 8822 20266 8840
rect 47634 8852 48634 8868
rect 48692 8852 49692 8868
rect 49750 8852 50750 8868
rect 50808 8852 51808 8868
rect 51866 8852 52866 8868
rect 54148 8864 55148 8882
rect 55206 8864 56206 8882
rect 56264 8864 57264 8882
rect 57322 8864 58322 8882
rect 58380 8864 59380 8882
rect 54148 8856 59380 8864
rect 15034 8814 20266 8822
rect 8528 8806 13760 8814
rect 2612 8360 2878 8798
rect 3352 8360 3618 8798
rect 4480 8360 4746 8798
rect 5398 8360 5664 8798
rect 6564 8360 6830 8798
rect 8902 8728 13454 8806
rect 11142 8368 11322 8728
rect 15492 8700 20048 8814
rect 21524 8804 22524 8824
rect 22582 8804 23582 8824
rect 23640 8804 24640 8824
rect 24698 8804 25698 8824
rect 25756 8804 26756 8824
rect 28046 8820 29046 8840
rect 29104 8820 30104 8840
rect 30162 8820 31162 8840
rect 31220 8820 32220 8840
rect 32278 8820 33278 8840
rect 34556 8828 35556 8846
rect 35614 8828 36614 8846
rect 36672 8828 37672 8846
rect 37730 8828 38730 8846
rect 38788 8828 39788 8846
rect 34556 8820 39788 8828
rect 41046 8826 42046 8846
rect 42104 8826 43104 8846
rect 43162 8826 44162 8846
rect 44220 8826 45220 8846
rect 45278 8826 46278 8846
rect 47634 8842 52866 8852
rect 41046 8820 46278 8826
rect 28046 8814 33278 8820
rect 21524 8798 26756 8804
rect 17604 8376 17814 8700
rect 22064 8536 26522 8798
rect 28490 8634 32784 8814
rect 2482 8318 7108 8360
rect 8996 8326 13622 8368
rect 15502 8334 20128 8376
rect 23138 8360 23344 8536
rect 30554 8376 30760 8634
rect 35074 8600 39566 8820
rect 41522 8602 46018 8820
rect 48096 8648 52572 8842
rect 54648 8668 59120 8856
rect 36926 8382 37132 8600
rect 42486 8382 42712 8602
rect 49102 8404 49328 8648
rect 55526 8418 55752 8668
rect 15052 8328 20284 8334
rect 8546 8320 13778 8326
rect 2032 8312 7264 8318
rect 2032 8292 3032 8312
rect 3090 8292 4090 8312
rect 4148 8292 5148 8312
rect 5206 8292 6206 8312
rect 6264 8292 7264 8312
rect 8546 8300 9546 8320
rect 9604 8300 10604 8320
rect 10662 8300 11662 8320
rect 11720 8300 12720 8320
rect 12778 8300 13778 8320
rect 15052 8308 16052 8328
rect 16110 8308 17110 8328
rect 17168 8308 18168 8328
rect 18226 8308 19226 8328
rect 19284 8308 20284 8328
rect 21992 8318 26618 8360
rect 28514 8334 33140 8376
rect 35024 8340 39650 8382
rect 41514 8340 46140 8382
rect 48102 8362 52728 8404
rect 54616 8376 59242 8418
rect 54166 8370 59398 8376
rect 47652 8356 52884 8362
rect 34574 8334 39806 8340
rect 28064 8328 33296 8334
rect 21542 8312 26774 8318
rect 21542 8292 22542 8312
rect 22600 8292 23600 8312
rect 23658 8292 24658 8312
rect 24716 8292 25716 8312
rect 25774 8292 26774 8312
rect 28064 8308 29064 8328
rect 29122 8308 30122 8328
rect 30180 8308 31180 8328
rect 31238 8308 32238 8328
rect 32296 8308 33296 8328
rect 34574 8314 35574 8334
rect 35632 8314 36632 8334
rect 36690 8314 37690 8334
rect 37748 8314 38748 8334
rect 38806 8314 39806 8334
rect 41064 8334 46296 8340
rect 47652 8336 48652 8356
rect 48710 8336 49710 8356
rect 49768 8336 50768 8356
rect 50826 8336 51826 8356
rect 51884 8336 52884 8356
rect 54166 8350 55166 8370
rect 55224 8350 56224 8370
rect 56282 8350 57282 8370
rect 57340 8350 58340 8370
rect 58398 8350 59398 8370
rect 41064 8314 42064 8334
rect 42122 8314 43122 8334
rect 43180 8314 44180 8334
rect 44238 8314 45238 8334
rect 45296 8314 46296 8334
rect 2032 7266 3032 7292
rect 3090 7266 4090 7292
rect 4148 7266 5148 7292
rect 5206 7266 6206 7292
rect 6264 7266 7264 7292
rect 8546 7274 9546 7300
rect 9604 7274 10604 7300
rect 10662 7274 11662 7300
rect 11720 7274 12720 7300
rect 12778 7274 13778 7300
rect 15052 7282 16052 7308
rect 16110 7282 17110 7308
rect 17168 7282 18168 7308
rect 18226 7282 19226 7308
rect 19284 7282 20284 7308
rect 2284 7224 2818 7266
rect 3322 7224 3856 7266
rect 4440 7224 4974 7266
rect 5456 7224 5990 7266
rect 6522 7224 7056 7266
rect 8798 7232 9332 7274
rect 9836 7232 10370 7274
rect 10954 7232 11488 7274
rect 11970 7232 12504 7274
rect 13036 7232 13570 7274
rect 15304 7240 15838 7282
rect 16342 7240 16876 7282
rect 17460 7240 17994 7282
rect 18476 7240 19010 7282
rect 19542 7240 20076 7282
rect 21542 7266 22542 7292
rect 22600 7266 23600 7292
rect 23658 7266 24658 7292
rect 24716 7266 25716 7292
rect 25774 7266 26774 7292
rect 28064 7282 29064 7308
rect 29122 7282 30122 7308
rect 30180 7282 31180 7308
rect 31238 7282 32238 7308
rect 32296 7282 33296 7308
rect 34574 7288 35574 7314
rect 35632 7288 36632 7314
rect 36690 7288 37690 7314
rect 37748 7288 38748 7314
rect 38806 7288 39806 7314
rect 41064 7288 42064 7314
rect 42122 7288 43122 7314
rect 43180 7288 44180 7314
rect 44238 7288 45238 7314
rect 45296 7288 46296 7314
rect 47652 7310 48652 7336
rect 48710 7310 49710 7336
rect 49768 7310 50768 7336
rect 50826 7310 51826 7336
rect 51884 7310 52884 7336
rect 54166 7324 55166 7350
rect 55224 7324 56224 7350
rect 56282 7324 57282 7350
rect 57340 7324 58340 7350
rect 58398 7324 59398 7350
rect 2032 7198 3032 7224
rect 3090 7198 4090 7224
rect 4148 7198 5148 7224
rect 5206 7198 6206 7224
rect 6264 7198 7264 7224
rect 8546 7206 9546 7232
rect 9604 7206 10604 7232
rect 10662 7206 11662 7232
rect 11720 7206 12720 7232
rect 12778 7206 13778 7232
rect 15052 7214 16052 7240
rect 16110 7214 17110 7240
rect 17168 7214 18168 7240
rect 18226 7214 19226 7240
rect 19284 7214 20284 7240
rect 21794 7224 22328 7266
rect 22832 7224 23366 7266
rect 23950 7224 24484 7266
rect 24966 7224 25500 7266
rect 26032 7224 26566 7266
rect 28316 7240 28850 7282
rect 29354 7240 29888 7282
rect 30472 7240 31006 7282
rect 31488 7240 32022 7282
rect 32554 7240 33088 7282
rect 34826 7246 35360 7288
rect 35864 7246 36398 7288
rect 36982 7246 37516 7288
rect 37998 7246 38532 7288
rect 39064 7246 39598 7288
rect 41316 7246 41850 7288
rect 42354 7246 42888 7288
rect 43472 7246 44006 7288
rect 44488 7246 45022 7288
rect 45554 7246 46088 7288
rect 47904 7268 48438 7310
rect 48942 7268 49476 7310
rect 50060 7268 50594 7310
rect 51076 7268 51610 7310
rect 52142 7268 52676 7310
rect 54418 7282 54952 7324
rect 55456 7282 55990 7324
rect 56574 7282 57108 7324
rect 57590 7282 58124 7324
rect 58656 7282 59190 7324
rect 2032 6172 3032 6198
rect 3090 6172 4090 6198
rect 4148 6172 5148 6198
rect 5206 6172 6206 6198
rect 6264 6172 7264 6198
rect 2320 6130 2854 6172
rect 3276 6130 3810 6172
rect 4384 6130 4918 6172
rect 5490 6130 6024 6172
rect 6520 6130 7054 6172
rect 2032 6104 3032 6130
rect 3090 6104 4090 6130
rect 4148 6104 5148 6130
rect 5206 6104 6206 6130
rect 6264 6104 7264 6130
rect 8546 6180 9546 6206
rect 9604 6180 10604 6206
rect 10662 6180 11662 6206
rect 11720 6180 12720 6206
rect 12778 6180 13778 6206
rect 8834 6138 9368 6180
rect 9790 6138 10324 6180
rect 10898 6138 11432 6180
rect 12004 6138 12538 6180
rect 13034 6138 13568 6180
rect 8546 6112 9546 6138
rect 9604 6112 10604 6138
rect 10662 6112 11662 6138
rect 11720 6112 12720 6138
rect 12778 6112 13778 6138
rect 2032 5078 3032 5104
rect 3090 5078 4090 5104
rect 4148 5078 5148 5104
rect 5206 5078 6206 5104
rect 6264 5078 7264 5104
rect 2256 5036 2790 5078
rect 3310 5036 3844 5078
rect 4362 5036 4896 5078
rect 5470 5036 6004 5078
rect 6526 5036 7060 5078
rect 2032 5010 3032 5036
rect 3090 5010 4090 5036
rect 4148 5010 5148 5036
rect 5206 5010 6206 5036
rect 6264 5010 7264 5036
rect 21542 7198 22542 7224
rect 22600 7198 23600 7224
rect 23658 7198 24658 7224
rect 24716 7198 25716 7224
rect 25774 7198 26774 7224
rect 28064 7214 29064 7240
rect 29122 7214 30122 7240
rect 30180 7214 31180 7240
rect 31238 7214 32238 7240
rect 32296 7214 33296 7240
rect 34574 7220 35574 7246
rect 35632 7220 36632 7246
rect 36690 7220 37690 7246
rect 37748 7220 38748 7246
rect 38806 7220 39806 7246
rect 41064 7220 42064 7246
rect 42122 7220 43122 7246
rect 43180 7220 44180 7246
rect 44238 7220 45238 7246
rect 45296 7220 46296 7246
rect 47652 7242 48652 7268
rect 48710 7242 49710 7268
rect 49768 7242 50768 7268
rect 50826 7242 51826 7268
rect 51884 7242 52884 7268
rect 54166 7256 55166 7282
rect 55224 7256 56224 7282
rect 56282 7256 57282 7282
rect 57340 7256 58340 7282
rect 58398 7256 59398 7282
rect 15052 6188 16052 6214
rect 16110 6188 17110 6214
rect 17168 6188 18168 6214
rect 18226 6188 19226 6214
rect 19284 6188 20284 6214
rect 15340 6146 15874 6188
rect 16296 6146 16830 6188
rect 17404 6146 17938 6188
rect 18510 6146 19044 6188
rect 19540 6146 20074 6188
rect 15052 6120 16052 6146
rect 16110 6120 17110 6146
rect 17168 6120 18168 6146
rect 18226 6120 19226 6146
rect 19284 6120 20284 6146
rect 8546 5086 9546 5112
rect 9604 5086 10604 5112
rect 10662 5086 11662 5112
rect 11720 5086 12720 5112
rect 12778 5086 13778 5112
rect 8770 5044 9304 5086
rect 9824 5044 10358 5086
rect 10876 5044 11410 5086
rect 11984 5044 12518 5086
rect 13040 5044 13574 5086
rect 8546 5018 9546 5044
rect 9604 5018 10604 5044
rect 10662 5018 11662 5044
rect 11720 5018 12720 5044
rect 12778 5018 13778 5044
rect 21542 6172 22542 6198
rect 22600 6172 23600 6198
rect 23658 6172 24658 6198
rect 24716 6172 25716 6198
rect 25774 6172 26774 6198
rect 21830 6130 22364 6172
rect 22786 6130 23320 6172
rect 23894 6130 24428 6172
rect 25000 6130 25534 6172
rect 26030 6130 26564 6172
rect 21542 6104 22542 6130
rect 22600 6104 23600 6130
rect 23658 6104 24658 6130
rect 24716 6104 25716 6130
rect 25774 6104 26774 6130
rect 15052 5094 16052 5120
rect 16110 5094 17110 5120
rect 17168 5094 18168 5120
rect 18226 5094 19226 5120
rect 19284 5094 20284 5120
rect 15276 5052 15810 5094
rect 16330 5052 16864 5094
rect 17382 5052 17916 5094
rect 18490 5052 19024 5094
rect 19546 5052 20080 5094
rect 15052 5026 16052 5052
rect 16110 5026 17110 5052
rect 17168 5026 18168 5052
rect 18226 5026 19226 5052
rect 19284 5026 20284 5052
rect 28064 6188 29064 6214
rect 29122 6188 30122 6214
rect 30180 6188 31180 6214
rect 31238 6188 32238 6214
rect 32296 6188 33296 6214
rect 28352 6146 28886 6188
rect 29308 6146 29842 6188
rect 30416 6146 30950 6188
rect 31522 6146 32056 6188
rect 32552 6146 33086 6188
rect 28064 6120 29064 6146
rect 29122 6120 30122 6146
rect 30180 6120 31180 6146
rect 31238 6120 32238 6146
rect 32296 6120 33296 6146
rect 21542 5078 22542 5104
rect 22600 5078 23600 5104
rect 23658 5078 24658 5104
rect 24716 5078 25716 5104
rect 25774 5078 26774 5104
rect 21766 5036 22300 5078
rect 22820 5036 23354 5078
rect 23872 5036 24406 5078
rect 24980 5036 25514 5078
rect 26036 5036 26570 5078
rect 21542 5010 22542 5036
rect 22600 5010 23600 5036
rect 23658 5010 24658 5036
rect 24716 5010 25716 5036
rect 25774 5010 26774 5036
rect 2032 3984 3032 4010
rect 3090 3984 4090 4010
rect 4148 3984 5148 4010
rect 5206 3984 6206 4010
rect 6264 3984 7264 4010
rect 8546 3992 9546 4018
rect 9604 3992 10604 4018
rect 10662 3992 11662 4018
rect 11720 3992 12720 4018
rect 12778 3992 13778 4018
rect 15052 4000 16052 4026
rect 16110 4000 17110 4026
rect 17168 4000 18168 4026
rect 18226 4000 19226 4026
rect 19284 4000 20284 4026
rect 34574 6194 35574 6220
rect 35632 6194 36632 6220
rect 36690 6194 37690 6220
rect 37748 6194 38748 6220
rect 38806 6194 39806 6220
rect 34862 6152 35396 6194
rect 35818 6152 36352 6194
rect 36926 6152 37460 6194
rect 38032 6152 38566 6194
rect 39062 6152 39596 6194
rect 34574 6126 35574 6152
rect 35632 6126 36632 6152
rect 36690 6126 37690 6152
rect 37748 6126 38748 6152
rect 38806 6126 39806 6152
rect 28064 5094 29064 5120
rect 29122 5094 30122 5120
rect 30180 5094 31180 5120
rect 31238 5094 32238 5120
rect 32296 5094 33296 5120
rect 28288 5052 28822 5094
rect 29342 5052 29876 5094
rect 30394 5052 30928 5094
rect 31502 5052 32036 5094
rect 32558 5052 33092 5094
rect 28064 5026 29064 5052
rect 29122 5026 30122 5052
rect 30180 5026 31180 5052
rect 31238 5026 32238 5052
rect 32296 5026 33296 5052
rect 41064 6194 42064 6220
rect 42122 6194 43122 6220
rect 43180 6194 44180 6220
rect 44238 6194 45238 6220
rect 45296 6194 46296 6220
rect 41352 6152 41886 6194
rect 42308 6152 42842 6194
rect 43416 6152 43950 6194
rect 44522 6152 45056 6194
rect 45552 6152 46086 6194
rect 41064 6126 42064 6152
rect 42122 6126 43122 6152
rect 43180 6126 44180 6152
rect 44238 6126 45238 6152
rect 45296 6126 46296 6152
rect 34574 5100 35574 5126
rect 35632 5100 36632 5126
rect 36690 5100 37690 5126
rect 37748 5100 38748 5126
rect 38806 5100 39806 5126
rect 34798 5058 35332 5100
rect 35852 5058 36386 5100
rect 36904 5058 37438 5100
rect 38012 5058 38546 5100
rect 39068 5058 39602 5100
rect 34574 5032 35574 5058
rect 35632 5032 36632 5058
rect 36690 5032 37690 5058
rect 37748 5032 38748 5058
rect 38806 5032 39806 5058
rect 47652 6216 48652 6242
rect 48710 6216 49710 6242
rect 49768 6216 50768 6242
rect 50826 6216 51826 6242
rect 51884 6216 52884 6242
rect 47940 6174 48474 6216
rect 48896 6174 49430 6216
rect 50004 6174 50538 6216
rect 51110 6174 51644 6216
rect 52140 6174 52674 6216
rect 47652 6148 48652 6174
rect 48710 6148 49710 6174
rect 49768 6148 50768 6174
rect 50826 6148 51826 6174
rect 51884 6148 52884 6174
rect 41064 5100 42064 5126
rect 42122 5100 43122 5126
rect 43180 5100 44180 5126
rect 44238 5100 45238 5126
rect 45296 5100 46296 5126
rect 41288 5058 41822 5100
rect 42342 5058 42876 5100
rect 43394 5058 43928 5100
rect 44502 5058 45036 5100
rect 45558 5058 46092 5100
rect 41064 5032 42064 5058
rect 42122 5032 43122 5058
rect 43180 5032 44180 5058
rect 44238 5032 45238 5058
rect 45296 5032 46296 5058
rect 54166 6230 55166 6256
rect 55224 6230 56224 6256
rect 56282 6230 57282 6256
rect 57340 6230 58340 6256
rect 58398 6230 59398 6256
rect 54454 6188 54988 6230
rect 55410 6188 55944 6230
rect 56518 6188 57052 6230
rect 57624 6188 58158 6230
rect 58654 6188 59188 6230
rect 54166 6162 55166 6188
rect 55224 6162 56224 6188
rect 56282 6162 57282 6188
rect 57340 6162 58340 6188
rect 58398 6162 59398 6188
rect 47652 5122 48652 5148
rect 48710 5122 49710 5148
rect 49768 5122 50768 5148
rect 50826 5122 51826 5148
rect 51884 5122 52884 5148
rect 47876 5080 48410 5122
rect 48930 5080 49464 5122
rect 49982 5080 50516 5122
rect 51090 5080 51624 5122
rect 52146 5080 52680 5122
rect 47652 5054 48652 5080
rect 48710 5054 49710 5080
rect 49768 5054 50768 5080
rect 50826 5054 51826 5080
rect 51884 5054 52884 5080
rect 54166 5136 55166 5162
rect 55224 5136 56224 5162
rect 56282 5136 57282 5162
rect 57340 5136 58340 5162
rect 58398 5136 59398 5162
rect 54390 5094 54924 5136
rect 55444 5094 55978 5136
rect 56496 5094 57030 5136
rect 57604 5094 58138 5136
rect 58660 5094 59194 5136
rect 54166 5068 55166 5094
rect 55224 5068 56224 5094
rect 56282 5068 57282 5094
rect 57340 5068 58340 5094
rect 58398 5068 59398 5094
rect 2284 3942 2818 3984
rect 3382 3942 3916 3984
rect 4410 3942 4944 3984
rect 5374 3942 5908 3984
rect 6474 3942 7008 3984
rect 8798 3950 9332 3992
rect 9896 3950 10430 3992
rect 10924 3950 11458 3992
rect 11888 3950 12422 3992
rect 12988 3950 13522 3992
rect 15304 3958 15838 4000
rect 16402 3958 16936 4000
rect 17430 3958 17964 4000
rect 18394 3958 18928 4000
rect 19494 3958 20028 4000
rect 21542 3984 22542 4010
rect 22600 3984 23600 4010
rect 23658 3984 24658 4010
rect 24716 3984 25716 4010
rect 25774 3984 26774 4010
rect 28064 4000 29064 4026
rect 29122 4000 30122 4026
rect 30180 4000 31180 4026
rect 31238 4000 32238 4026
rect 32296 4000 33296 4026
rect 34574 4006 35574 4032
rect 35632 4006 36632 4032
rect 36690 4006 37690 4032
rect 37748 4006 38748 4032
rect 38806 4006 39806 4032
rect 41064 4006 42064 4032
rect 42122 4006 43122 4032
rect 43180 4006 44180 4032
rect 44238 4006 45238 4032
rect 45296 4006 46296 4032
rect 47652 4028 48652 4054
rect 48710 4028 49710 4054
rect 49768 4028 50768 4054
rect 50826 4028 51826 4054
rect 51884 4028 52884 4054
rect 54166 4042 55166 4068
rect 55224 4042 56224 4068
rect 56282 4042 57282 4068
rect 57340 4042 58340 4068
rect 58398 4042 59398 4068
rect 2032 3916 3032 3942
rect 3090 3916 4090 3942
rect 4148 3916 5148 3942
rect 5206 3916 6206 3942
rect 6264 3916 7264 3942
rect 8546 3924 9546 3950
rect 9604 3924 10604 3950
rect 10662 3924 11662 3950
rect 11720 3924 12720 3950
rect 12778 3924 13778 3950
rect 15052 3932 16052 3958
rect 16110 3932 17110 3958
rect 17168 3932 18168 3958
rect 18226 3932 19226 3958
rect 19284 3932 20284 3958
rect 21794 3942 22328 3984
rect 22892 3942 23426 3984
rect 23920 3942 24454 3984
rect 24884 3942 25418 3984
rect 25984 3942 26518 3984
rect 28316 3958 28850 4000
rect 29414 3958 29948 4000
rect 30442 3958 30976 4000
rect 31406 3958 31940 4000
rect 32506 3958 33040 4000
rect 34826 3964 35360 4006
rect 35924 3964 36458 4006
rect 36952 3964 37486 4006
rect 37916 3964 38450 4006
rect 39016 3964 39550 4006
rect 41316 3964 41850 4006
rect 42414 3964 42948 4006
rect 43442 3964 43976 4006
rect 44406 3964 44940 4006
rect 45506 3964 46040 4006
rect 47904 3986 48438 4028
rect 49002 3986 49536 4028
rect 50030 3986 50564 4028
rect 50994 3986 51528 4028
rect 52094 3986 52628 4028
rect 54418 4000 54952 4042
rect 55516 4000 56050 4042
rect 56544 4000 57078 4042
rect 57508 4000 58042 4042
rect 58608 4000 59142 4042
rect 21542 3916 22542 3942
rect 22600 3916 23600 3942
rect 23658 3916 24658 3942
rect 24716 3916 25716 3942
rect 25774 3916 26774 3942
rect 28064 3932 29064 3958
rect 29122 3932 30122 3958
rect 30180 3932 31180 3958
rect 31238 3932 32238 3958
rect 32296 3932 33296 3958
rect 34574 3938 35574 3964
rect 35632 3938 36632 3964
rect 36690 3938 37690 3964
rect 37748 3938 38748 3964
rect 38806 3938 39806 3964
rect 41064 3938 42064 3964
rect 42122 3938 43122 3964
rect 43180 3938 44180 3964
rect 44238 3938 45238 3964
rect 45296 3938 46296 3964
rect 47652 3960 48652 3986
rect 48710 3960 49710 3986
rect 49768 3960 50768 3986
rect 50826 3960 51826 3986
rect 51884 3960 52884 3986
rect 54166 3974 55166 4000
rect 55224 3974 56224 4000
rect 56282 3974 57282 4000
rect 57340 3974 58340 4000
rect 58398 3974 59398 4000
rect 2032 2890 3032 2916
rect 3090 2890 4090 2916
rect 4148 2890 5148 2916
rect 5206 2890 6206 2916
rect 6264 2890 7264 2916
rect 8546 2898 9546 2924
rect 9604 2898 10604 2924
rect 10662 2898 11662 2924
rect 11720 2898 12720 2924
rect 12778 2898 13778 2924
rect 15052 2906 16052 2932
rect 16110 2906 17110 2932
rect 17168 2906 18168 2932
rect 18226 2906 19226 2932
rect 19284 2906 20284 2932
rect 21542 2890 22542 2916
rect 22600 2890 23600 2916
rect 23658 2890 24658 2916
rect 24716 2890 25716 2916
rect 25774 2890 26774 2916
rect 28064 2906 29064 2932
rect 29122 2906 30122 2932
rect 30180 2906 31180 2932
rect 31238 2906 32238 2932
rect 32296 2906 33296 2932
rect 34574 2912 35574 2938
rect 35632 2912 36632 2938
rect 36690 2912 37690 2938
rect 37748 2912 38748 2938
rect 38806 2912 39806 2938
rect 41064 2912 42064 2938
rect 42122 2912 43122 2938
rect 43180 2912 44180 2938
rect 44238 2912 45238 2938
rect 45296 2912 46296 2938
rect 47652 2934 48652 2960
rect 48710 2934 49710 2960
rect 49768 2934 50768 2960
rect 50826 2934 51826 2960
rect 51884 2934 52884 2960
rect 54166 2948 55166 2974
rect 55224 2948 56224 2974
rect 56282 2948 57282 2974
rect 57340 2948 58340 2974
rect 58398 2948 59398 2974
rect 69354 26372 69558 26376
rect 69354 26368 69576 26372
rect 65526 26320 69576 26368
rect 80178 26340 81252 26704
rect 82510 26344 82714 26348
rect 82510 26340 82732 26344
rect 65526 26188 67586 26320
rect 68284 26188 69576 26320
rect 65526 26154 69576 26188
rect 65534 25990 66048 26154
rect 62608 25948 67234 25990
rect 69354 25988 69576 26154
rect 78682 26126 82732 26340
rect 95744 26336 95948 26340
rect 95744 26332 95966 26336
rect 62158 25942 67390 25948
rect 69070 25946 73696 25988
rect 78690 25962 79204 26126
rect 62158 25922 63158 25942
rect 63216 25922 64216 25942
rect 64274 25922 65274 25942
rect 65332 25922 66332 25942
rect 66390 25922 67390 25942
rect 68620 25940 73852 25946
rect 68620 25920 69620 25940
rect 69678 25920 70678 25940
rect 70736 25920 71736 25940
rect 71794 25920 72794 25940
rect 72852 25920 73852 25940
rect 75764 25920 80390 25962
rect 82510 25960 82732 26126
rect 91916 26288 95966 26332
rect 91916 26156 93994 26288
rect 94426 26156 95966 26288
rect 91916 26118 95966 26156
rect 62158 24896 63158 24922
rect 63216 24896 64216 24922
rect 64274 24896 65274 24922
rect 65332 24896 66332 24922
rect 66390 24896 67390 24922
rect 75314 25914 80546 25920
rect 82226 25918 86852 25960
rect 91924 25954 92438 26118
rect 75314 25894 76314 25914
rect 76372 25894 77372 25914
rect 77430 25894 78430 25914
rect 78488 25894 79488 25914
rect 79546 25894 80546 25914
rect 81776 25912 87008 25918
rect 88998 25912 93624 25954
rect 95744 25952 95966 26118
rect 62410 24854 62944 24896
rect 63448 24854 63982 24896
rect 64566 24854 65100 24896
rect 65582 24854 66116 24896
rect 66648 24854 67182 24896
rect 68620 24894 69620 24920
rect 69678 24894 70678 24920
rect 70736 24894 71736 24920
rect 71794 24894 72794 24920
rect 72852 24894 73852 24920
rect 81776 25892 82776 25912
rect 82834 25892 83834 25912
rect 83892 25892 84892 25912
rect 84950 25892 85950 25912
rect 86008 25892 87008 25912
rect 88548 25906 93780 25912
rect 95460 25910 100086 25952
rect 62158 24828 63158 24854
rect 63216 24828 64216 24854
rect 64274 24828 65274 24854
rect 65332 24828 66332 24854
rect 66390 24828 67390 24854
rect 68872 24852 69406 24894
rect 69910 24852 70444 24894
rect 71028 24852 71562 24894
rect 72044 24852 72578 24894
rect 73110 24852 73644 24894
rect 75314 24868 76314 24894
rect 76372 24868 77372 24894
rect 77430 24868 78430 24894
rect 78488 24868 79488 24894
rect 79546 24868 80546 24894
rect 88548 25886 89548 25906
rect 89606 25886 90606 25906
rect 90664 25886 91664 25906
rect 91722 25886 92722 25906
rect 92780 25886 93780 25906
rect 95010 25904 100242 25910
rect 68620 24826 69620 24852
rect 69678 24826 70678 24852
rect 70736 24826 71736 24852
rect 71794 24826 72794 24852
rect 72852 24826 73852 24852
rect 75566 24826 76100 24868
rect 76604 24826 77138 24868
rect 77722 24826 78256 24868
rect 78738 24826 79272 24868
rect 79804 24826 80338 24868
rect 81776 24866 82776 24892
rect 82834 24866 83834 24892
rect 83892 24866 84892 24892
rect 84950 24866 85950 24892
rect 86008 24866 87008 24892
rect 95010 25884 96010 25904
rect 96068 25884 97068 25904
rect 97126 25884 98126 25904
rect 98184 25884 99184 25904
rect 99242 25884 100242 25904
rect 62158 23802 63158 23828
rect 63216 23802 64216 23828
rect 64274 23802 65274 23828
rect 65332 23802 66332 23828
rect 66390 23802 67390 23828
rect 62446 23760 62980 23802
rect 63402 23760 63936 23802
rect 64510 23760 65044 23802
rect 65616 23760 66150 23802
rect 66646 23760 67180 23802
rect 62158 23734 63158 23760
rect 63216 23734 64216 23760
rect 64274 23734 65274 23760
rect 65332 23734 66332 23760
rect 66390 23734 67390 23760
rect 75314 24800 76314 24826
rect 76372 24800 77372 24826
rect 77430 24800 78430 24826
rect 78488 24800 79488 24826
rect 79546 24800 80546 24826
rect 82028 24824 82562 24866
rect 83066 24824 83600 24866
rect 84184 24824 84718 24866
rect 85200 24824 85734 24866
rect 86266 24824 86800 24866
rect 88548 24860 89548 24886
rect 89606 24860 90606 24886
rect 90664 24860 91664 24886
rect 91722 24860 92722 24886
rect 92780 24860 93780 24886
rect 68620 23800 69620 23826
rect 69678 23800 70678 23826
rect 70736 23800 71736 23826
rect 71794 23800 72794 23826
rect 72852 23800 73852 23826
rect 68908 23758 69442 23800
rect 69864 23758 70398 23800
rect 70972 23758 71506 23800
rect 72078 23758 72612 23800
rect 73108 23758 73642 23800
rect 68620 23732 69620 23758
rect 69678 23732 70678 23758
rect 70736 23732 71736 23758
rect 71794 23732 72794 23758
rect 72852 23732 73852 23758
rect 62158 22708 63158 22734
rect 63216 22708 64216 22734
rect 64274 22708 65274 22734
rect 65332 22708 66332 22734
rect 66390 22708 67390 22734
rect 62382 22666 62916 22708
rect 63436 22666 63970 22708
rect 64488 22666 65022 22708
rect 65596 22666 66130 22708
rect 66652 22666 67186 22708
rect 62158 22640 63158 22666
rect 63216 22640 64216 22666
rect 64274 22640 65274 22666
rect 65332 22640 66332 22666
rect 66390 22640 67390 22666
rect 81776 24798 82776 24824
rect 82834 24798 83834 24824
rect 83892 24798 84892 24824
rect 84950 24798 85950 24824
rect 86008 24798 87008 24824
rect 88800 24818 89334 24860
rect 89838 24818 90372 24860
rect 90956 24818 91490 24860
rect 91972 24818 92506 24860
rect 93038 24818 93572 24860
rect 95010 24858 96010 24884
rect 96068 24858 97068 24884
rect 97126 24858 98126 24884
rect 98184 24858 99184 24884
rect 99242 24858 100242 24884
rect 75314 23774 76314 23800
rect 76372 23774 77372 23800
rect 77430 23774 78430 23800
rect 78488 23774 79488 23800
rect 79546 23774 80546 23800
rect 75602 23732 76136 23774
rect 76558 23732 77092 23774
rect 77666 23732 78200 23774
rect 78772 23732 79306 23774
rect 79802 23732 80336 23774
rect 75314 23706 76314 23732
rect 76372 23706 77372 23732
rect 77430 23706 78430 23732
rect 78488 23706 79488 23732
rect 79546 23706 80546 23732
rect 68620 22706 69620 22732
rect 69678 22706 70678 22732
rect 70736 22706 71736 22732
rect 71794 22706 72794 22732
rect 72852 22706 73852 22732
rect 68844 22664 69378 22706
rect 69898 22664 70432 22706
rect 70950 22664 71484 22706
rect 72058 22664 72592 22706
rect 73114 22664 73648 22706
rect 68620 22638 69620 22664
rect 69678 22638 70678 22664
rect 70736 22638 71736 22664
rect 71794 22638 72794 22664
rect 72852 22638 73852 22664
rect 62158 21614 63158 21640
rect 63216 21614 64216 21640
rect 64274 21614 65274 21640
rect 65332 21614 66332 21640
rect 66390 21614 67390 21640
rect 88548 24792 89548 24818
rect 89606 24792 90606 24818
rect 90664 24792 91664 24818
rect 91722 24792 92722 24818
rect 92780 24792 93780 24818
rect 95262 24816 95796 24858
rect 96300 24816 96834 24858
rect 97418 24816 97952 24858
rect 98434 24816 98968 24858
rect 99500 24816 100034 24858
rect 81776 23772 82776 23798
rect 82834 23772 83834 23798
rect 83892 23772 84892 23798
rect 84950 23772 85950 23798
rect 86008 23772 87008 23798
rect 82064 23730 82598 23772
rect 83020 23730 83554 23772
rect 84128 23730 84662 23772
rect 85234 23730 85768 23772
rect 86264 23730 86798 23772
rect 81776 23704 82776 23730
rect 82834 23704 83834 23730
rect 83892 23704 84892 23730
rect 84950 23704 85950 23730
rect 86008 23704 87008 23730
rect 75314 22680 76314 22706
rect 76372 22680 77372 22706
rect 77430 22680 78430 22706
rect 78488 22680 79488 22706
rect 79546 22680 80546 22706
rect 75538 22638 76072 22680
rect 76592 22638 77126 22680
rect 77644 22638 78178 22680
rect 78752 22638 79286 22680
rect 79808 22638 80342 22680
rect 75314 22612 76314 22638
rect 76372 22612 77372 22638
rect 77430 22612 78430 22638
rect 78488 22612 79488 22638
rect 79546 22612 80546 22638
rect 62410 21572 62944 21614
rect 63508 21572 64042 21614
rect 64536 21572 65070 21614
rect 65500 21572 66034 21614
rect 66600 21572 67134 21614
rect 68620 21612 69620 21638
rect 69678 21612 70678 21638
rect 70736 21612 71736 21638
rect 71794 21612 72794 21638
rect 72852 21612 73852 21638
rect 95010 24790 96010 24816
rect 96068 24790 97068 24816
rect 97126 24790 98126 24816
rect 98184 24790 99184 24816
rect 99242 24790 100242 24816
rect 88548 23766 89548 23792
rect 89606 23766 90606 23792
rect 90664 23766 91664 23792
rect 91722 23766 92722 23792
rect 92780 23766 93780 23792
rect 88836 23724 89370 23766
rect 89792 23724 90326 23766
rect 90900 23724 91434 23766
rect 92006 23724 92540 23766
rect 93036 23724 93570 23766
rect 88548 23698 89548 23724
rect 89606 23698 90606 23724
rect 90664 23698 91664 23724
rect 91722 23698 92722 23724
rect 92780 23698 93780 23724
rect 81776 22678 82776 22704
rect 82834 22678 83834 22704
rect 83892 22678 84892 22704
rect 84950 22678 85950 22704
rect 86008 22678 87008 22704
rect 82000 22636 82534 22678
rect 83054 22636 83588 22678
rect 84106 22636 84640 22678
rect 85214 22636 85748 22678
rect 86270 22636 86804 22678
rect 81776 22610 82776 22636
rect 82834 22610 83834 22636
rect 83892 22610 84892 22636
rect 84950 22610 85950 22636
rect 86008 22610 87008 22636
rect 62158 21546 63158 21572
rect 63216 21546 64216 21572
rect 64274 21546 65274 21572
rect 65332 21546 66332 21572
rect 66390 21546 67390 21572
rect 68872 21570 69406 21612
rect 69970 21570 70504 21612
rect 70998 21570 71532 21612
rect 71962 21570 72496 21612
rect 73062 21570 73596 21612
rect 75314 21586 76314 21612
rect 76372 21586 77372 21612
rect 77430 21586 78430 21612
rect 78488 21586 79488 21612
rect 79546 21586 80546 21612
rect 95010 23764 96010 23790
rect 96068 23764 97068 23790
rect 97126 23764 98126 23790
rect 98184 23764 99184 23790
rect 99242 23764 100242 23790
rect 95298 23722 95832 23764
rect 96254 23722 96788 23764
rect 97362 23722 97896 23764
rect 98468 23722 99002 23764
rect 99498 23722 100032 23764
rect 95010 23696 96010 23722
rect 96068 23696 97068 23722
rect 97126 23696 98126 23722
rect 98184 23696 99184 23722
rect 99242 23696 100242 23722
rect 88548 22672 89548 22698
rect 89606 22672 90606 22698
rect 90664 22672 91664 22698
rect 91722 22672 92722 22698
rect 92780 22672 93780 22698
rect 88772 22630 89306 22672
rect 89826 22630 90360 22672
rect 90878 22630 91412 22672
rect 91986 22630 92520 22672
rect 93042 22630 93576 22672
rect 88548 22604 89548 22630
rect 89606 22604 90606 22630
rect 90664 22604 91664 22630
rect 91722 22604 92722 22630
rect 92780 22604 93780 22630
rect 68620 21544 69620 21570
rect 69678 21544 70678 21570
rect 70736 21544 71736 21570
rect 71794 21544 72794 21570
rect 72852 21544 73852 21570
rect 75566 21544 76100 21586
rect 76664 21544 77198 21586
rect 77692 21544 78226 21586
rect 78656 21544 79190 21586
rect 79756 21544 80290 21586
rect 81776 21584 82776 21610
rect 82834 21584 83834 21610
rect 83892 21584 84892 21610
rect 84950 21584 85950 21610
rect 86008 21584 87008 21610
rect 95010 22670 96010 22696
rect 96068 22670 97068 22696
rect 97126 22670 98126 22696
rect 98184 22670 99184 22696
rect 99242 22670 100242 22696
rect 95234 22628 95768 22670
rect 96288 22628 96822 22670
rect 97340 22628 97874 22670
rect 98448 22628 98982 22670
rect 99504 22628 100038 22670
rect 95010 22602 96010 22628
rect 96068 22602 97068 22628
rect 97126 22602 98126 22628
rect 98184 22602 99184 22628
rect 99242 22602 100242 22628
rect 62158 20520 63158 20546
rect 63216 20520 64216 20546
rect 64274 20520 65274 20546
rect 65332 20520 66332 20546
rect 66390 20520 67390 20546
rect 75314 21518 76314 21544
rect 76372 21518 77372 21544
rect 77430 21518 78430 21544
rect 78488 21518 79488 21544
rect 79546 21518 80546 21544
rect 82028 21542 82562 21584
rect 83126 21542 83660 21584
rect 84154 21542 84688 21584
rect 85118 21542 85652 21584
rect 86218 21542 86752 21584
rect 88548 21578 89548 21604
rect 89606 21578 90606 21604
rect 90664 21578 91664 21604
rect 91722 21578 92722 21604
rect 92780 21578 93780 21604
rect 62706 20152 63006 20520
rect 63568 20152 63868 20520
rect 64676 20152 64976 20520
rect 65630 20152 65930 20520
rect 66598 20152 66898 20520
rect 68620 20518 69620 20544
rect 69678 20518 70678 20544
rect 70736 20518 71736 20544
rect 71794 20518 72794 20544
rect 72852 20518 73852 20544
rect 81776 21516 82776 21542
rect 82834 21516 83834 21542
rect 83892 21516 84892 21542
rect 84950 21516 85950 21542
rect 86008 21516 87008 21542
rect 88800 21536 89334 21578
rect 89898 21536 90432 21578
rect 90926 21536 91460 21578
rect 91890 21536 92424 21578
rect 92990 21536 93524 21578
rect 95010 21576 96010 21602
rect 96068 21576 97068 21602
rect 97126 21576 98126 21602
rect 98184 21576 99184 21602
rect 99242 21576 100242 21602
rect 69122 20164 69390 20518
rect 69974 20164 70242 20518
rect 71194 20164 71462 20518
rect 72142 20164 72410 20518
rect 73070 20164 73338 20518
rect 75314 20492 76314 20518
rect 76372 20492 77372 20518
rect 77430 20492 78430 20518
rect 78488 20492 79488 20518
rect 79546 20492 80546 20518
rect 88548 21510 89548 21536
rect 89606 21510 90606 21536
rect 90664 21510 91664 21536
rect 91722 21510 92722 21536
rect 92780 21510 93780 21536
rect 95262 21534 95796 21576
rect 96360 21534 96894 21576
rect 97388 21534 97922 21576
rect 98352 21534 98886 21576
rect 99452 21534 99986 21576
rect 62614 20110 67240 20152
rect 69078 20122 73704 20164
rect 75862 20124 76162 20492
rect 76724 20124 77024 20492
rect 77832 20124 78132 20492
rect 78786 20124 79086 20492
rect 79754 20124 80054 20492
rect 81776 20490 82776 20516
rect 82834 20490 83834 20516
rect 83892 20490 84892 20516
rect 84950 20490 85950 20516
rect 86008 20490 87008 20516
rect 95010 21508 96010 21534
rect 96068 21508 97068 21534
rect 97126 21508 98126 21534
rect 98184 21508 99184 21534
rect 99242 21508 100242 21534
rect 82278 20136 82546 20490
rect 83130 20136 83398 20490
rect 84350 20136 84618 20490
rect 85298 20136 85566 20490
rect 86226 20136 86494 20490
rect 88548 20484 89548 20510
rect 89606 20484 90606 20510
rect 90664 20484 91664 20510
rect 91722 20484 92722 20510
rect 92780 20484 93780 20510
rect 68628 20116 73860 20122
rect 62164 20104 67396 20110
rect 62164 20084 63164 20104
rect 63222 20084 64222 20104
rect 64280 20084 65280 20104
rect 65338 20084 66338 20104
rect 66396 20084 67396 20104
rect 68628 20096 69628 20116
rect 69686 20096 70686 20116
rect 70744 20096 71744 20116
rect 71802 20096 72802 20116
rect 72860 20096 73860 20116
rect 75770 20082 80396 20124
rect 82234 20094 86860 20136
rect 89096 20116 89396 20484
rect 89958 20116 90258 20484
rect 91066 20116 91366 20484
rect 92020 20116 92320 20484
rect 92988 20116 93288 20484
rect 95010 20482 96010 20508
rect 96068 20482 97068 20508
rect 97126 20482 98126 20508
rect 98184 20482 99184 20508
rect 99242 20482 100242 20508
rect 95512 20128 95780 20482
rect 96364 20128 96632 20482
rect 97584 20128 97852 20482
rect 98532 20128 98800 20482
rect 99460 20128 99728 20482
rect 81784 20088 87016 20094
rect 75320 20076 80552 20082
rect 75320 20056 76320 20076
rect 76378 20056 77378 20076
rect 77436 20056 78436 20076
rect 78494 20056 79494 20076
rect 79552 20056 80552 20076
rect 81784 20068 82784 20088
rect 82842 20068 83842 20088
rect 83900 20068 84900 20088
rect 84958 20068 85958 20088
rect 86016 20068 87016 20088
rect 89004 20074 93630 20116
rect 95468 20086 100094 20128
rect 95018 20080 100250 20086
rect 88554 20068 93786 20074
rect 62164 19058 63164 19084
rect 63222 19058 64222 19084
rect 64280 19058 65280 19084
rect 65338 19058 66338 19084
rect 66396 19058 67396 19084
rect 68628 19070 69628 19096
rect 69686 19070 70686 19096
rect 70744 19070 71744 19096
rect 71802 19070 72802 19096
rect 72860 19070 73860 19096
rect 62416 19016 62950 19058
rect 63454 19016 63988 19058
rect 64572 19016 65106 19058
rect 65588 19016 66122 19058
rect 66654 19016 67188 19058
rect 68880 19028 69414 19070
rect 69918 19028 70452 19070
rect 71036 19028 71570 19070
rect 72052 19028 72586 19070
rect 73118 19028 73652 19070
rect 88554 20048 89554 20068
rect 89612 20048 90612 20068
rect 90670 20048 91670 20068
rect 91728 20048 92728 20068
rect 92786 20048 93786 20068
rect 95018 20060 96018 20080
rect 96076 20060 97076 20080
rect 97134 20060 98134 20080
rect 98192 20060 99192 20080
rect 99250 20060 100250 20080
rect 75320 19030 76320 19056
rect 76378 19030 77378 19056
rect 77436 19030 78436 19056
rect 78494 19030 79494 19056
rect 79552 19030 80552 19056
rect 81784 19042 82784 19068
rect 82842 19042 83842 19068
rect 83900 19042 84900 19068
rect 84958 19042 85958 19068
rect 86016 19042 87016 19068
rect 62164 18990 63164 19016
rect 63222 18990 64222 19016
rect 64280 18990 65280 19016
rect 65338 18990 66338 19016
rect 66396 18990 67396 19016
rect 68628 19002 69628 19028
rect 69686 19002 70686 19028
rect 70744 19002 71744 19028
rect 71802 19002 72802 19028
rect 72860 19002 73860 19028
rect 62164 17964 63164 17990
rect 63222 17964 64222 17990
rect 64280 17964 65280 17990
rect 65338 17964 66338 17990
rect 66396 17964 67396 17990
rect 62452 17922 62986 17964
rect 63408 17922 63942 17964
rect 64516 17922 65050 17964
rect 65622 17922 66156 17964
rect 66652 17922 67186 17964
rect 62164 17896 63164 17922
rect 63222 17896 64222 17922
rect 64280 17896 65280 17922
rect 65338 17896 66338 17922
rect 66396 17896 67396 17922
rect 75572 18988 76106 19030
rect 76610 18988 77144 19030
rect 77728 18988 78262 19030
rect 78744 18988 79278 19030
rect 79810 18988 80344 19030
rect 82036 19000 82570 19042
rect 83074 19000 83608 19042
rect 84192 19000 84726 19042
rect 85208 19000 85742 19042
rect 86274 19000 86808 19042
rect 88554 19022 89554 19048
rect 89612 19022 90612 19048
rect 90670 19022 91670 19048
rect 91728 19022 92728 19048
rect 92786 19022 93786 19048
rect 95018 19034 96018 19060
rect 96076 19034 97076 19060
rect 97134 19034 98134 19060
rect 98192 19034 99192 19060
rect 99250 19034 100250 19060
rect 75320 18962 76320 18988
rect 76378 18962 77378 18988
rect 77436 18962 78436 18988
rect 78494 18962 79494 18988
rect 79552 18962 80552 18988
rect 81784 18974 82784 19000
rect 82842 18974 83842 19000
rect 83900 18974 84900 19000
rect 84958 18974 85958 19000
rect 86016 18974 87016 19000
rect 88806 18980 89340 19022
rect 89844 18980 90378 19022
rect 90962 18980 91496 19022
rect 91978 18980 92512 19022
rect 93044 18980 93578 19022
rect 95270 18992 95804 19034
rect 96308 18992 96842 19034
rect 97426 18992 97960 19034
rect 98442 18992 98976 19034
rect 99508 18992 100042 19034
rect 68628 17976 69628 18002
rect 69686 17976 70686 18002
rect 70744 17976 71744 18002
rect 71802 17976 72802 18002
rect 72860 17976 73860 18002
rect 68916 17934 69450 17976
rect 69872 17934 70406 17976
rect 70980 17934 71514 17976
rect 72086 17934 72620 17976
rect 73116 17934 73650 17976
rect 68628 17908 69628 17934
rect 69686 17908 70686 17934
rect 70744 17908 71744 17934
rect 71802 17908 72802 17934
rect 72860 17908 73860 17934
rect 62164 16870 63164 16896
rect 63222 16870 64222 16896
rect 64280 16870 65280 16896
rect 65338 16870 66338 16896
rect 66396 16870 67396 16896
rect 62388 16828 62922 16870
rect 63442 16828 63976 16870
rect 64494 16828 65028 16870
rect 65602 16828 66136 16870
rect 66658 16828 67192 16870
rect 62164 16802 63164 16828
rect 63222 16802 64222 16828
rect 64280 16802 65280 16828
rect 65338 16802 66338 16828
rect 66396 16802 67396 16828
rect 75320 17936 76320 17962
rect 76378 17936 77378 17962
rect 77436 17936 78436 17962
rect 78494 17936 79494 17962
rect 79552 17936 80552 17962
rect 75608 17894 76142 17936
rect 76564 17894 77098 17936
rect 77672 17894 78206 17936
rect 78778 17894 79312 17936
rect 79808 17894 80342 17936
rect 75320 17868 76320 17894
rect 76378 17868 77378 17894
rect 77436 17868 78436 17894
rect 78494 17868 79494 17894
rect 79552 17868 80552 17894
rect 68628 16882 69628 16908
rect 69686 16882 70686 16908
rect 70744 16882 71744 16908
rect 71802 16882 72802 16908
rect 72860 16882 73860 16908
rect 68852 16840 69386 16882
rect 69906 16840 70440 16882
rect 70958 16840 71492 16882
rect 72066 16840 72600 16882
rect 73122 16840 73656 16882
rect 68628 16814 69628 16840
rect 69686 16814 70686 16840
rect 70744 16814 71744 16840
rect 71802 16814 72802 16840
rect 72860 16814 73860 16840
rect 88554 18954 89554 18980
rect 89612 18954 90612 18980
rect 90670 18954 91670 18980
rect 91728 18954 92728 18980
rect 92786 18954 93786 18980
rect 95018 18966 96018 18992
rect 96076 18966 97076 18992
rect 97134 18966 98134 18992
rect 98192 18966 99192 18992
rect 99250 18966 100250 18992
rect 81784 17948 82784 17974
rect 82842 17948 83842 17974
rect 83900 17948 84900 17974
rect 84958 17948 85958 17974
rect 86016 17948 87016 17974
rect 82072 17906 82606 17948
rect 83028 17906 83562 17948
rect 84136 17906 84670 17948
rect 85242 17906 85776 17948
rect 86272 17906 86806 17948
rect 81784 17880 82784 17906
rect 82842 17880 83842 17906
rect 83900 17880 84900 17906
rect 84958 17880 85958 17906
rect 86016 17880 87016 17906
rect 75320 16842 76320 16868
rect 76378 16842 77378 16868
rect 77436 16842 78436 16868
rect 78494 16842 79494 16868
rect 79552 16842 80552 16868
rect 75544 16800 76078 16842
rect 76598 16800 77132 16842
rect 77650 16800 78184 16842
rect 78758 16800 79292 16842
rect 79814 16800 80348 16842
rect 75320 16774 76320 16800
rect 76378 16774 77378 16800
rect 77436 16774 78436 16800
rect 78494 16774 79494 16800
rect 79552 16774 80552 16800
rect 62164 15776 63164 15802
rect 63222 15776 64222 15802
rect 64280 15776 65280 15802
rect 65338 15776 66338 15802
rect 66396 15776 67396 15802
rect 68628 15788 69628 15814
rect 69686 15788 70686 15814
rect 70744 15788 71744 15814
rect 71802 15788 72802 15814
rect 72860 15788 73860 15814
rect 62416 15734 62950 15776
rect 63514 15734 64048 15776
rect 64542 15734 65076 15776
rect 65506 15734 66040 15776
rect 66606 15734 67140 15776
rect 68880 15746 69414 15788
rect 69978 15746 70512 15788
rect 71006 15746 71540 15788
rect 71970 15746 72504 15788
rect 73070 15746 73604 15788
rect 88554 17928 89554 17954
rect 89612 17928 90612 17954
rect 90670 17928 91670 17954
rect 91728 17928 92728 17954
rect 92786 17928 93786 17954
rect 88842 17886 89376 17928
rect 89798 17886 90332 17928
rect 90906 17886 91440 17928
rect 92012 17886 92546 17928
rect 93042 17886 93576 17928
rect 88554 17860 89554 17886
rect 89612 17860 90612 17886
rect 90670 17860 91670 17886
rect 91728 17860 92728 17886
rect 92786 17860 93786 17886
rect 81784 16854 82784 16880
rect 82842 16854 83842 16880
rect 83900 16854 84900 16880
rect 84958 16854 85958 16880
rect 86016 16854 87016 16880
rect 82008 16812 82542 16854
rect 83062 16812 83596 16854
rect 84114 16812 84648 16854
rect 85222 16812 85756 16854
rect 86278 16812 86812 16854
rect 81784 16786 82784 16812
rect 82842 16786 83842 16812
rect 83900 16786 84900 16812
rect 84958 16786 85958 16812
rect 86016 16786 87016 16812
rect 95018 17940 96018 17966
rect 96076 17940 97076 17966
rect 97134 17940 98134 17966
rect 98192 17940 99192 17966
rect 99250 17940 100250 17966
rect 95306 17898 95840 17940
rect 96262 17898 96796 17940
rect 97370 17898 97904 17940
rect 98476 17898 99010 17940
rect 99506 17898 100040 17940
rect 95018 17872 96018 17898
rect 96076 17872 97076 17898
rect 97134 17872 98134 17898
rect 98192 17872 99192 17898
rect 99250 17872 100250 17898
rect 88554 16834 89554 16860
rect 89612 16834 90612 16860
rect 90670 16834 91670 16860
rect 91728 16834 92728 16860
rect 92786 16834 93786 16860
rect 88778 16792 89312 16834
rect 89832 16792 90366 16834
rect 90884 16792 91418 16834
rect 91992 16792 92526 16834
rect 93048 16792 93582 16834
rect 88554 16766 89554 16792
rect 89612 16766 90612 16792
rect 90670 16766 91670 16792
rect 91728 16766 92728 16792
rect 92786 16766 93786 16792
rect 75320 15748 76320 15774
rect 76378 15748 77378 15774
rect 77436 15748 78436 15774
rect 78494 15748 79494 15774
rect 79552 15748 80552 15774
rect 81784 15760 82784 15786
rect 82842 15760 83842 15786
rect 83900 15760 84900 15786
rect 84958 15760 85958 15786
rect 86016 15760 87016 15786
rect 95018 16846 96018 16872
rect 96076 16846 97076 16872
rect 97134 16846 98134 16872
rect 98192 16846 99192 16872
rect 99250 16846 100250 16872
rect 95242 16804 95776 16846
rect 96296 16804 96830 16846
rect 97348 16804 97882 16846
rect 98456 16804 98990 16846
rect 99512 16804 100046 16846
rect 95018 16778 96018 16804
rect 96076 16778 97076 16804
rect 97134 16778 98134 16804
rect 98192 16778 99192 16804
rect 99250 16778 100250 16804
rect 62164 15708 63164 15734
rect 63222 15708 64222 15734
rect 64280 15708 65280 15734
rect 65338 15708 66338 15734
rect 66396 15708 67396 15734
rect 68628 15720 69628 15746
rect 69686 15720 70686 15746
rect 70744 15720 71744 15746
rect 71802 15720 72802 15746
rect 72860 15720 73860 15746
rect 75572 15706 76106 15748
rect 76670 15706 77204 15748
rect 77698 15706 78232 15748
rect 78662 15706 79196 15748
rect 79762 15706 80296 15748
rect 82036 15718 82570 15760
rect 83134 15718 83668 15760
rect 84162 15718 84696 15760
rect 85126 15718 85660 15760
rect 86226 15718 86760 15760
rect 88554 15740 89554 15766
rect 89612 15740 90612 15766
rect 90670 15740 91670 15766
rect 91728 15740 92728 15766
rect 92786 15740 93786 15766
rect 95018 15752 96018 15778
rect 96076 15752 97076 15778
rect 97134 15752 98134 15778
rect 98192 15752 99192 15778
rect 99250 15752 100250 15778
rect 75320 15680 76320 15706
rect 76378 15680 77378 15706
rect 77436 15680 78436 15706
rect 78494 15680 79494 15706
rect 79552 15680 80552 15706
rect 81784 15692 82784 15718
rect 82842 15692 83842 15718
rect 83900 15692 84900 15718
rect 84958 15692 85958 15718
rect 86016 15692 87016 15718
rect 88806 15698 89340 15740
rect 89904 15698 90438 15740
rect 90932 15698 91466 15740
rect 91896 15698 92430 15740
rect 92996 15698 93530 15740
rect 95270 15710 95804 15752
rect 96368 15710 96902 15752
rect 97396 15710 97930 15752
rect 98360 15710 98894 15752
rect 99460 15710 99994 15752
rect 62164 14682 63164 14708
rect 63222 14682 64222 14708
rect 64280 14682 65280 14708
rect 65338 14682 66338 14708
rect 66396 14682 67396 14708
rect 68628 14694 69628 14720
rect 69686 14694 70686 14720
rect 70744 14694 71744 14720
rect 71802 14694 72802 14720
rect 72860 14694 73860 14720
rect 62718 14294 63026 14682
rect 63436 14294 63744 14682
rect 64794 14294 65102 14682
rect 65526 14294 65834 14682
rect 66630 14294 66938 14682
rect 62614 14252 67240 14294
rect 69138 14292 69428 14694
rect 69970 14292 70276 14694
rect 71012 14292 71318 14694
rect 72118 14292 72424 14694
rect 73194 14292 73500 14694
rect 88554 15672 89554 15698
rect 89612 15672 90612 15698
rect 90670 15672 91670 15698
rect 91728 15672 92728 15698
rect 92786 15672 93786 15698
rect 95018 15684 96018 15710
rect 96076 15684 97076 15710
rect 97134 15684 98134 15710
rect 98192 15684 99192 15710
rect 99250 15684 100250 15710
rect 75320 14654 76320 14680
rect 76378 14654 77378 14680
rect 77436 14654 78436 14680
rect 78494 14654 79494 14680
rect 79552 14654 80552 14680
rect 81784 14666 82784 14692
rect 82842 14666 83842 14692
rect 83900 14666 84900 14692
rect 84958 14666 85958 14692
rect 86016 14666 87016 14692
rect 62164 14246 67396 14252
rect 69082 14250 73708 14292
rect 75874 14266 76182 14654
rect 76592 14266 76900 14654
rect 77950 14266 78258 14654
rect 78682 14266 78990 14654
rect 79786 14266 80094 14654
rect 62164 14226 63164 14246
rect 63222 14226 64222 14246
rect 64280 14226 65280 14246
rect 65338 14226 66338 14246
rect 66396 14226 67396 14246
rect 68632 14244 73864 14250
rect 68632 14224 69632 14244
rect 69690 14224 70690 14244
rect 70748 14224 71748 14244
rect 71806 14224 72806 14244
rect 72864 14224 73864 14244
rect 75770 14224 80396 14266
rect 82294 14264 82584 14666
rect 83126 14264 83432 14666
rect 84168 14264 84474 14666
rect 85274 14264 85580 14666
rect 86350 14264 86656 14666
rect 88554 14646 89554 14672
rect 89612 14646 90612 14672
rect 90670 14646 91670 14672
rect 91728 14646 92728 14672
rect 92786 14646 93786 14672
rect 95018 14658 96018 14684
rect 96076 14658 97076 14684
rect 97134 14658 98134 14684
rect 98192 14658 99192 14684
rect 99250 14658 100250 14684
rect 62164 13200 63164 13226
rect 63222 13200 64222 13226
rect 64280 13200 65280 13226
rect 65338 13200 66338 13226
rect 66396 13200 67396 13226
rect 75320 14218 80552 14224
rect 82238 14222 86864 14264
rect 89108 14258 89416 14646
rect 89826 14258 90134 14646
rect 91184 14258 91492 14646
rect 91916 14258 92224 14646
rect 93020 14258 93328 14646
rect 75320 14198 76320 14218
rect 76378 14198 77378 14218
rect 77436 14198 78436 14218
rect 78494 14198 79494 14218
rect 79552 14198 80552 14218
rect 81788 14216 87020 14222
rect 89004 14216 93630 14258
rect 95528 14256 95818 14658
rect 96360 14256 96666 14658
rect 97402 14256 97708 14658
rect 98508 14256 98814 14658
rect 99584 14256 99890 14658
rect 62416 13158 62950 13200
rect 63454 13158 63988 13200
rect 64572 13158 65106 13200
rect 65588 13158 66122 13200
rect 66654 13158 67188 13200
rect 68632 13198 69632 13224
rect 69690 13198 70690 13224
rect 70748 13198 71748 13224
rect 71806 13198 72806 13224
rect 72864 13198 73864 13224
rect 81788 14196 82788 14216
rect 82846 14196 83846 14216
rect 83904 14196 84904 14216
rect 84962 14196 85962 14216
rect 86020 14196 87020 14216
rect 88554 14210 93786 14216
rect 95472 14214 100098 14256
rect 62164 13132 63164 13158
rect 63222 13132 64222 13158
rect 64280 13132 65280 13158
rect 65338 13132 66338 13158
rect 66396 13132 67396 13158
rect 68884 13156 69418 13198
rect 69922 13156 70456 13198
rect 71040 13156 71574 13198
rect 72056 13156 72590 13198
rect 73122 13156 73656 13198
rect 75320 13172 76320 13198
rect 76378 13172 77378 13198
rect 77436 13172 78436 13198
rect 78494 13172 79494 13198
rect 79552 13172 80552 13198
rect 88554 14190 89554 14210
rect 89612 14190 90612 14210
rect 90670 14190 91670 14210
rect 91728 14190 92728 14210
rect 92786 14190 93786 14210
rect 95022 14208 100254 14214
rect 68632 13130 69632 13156
rect 69690 13130 70690 13156
rect 70748 13130 71748 13156
rect 71806 13130 72806 13156
rect 72864 13130 73864 13156
rect 75572 13130 76106 13172
rect 76610 13130 77144 13172
rect 77728 13130 78262 13172
rect 78744 13130 79278 13172
rect 79810 13130 80344 13172
rect 81788 13170 82788 13196
rect 82846 13170 83846 13196
rect 83904 13170 84904 13196
rect 84962 13170 85962 13196
rect 86020 13170 87020 13196
rect 95022 14188 96022 14208
rect 96080 14188 97080 14208
rect 97138 14188 98138 14208
rect 98196 14188 99196 14208
rect 99254 14188 100254 14208
rect 62164 12106 63164 12132
rect 63222 12106 64222 12132
rect 64280 12106 65280 12132
rect 65338 12106 66338 12132
rect 66396 12106 67396 12132
rect 62452 12064 62986 12106
rect 63408 12064 63942 12106
rect 64516 12064 65050 12106
rect 65622 12064 66156 12106
rect 66652 12064 67186 12106
rect 62164 12038 63164 12064
rect 63222 12038 64222 12064
rect 64280 12038 65280 12064
rect 65338 12038 66338 12064
rect 66396 12038 67396 12064
rect 75320 13104 76320 13130
rect 76378 13104 77378 13130
rect 77436 13104 78436 13130
rect 78494 13104 79494 13130
rect 79552 13104 80552 13130
rect 82040 13128 82574 13170
rect 83078 13128 83612 13170
rect 84196 13128 84730 13170
rect 85212 13128 85746 13170
rect 86278 13128 86812 13170
rect 88554 13164 89554 13190
rect 89612 13164 90612 13190
rect 90670 13164 91670 13190
rect 91728 13164 92728 13190
rect 92786 13164 93786 13190
rect 68632 12104 69632 12130
rect 69690 12104 70690 12130
rect 70748 12104 71748 12130
rect 71806 12104 72806 12130
rect 72864 12104 73864 12130
rect 68920 12062 69454 12104
rect 69876 12062 70410 12104
rect 70984 12062 71518 12104
rect 72090 12062 72624 12104
rect 73120 12062 73654 12104
rect 68632 12036 69632 12062
rect 69690 12036 70690 12062
rect 70748 12036 71748 12062
rect 71806 12036 72806 12062
rect 72864 12036 73864 12062
rect 62164 11012 63164 11038
rect 63222 11012 64222 11038
rect 64280 11012 65280 11038
rect 65338 11012 66338 11038
rect 66396 11012 67396 11038
rect 62388 10970 62922 11012
rect 63442 10970 63976 11012
rect 64494 10970 65028 11012
rect 65602 10970 66136 11012
rect 66658 10970 67192 11012
rect 62164 10944 63164 10970
rect 63222 10944 64222 10970
rect 64280 10944 65280 10970
rect 65338 10944 66338 10970
rect 66396 10944 67396 10970
rect 81788 13102 82788 13128
rect 82846 13102 83846 13128
rect 83904 13102 84904 13128
rect 84962 13102 85962 13128
rect 86020 13102 87020 13128
rect 88806 13122 89340 13164
rect 89844 13122 90378 13164
rect 90962 13122 91496 13164
rect 91978 13122 92512 13164
rect 93044 13122 93578 13164
rect 95022 13162 96022 13188
rect 96080 13162 97080 13188
rect 97138 13162 98138 13188
rect 98196 13162 99196 13188
rect 99254 13162 100254 13188
rect 75320 12078 76320 12104
rect 76378 12078 77378 12104
rect 77436 12078 78436 12104
rect 78494 12078 79494 12104
rect 79552 12078 80552 12104
rect 75608 12036 76142 12078
rect 76564 12036 77098 12078
rect 77672 12036 78206 12078
rect 78778 12036 79312 12078
rect 79808 12036 80342 12078
rect 75320 12010 76320 12036
rect 76378 12010 77378 12036
rect 77436 12010 78436 12036
rect 78494 12010 79494 12036
rect 79552 12010 80552 12036
rect 68632 11010 69632 11036
rect 69690 11010 70690 11036
rect 70748 11010 71748 11036
rect 71806 11010 72806 11036
rect 72864 11010 73864 11036
rect 68856 10968 69390 11010
rect 69910 10968 70444 11010
rect 70962 10968 71496 11010
rect 72070 10968 72604 11010
rect 73126 10968 73660 11010
rect 68632 10942 69632 10968
rect 69690 10942 70690 10968
rect 70748 10942 71748 10968
rect 71806 10942 72806 10968
rect 72864 10942 73864 10968
rect 62164 9918 63164 9944
rect 63222 9918 64222 9944
rect 64280 9918 65280 9944
rect 65338 9918 66338 9944
rect 66396 9918 67396 9944
rect 88554 13096 89554 13122
rect 89612 13096 90612 13122
rect 90670 13096 91670 13122
rect 91728 13096 92728 13122
rect 92786 13096 93786 13122
rect 95274 13120 95808 13162
rect 96312 13120 96846 13162
rect 97430 13120 97964 13162
rect 98446 13120 98980 13162
rect 99512 13120 100046 13162
rect 81788 12076 82788 12102
rect 82846 12076 83846 12102
rect 83904 12076 84904 12102
rect 84962 12076 85962 12102
rect 86020 12076 87020 12102
rect 82076 12034 82610 12076
rect 83032 12034 83566 12076
rect 84140 12034 84674 12076
rect 85246 12034 85780 12076
rect 86276 12034 86810 12076
rect 81788 12008 82788 12034
rect 82846 12008 83846 12034
rect 83904 12008 84904 12034
rect 84962 12008 85962 12034
rect 86020 12008 87020 12034
rect 75320 10984 76320 11010
rect 76378 10984 77378 11010
rect 77436 10984 78436 11010
rect 78494 10984 79494 11010
rect 79552 10984 80552 11010
rect 75544 10942 76078 10984
rect 76598 10942 77132 10984
rect 77650 10942 78184 10984
rect 78758 10942 79292 10984
rect 79814 10942 80348 10984
rect 75320 10916 76320 10942
rect 76378 10916 77378 10942
rect 77436 10916 78436 10942
rect 78494 10916 79494 10942
rect 79552 10916 80552 10942
rect 62416 9876 62950 9918
rect 63514 9876 64048 9918
rect 64542 9876 65076 9918
rect 65506 9876 66040 9918
rect 66606 9876 67140 9918
rect 68632 9916 69632 9942
rect 69690 9916 70690 9942
rect 70748 9916 71748 9942
rect 71806 9916 72806 9942
rect 72864 9916 73864 9942
rect 95022 13094 96022 13120
rect 96080 13094 97080 13120
rect 97138 13094 98138 13120
rect 98196 13094 99196 13120
rect 99254 13094 100254 13120
rect 88554 12070 89554 12096
rect 89612 12070 90612 12096
rect 90670 12070 91670 12096
rect 91728 12070 92728 12096
rect 92786 12070 93786 12096
rect 88842 12028 89376 12070
rect 89798 12028 90332 12070
rect 90906 12028 91440 12070
rect 92012 12028 92546 12070
rect 93042 12028 93576 12070
rect 88554 12002 89554 12028
rect 89612 12002 90612 12028
rect 90670 12002 91670 12028
rect 91728 12002 92728 12028
rect 92786 12002 93786 12028
rect 81788 10982 82788 11008
rect 82846 10982 83846 11008
rect 83904 10982 84904 11008
rect 84962 10982 85962 11008
rect 86020 10982 87020 11008
rect 82012 10940 82546 10982
rect 83066 10940 83600 10982
rect 84118 10940 84652 10982
rect 85226 10940 85760 10982
rect 86282 10940 86816 10982
rect 81788 10914 82788 10940
rect 82846 10914 83846 10940
rect 83904 10914 84904 10940
rect 84962 10914 85962 10940
rect 86020 10914 87020 10940
rect 62164 9850 63164 9876
rect 63222 9850 64222 9876
rect 64280 9850 65280 9876
rect 65338 9850 66338 9876
rect 66396 9850 67396 9876
rect 68884 9874 69418 9916
rect 69982 9874 70516 9916
rect 71010 9874 71544 9916
rect 71974 9874 72508 9916
rect 73074 9874 73608 9916
rect 75320 9890 76320 9916
rect 76378 9890 77378 9916
rect 77436 9890 78436 9916
rect 78494 9890 79494 9916
rect 79552 9890 80552 9916
rect 95022 12068 96022 12094
rect 96080 12068 97080 12094
rect 97138 12068 98138 12094
rect 98196 12068 99196 12094
rect 99254 12068 100254 12094
rect 95310 12026 95844 12068
rect 96266 12026 96800 12068
rect 97374 12026 97908 12068
rect 98480 12026 99014 12068
rect 99510 12026 100044 12068
rect 95022 12000 96022 12026
rect 96080 12000 97080 12026
rect 97138 12000 98138 12026
rect 98196 12000 99196 12026
rect 99254 12000 100254 12026
rect 88554 10976 89554 11002
rect 89612 10976 90612 11002
rect 90670 10976 91670 11002
rect 91728 10976 92728 11002
rect 92786 10976 93786 11002
rect 88778 10934 89312 10976
rect 89832 10934 90366 10976
rect 90884 10934 91418 10976
rect 91992 10934 92526 10976
rect 93048 10934 93582 10976
rect 88554 10908 89554 10934
rect 89612 10908 90612 10934
rect 90670 10908 91670 10934
rect 91728 10908 92728 10934
rect 92786 10908 93786 10934
rect 68632 9848 69632 9874
rect 69690 9848 70690 9874
rect 70748 9848 71748 9874
rect 71806 9848 72806 9874
rect 72864 9848 73864 9874
rect 75572 9848 76106 9890
rect 76670 9848 77204 9890
rect 77698 9848 78232 9890
rect 78662 9848 79196 9890
rect 79762 9848 80296 9890
rect 81788 9888 82788 9914
rect 82846 9888 83846 9914
rect 83904 9888 84904 9914
rect 84962 9888 85962 9914
rect 86020 9888 87020 9914
rect 95022 10974 96022 11000
rect 96080 10974 97080 11000
rect 97138 10974 98138 11000
rect 98196 10974 99196 11000
rect 99254 10974 100254 11000
rect 95246 10932 95780 10974
rect 96300 10932 96834 10974
rect 97352 10932 97886 10974
rect 98460 10932 98994 10974
rect 99516 10932 100050 10974
rect 95022 10906 96022 10932
rect 96080 10906 97080 10932
rect 97138 10906 98138 10932
rect 98196 10906 99196 10932
rect 99254 10906 100254 10932
rect 62164 8824 63164 8850
rect 63222 8824 64222 8850
rect 64280 8824 65280 8850
rect 65338 8824 66338 8850
rect 66396 8824 67396 8850
rect 75320 9822 76320 9848
rect 76378 9822 77378 9848
rect 77436 9822 78436 9848
rect 78494 9822 79494 9848
rect 79552 9822 80552 9848
rect 82040 9846 82574 9888
rect 83138 9846 83672 9888
rect 84166 9846 84700 9888
rect 85130 9846 85664 9888
rect 86230 9846 86764 9888
rect 88554 9882 89554 9908
rect 89612 9882 90612 9908
rect 90670 9882 91670 9908
rect 91728 9882 92728 9908
rect 92786 9882 93786 9908
rect 62666 8436 62974 8824
rect 63504 8436 63812 8824
rect 64574 8436 64882 8824
rect 65622 8436 65930 8824
rect 66844 8436 67152 8824
rect 68632 8822 69632 8848
rect 69690 8822 70690 8848
rect 70748 8822 71748 8848
rect 71806 8822 72806 8848
rect 72864 8822 73864 8848
rect 81788 9820 82788 9846
rect 82846 9820 83846 9846
rect 83904 9820 84904 9846
rect 84962 9820 85962 9846
rect 86020 9820 87020 9846
rect 88806 9840 89340 9882
rect 89904 9840 90438 9882
rect 90932 9840 91466 9882
rect 91896 9840 92430 9882
rect 92996 9840 93530 9882
rect 95022 9880 96022 9906
rect 96080 9880 97080 9906
rect 97138 9880 98138 9906
rect 98196 9880 99196 9906
rect 99254 9880 100254 9906
rect 62614 8394 67240 8436
rect 69134 8434 69440 8822
rect 70100 8434 70406 8822
rect 70964 8434 71270 8822
rect 72126 8434 72432 8822
rect 73170 8434 73476 8822
rect 75320 8796 76320 8822
rect 76378 8796 77378 8822
rect 77436 8796 78436 8822
rect 78494 8796 79494 8822
rect 79552 8796 80552 8822
rect 88554 9814 89554 9840
rect 89612 9814 90612 9840
rect 90670 9814 91670 9840
rect 91728 9814 92728 9840
rect 92786 9814 93786 9840
rect 95274 9838 95808 9880
rect 96372 9838 96906 9880
rect 97400 9838 97934 9880
rect 98364 9838 98898 9880
rect 99464 9838 99998 9880
rect 62164 8388 67396 8394
rect 69086 8392 73712 8434
rect 75822 8408 76130 8796
rect 76660 8408 76968 8796
rect 77730 8408 78038 8796
rect 78778 8408 79086 8796
rect 80000 8408 80308 8796
rect 81788 8794 82788 8820
rect 82846 8794 83846 8820
rect 83904 8794 84904 8820
rect 84962 8794 85962 8820
rect 86020 8794 87020 8820
rect 95022 9812 96022 9838
rect 96080 9812 97080 9838
rect 97138 9812 98138 9838
rect 98196 9812 99196 9838
rect 99254 9812 100254 9838
rect 62164 8368 63164 8388
rect 63222 8368 64222 8388
rect 64280 8368 65280 8388
rect 65338 8368 66338 8388
rect 66396 8368 67396 8388
rect 68636 8386 73868 8392
rect 68636 8366 69636 8386
rect 69694 8366 70694 8386
rect 70752 8366 71752 8386
rect 71810 8366 72810 8386
rect 72868 8366 73868 8386
rect 75770 8366 80396 8408
rect 82290 8406 82596 8794
rect 83256 8406 83562 8794
rect 84120 8406 84426 8794
rect 85282 8406 85588 8794
rect 86326 8406 86632 8794
rect 88554 8788 89554 8814
rect 89612 8788 90612 8814
rect 90670 8788 91670 8814
rect 91728 8788 92728 8814
rect 92786 8788 93786 8814
rect 62164 7342 63164 7368
rect 63222 7342 64222 7368
rect 64280 7342 65280 7368
rect 65338 7342 66338 7368
rect 66396 7342 67396 7368
rect 75320 8360 80552 8366
rect 82242 8364 86868 8406
rect 89056 8400 89364 8788
rect 89894 8400 90202 8788
rect 90964 8400 91272 8788
rect 92012 8400 92320 8788
rect 93234 8400 93542 8788
rect 95022 8786 96022 8812
rect 96080 8786 97080 8812
rect 97138 8786 98138 8812
rect 98196 8786 99196 8812
rect 99254 8786 100254 8812
rect 75320 8340 76320 8360
rect 76378 8340 77378 8360
rect 77436 8340 78436 8360
rect 78494 8340 79494 8360
rect 79552 8340 80552 8360
rect 81792 8358 87024 8364
rect 89004 8358 93630 8400
rect 95524 8398 95830 8786
rect 96490 8398 96796 8786
rect 97354 8398 97660 8786
rect 98516 8398 98822 8786
rect 99560 8398 99866 8786
rect 62416 7300 62950 7342
rect 63454 7300 63988 7342
rect 64572 7300 65106 7342
rect 65588 7300 66122 7342
rect 66654 7300 67188 7342
rect 68636 7340 69636 7366
rect 69694 7340 70694 7366
rect 70752 7340 71752 7366
rect 71810 7340 72810 7366
rect 72868 7340 73868 7366
rect 81792 8338 82792 8358
rect 82850 8338 83850 8358
rect 83908 8338 84908 8358
rect 84966 8338 85966 8358
rect 86024 8338 87024 8358
rect 88554 8352 93786 8358
rect 95476 8356 100102 8398
rect 62164 7274 63164 7300
rect 63222 7274 64222 7300
rect 64280 7274 65280 7300
rect 65338 7274 66338 7300
rect 66396 7274 67396 7300
rect 68888 7298 69422 7340
rect 69926 7298 70460 7340
rect 71044 7298 71578 7340
rect 72060 7298 72594 7340
rect 73126 7298 73660 7340
rect 75320 7314 76320 7340
rect 76378 7314 77378 7340
rect 77436 7314 78436 7340
rect 78494 7314 79494 7340
rect 79552 7314 80552 7340
rect 88554 8332 89554 8352
rect 89612 8332 90612 8352
rect 90670 8332 91670 8352
rect 91728 8332 92728 8352
rect 92786 8332 93786 8352
rect 95026 8350 100258 8356
rect 68636 7272 69636 7298
rect 69694 7272 70694 7298
rect 70752 7272 71752 7298
rect 71810 7272 72810 7298
rect 72868 7272 73868 7298
rect 75572 7272 76106 7314
rect 76610 7272 77144 7314
rect 77728 7272 78262 7314
rect 78744 7272 79278 7314
rect 79810 7272 80344 7314
rect 81792 7312 82792 7338
rect 82850 7312 83850 7338
rect 83908 7312 84908 7338
rect 84966 7312 85966 7338
rect 86024 7312 87024 7338
rect 95026 8330 96026 8350
rect 96084 8330 97084 8350
rect 97142 8330 98142 8350
rect 98200 8330 99200 8350
rect 99258 8330 100258 8350
rect 62164 6248 63164 6274
rect 63222 6248 64222 6274
rect 64280 6248 65280 6274
rect 65338 6248 66338 6274
rect 66396 6248 67396 6274
rect 62452 6206 62986 6248
rect 63408 6206 63942 6248
rect 64516 6206 65050 6248
rect 65622 6206 66156 6248
rect 66652 6206 67186 6248
rect 62164 6180 63164 6206
rect 63222 6180 64222 6206
rect 64280 6180 65280 6206
rect 65338 6180 66338 6206
rect 66396 6180 67396 6206
rect 75320 7246 76320 7272
rect 76378 7246 77378 7272
rect 77436 7246 78436 7272
rect 78494 7246 79494 7272
rect 79552 7246 80552 7272
rect 82044 7270 82578 7312
rect 83082 7270 83616 7312
rect 84200 7270 84734 7312
rect 85216 7270 85750 7312
rect 86282 7270 86816 7312
rect 88554 7306 89554 7332
rect 89612 7306 90612 7332
rect 90670 7306 91670 7332
rect 91728 7306 92728 7332
rect 92786 7306 93786 7332
rect 68636 6246 69636 6272
rect 69694 6246 70694 6272
rect 70752 6246 71752 6272
rect 71810 6246 72810 6272
rect 72868 6246 73868 6272
rect 68924 6204 69458 6246
rect 69880 6204 70414 6246
rect 70988 6204 71522 6246
rect 72094 6204 72628 6246
rect 73124 6204 73658 6246
rect 68636 6178 69636 6204
rect 69694 6178 70694 6204
rect 70752 6178 71752 6204
rect 71810 6178 72810 6204
rect 72868 6178 73868 6204
rect 62164 5154 63164 5180
rect 63222 5154 64222 5180
rect 64280 5154 65280 5180
rect 65338 5154 66338 5180
rect 66396 5154 67396 5180
rect 62388 5112 62922 5154
rect 63442 5112 63976 5154
rect 64494 5112 65028 5154
rect 65602 5112 66136 5154
rect 66658 5112 67192 5154
rect 62164 5086 63164 5112
rect 63222 5086 64222 5112
rect 64280 5086 65280 5112
rect 65338 5086 66338 5112
rect 66396 5086 67396 5112
rect 81792 7244 82792 7270
rect 82850 7244 83850 7270
rect 83908 7244 84908 7270
rect 84966 7244 85966 7270
rect 86024 7244 87024 7270
rect 88806 7264 89340 7306
rect 89844 7264 90378 7306
rect 90962 7264 91496 7306
rect 91978 7264 92512 7306
rect 93044 7264 93578 7306
rect 95026 7304 96026 7330
rect 96084 7304 97084 7330
rect 97142 7304 98142 7330
rect 98200 7304 99200 7330
rect 99258 7304 100258 7330
rect 75320 6220 76320 6246
rect 76378 6220 77378 6246
rect 77436 6220 78436 6246
rect 78494 6220 79494 6246
rect 79552 6220 80552 6246
rect 75608 6178 76142 6220
rect 76564 6178 77098 6220
rect 77672 6178 78206 6220
rect 78778 6178 79312 6220
rect 79808 6178 80342 6220
rect 75320 6152 76320 6178
rect 76378 6152 77378 6178
rect 77436 6152 78436 6178
rect 78494 6152 79494 6178
rect 79552 6152 80552 6178
rect 68636 5152 69636 5178
rect 69694 5152 70694 5178
rect 70752 5152 71752 5178
rect 71810 5152 72810 5178
rect 72868 5152 73868 5178
rect 68860 5110 69394 5152
rect 69914 5110 70448 5152
rect 70966 5110 71500 5152
rect 72074 5110 72608 5152
rect 73130 5110 73664 5152
rect 68636 5084 69636 5110
rect 69694 5084 70694 5110
rect 70752 5084 71752 5110
rect 71810 5084 72810 5110
rect 72868 5084 73868 5110
rect 62164 4060 63164 4086
rect 63222 4060 64222 4086
rect 64280 4060 65280 4086
rect 65338 4060 66338 4086
rect 66396 4060 67396 4086
rect 88554 7238 89554 7264
rect 89612 7238 90612 7264
rect 90670 7238 91670 7264
rect 91728 7238 92728 7264
rect 92786 7238 93786 7264
rect 95278 7262 95812 7304
rect 96316 7262 96850 7304
rect 97434 7262 97968 7304
rect 98450 7262 98984 7304
rect 99516 7262 100050 7304
rect 81792 6218 82792 6244
rect 82850 6218 83850 6244
rect 83908 6218 84908 6244
rect 84966 6218 85966 6244
rect 86024 6218 87024 6244
rect 82080 6176 82614 6218
rect 83036 6176 83570 6218
rect 84144 6176 84678 6218
rect 85250 6176 85784 6218
rect 86280 6176 86814 6218
rect 81792 6150 82792 6176
rect 82850 6150 83850 6176
rect 83908 6150 84908 6176
rect 84966 6150 85966 6176
rect 86024 6150 87024 6176
rect 75320 5126 76320 5152
rect 76378 5126 77378 5152
rect 77436 5126 78436 5152
rect 78494 5126 79494 5152
rect 79552 5126 80552 5152
rect 75544 5084 76078 5126
rect 76598 5084 77132 5126
rect 77650 5084 78184 5126
rect 78758 5084 79292 5126
rect 79814 5084 80348 5126
rect 75320 5058 76320 5084
rect 76378 5058 77378 5084
rect 77436 5058 78436 5084
rect 78494 5058 79494 5084
rect 79552 5058 80552 5084
rect 62416 4018 62950 4060
rect 63514 4018 64048 4060
rect 64542 4018 65076 4060
rect 65506 4018 66040 4060
rect 66606 4018 67140 4060
rect 68636 4058 69636 4084
rect 69694 4058 70694 4084
rect 70752 4058 71752 4084
rect 71810 4058 72810 4084
rect 72868 4058 73868 4084
rect 95026 7236 96026 7262
rect 96084 7236 97084 7262
rect 97142 7236 98142 7262
rect 98200 7236 99200 7262
rect 99258 7236 100258 7262
rect 88554 6212 89554 6238
rect 89612 6212 90612 6238
rect 90670 6212 91670 6238
rect 91728 6212 92728 6238
rect 92786 6212 93786 6238
rect 88842 6170 89376 6212
rect 89798 6170 90332 6212
rect 90906 6170 91440 6212
rect 92012 6170 92546 6212
rect 93042 6170 93576 6212
rect 88554 6144 89554 6170
rect 89612 6144 90612 6170
rect 90670 6144 91670 6170
rect 91728 6144 92728 6170
rect 92786 6144 93786 6170
rect 81792 5124 82792 5150
rect 82850 5124 83850 5150
rect 83908 5124 84908 5150
rect 84966 5124 85966 5150
rect 86024 5124 87024 5150
rect 82016 5082 82550 5124
rect 83070 5082 83604 5124
rect 84122 5082 84656 5124
rect 85230 5082 85764 5124
rect 86286 5082 86820 5124
rect 81792 5056 82792 5082
rect 82850 5056 83850 5082
rect 83908 5056 84908 5082
rect 84966 5056 85966 5082
rect 86024 5056 87024 5082
rect 62164 3992 63164 4018
rect 63222 3992 64222 4018
rect 64280 3992 65280 4018
rect 65338 3992 66338 4018
rect 66396 3992 67396 4018
rect 68888 4016 69422 4058
rect 69986 4016 70520 4058
rect 71014 4016 71548 4058
rect 71978 4016 72512 4058
rect 73078 4016 73612 4058
rect 75320 4032 76320 4058
rect 76378 4032 77378 4058
rect 77436 4032 78436 4058
rect 78494 4032 79494 4058
rect 79552 4032 80552 4058
rect 95026 6210 96026 6236
rect 96084 6210 97084 6236
rect 97142 6210 98142 6236
rect 98200 6210 99200 6236
rect 99258 6210 100258 6236
rect 95314 6168 95848 6210
rect 96270 6168 96804 6210
rect 97378 6168 97912 6210
rect 98484 6168 99018 6210
rect 99514 6168 100048 6210
rect 95026 6142 96026 6168
rect 96084 6142 97084 6168
rect 97142 6142 98142 6168
rect 98200 6142 99200 6168
rect 99258 6142 100258 6168
rect 88554 5118 89554 5144
rect 89612 5118 90612 5144
rect 90670 5118 91670 5144
rect 91728 5118 92728 5144
rect 92786 5118 93786 5144
rect 88778 5076 89312 5118
rect 89832 5076 90366 5118
rect 90884 5076 91418 5118
rect 91992 5076 92526 5118
rect 93048 5076 93582 5118
rect 88554 5050 89554 5076
rect 89612 5050 90612 5076
rect 90670 5050 91670 5076
rect 91728 5050 92728 5076
rect 92786 5050 93786 5076
rect 68636 3990 69636 4016
rect 69694 3990 70694 4016
rect 70752 3990 71752 4016
rect 71810 3990 72810 4016
rect 72868 3990 73868 4016
rect 75572 3990 76106 4032
rect 76670 3990 77204 4032
rect 77698 3990 78232 4032
rect 78662 3990 79196 4032
rect 79762 3990 80296 4032
rect 81792 4030 82792 4056
rect 82850 4030 83850 4056
rect 83908 4030 84908 4056
rect 84966 4030 85966 4056
rect 86024 4030 87024 4056
rect 95026 5116 96026 5142
rect 96084 5116 97084 5142
rect 97142 5116 98142 5142
rect 98200 5116 99200 5142
rect 99258 5116 100258 5142
rect 95250 5074 95784 5116
rect 96304 5074 96838 5116
rect 97356 5074 97890 5116
rect 98464 5074 98998 5116
rect 99520 5074 100054 5116
rect 95026 5048 96026 5074
rect 96084 5048 97084 5074
rect 97142 5048 98142 5074
rect 98200 5048 99200 5074
rect 99258 5048 100258 5074
rect 62164 2966 63164 2992
rect 63222 2966 64222 2992
rect 64280 2966 65280 2992
rect 65338 2966 66338 2992
rect 66396 2966 67396 2992
rect 75320 3964 76320 3990
rect 76378 3964 77378 3990
rect 77436 3964 78436 3990
rect 78494 3964 79494 3990
rect 79552 3964 80552 3990
rect 82044 3988 82578 4030
rect 83142 3988 83676 4030
rect 84170 3988 84704 4030
rect 85134 3988 85668 4030
rect 86234 3988 86768 4030
rect 88554 4024 89554 4050
rect 89612 4024 90612 4050
rect 90670 4024 91670 4050
rect 91728 4024 92728 4050
rect 92786 4024 93786 4050
rect 68636 2964 69636 2990
rect 69694 2964 70694 2990
rect 70752 2964 71752 2990
rect 71810 2964 72810 2990
rect 72868 2964 73868 2990
rect 81792 3962 82792 3988
rect 82850 3962 83850 3988
rect 83908 3962 84908 3988
rect 84966 3962 85966 3988
rect 86024 3962 87024 3988
rect 88806 3982 89340 4024
rect 89904 3982 90438 4024
rect 90932 3982 91466 4024
rect 91896 3982 92430 4024
rect 92996 3982 93530 4024
rect 95026 4022 96026 4048
rect 96084 4022 97084 4048
rect 97142 4022 98142 4048
rect 98200 4022 99200 4048
rect 99258 4022 100258 4048
rect 75320 2938 76320 2964
rect 76378 2938 77378 2964
rect 77436 2938 78436 2964
rect 78494 2938 79494 2964
rect 79552 2938 80552 2964
rect 88554 3956 89554 3982
rect 89612 3956 90612 3982
rect 90670 3956 91670 3982
rect 91728 3956 92728 3982
rect 92786 3956 93786 3982
rect 95278 3980 95812 4022
rect 96376 3980 96910 4022
rect 97404 3980 97938 4022
rect 98368 3980 98902 4022
rect 99468 3980 100002 4022
rect 81792 2936 82792 2962
rect 82850 2936 83850 2962
rect 83908 2936 84908 2962
rect 84966 2936 85966 2962
rect 86024 2936 87024 2962
rect 95026 3954 96026 3980
rect 96084 3954 97084 3980
rect 97142 3954 98142 3980
rect 98200 3954 99200 3980
rect 99258 3954 100258 3980
rect 88554 2930 89554 2956
rect 89612 2930 90612 2956
rect 90670 2930 91670 2956
rect 91728 2930 92728 2956
rect 92786 2930 93786 2956
rect 95026 2928 96026 2954
rect 96084 2928 97084 2954
rect 97142 2928 98142 2954
rect 98200 2928 99200 2954
rect 99258 2928 100258 2954
<< polycont >>
rect 72590 74370 72878 74496
rect 80390 74406 80836 74590
rect 57710 69438 57854 69722
rect 20714 64054 20798 64128
rect 20678 54424 20792 54660
rect 20678 48690 20750 48742
rect 41814 64098 42072 64334
rect 57780 60506 57972 61190
rect 30340 56768 30394 56854
rect 23294 54418 23382 54734
rect 30374 52928 30470 53076
rect 57626 51974 57772 52376
rect 83536 53723 83570 53757
rect 83536 53655 83570 53689
rect 83400 53587 83434 53621
rect 83400 53519 83434 53553
rect 84123 53818 84157 53852
rect 84284 53818 84318 53852
rect 83827 53676 83861 53710
rect 83827 53608 83861 53642
rect 83971 53639 84005 53673
rect 83971 53571 84005 53605
rect 84456 53702 84490 53736
rect 84283 53633 84317 53667
rect 84283 53565 84317 53599
rect 84456 53634 84490 53668
rect 84609 53633 84643 53667
rect 85088 53729 85122 53763
rect 85088 53661 85122 53695
rect 85213 53705 85247 53739
rect 85449 53630 85483 53664
rect 84844 53563 84878 53597
rect 85281 53569 85315 53603
rect 85281 53501 85315 53535
rect 85449 53562 85483 53596
rect 85721 53705 85755 53739
rect 85579 53565 85613 53599
rect 85579 53497 85613 53531
rect 86166 53619 86200 53653
rect 77348 50826 77656 51022
rect 11050 43606 11240 43736
rect 49550 43672 49974 43936
rect 63810 43466 64200 43632
rect 67818 43438 68110 43584
rect 71596 43444 71844 43614
rect 78536 39406 78796 39510
rect 80866 39410 81116 39538
rect 85060 39412 85316 39524
rect 67586 26188 68284 26320
rect 93994 26156 94426 26288
<< locali >>
rect 80314 74590 80914 74608
rect 72564 74496 72908 74538
rect 72564 74370 72590 74496
rect 72878 74370 72908 74496
rect 72564 74328 72908 74370
rect 80314 74406 80390 74590
rect 80836 74406 80914 74590
rect 80314 74366 80914 74406
rect 72628 74210 72754 74328
rect 73954 74210 74030 74214
rect 71328 74206 74030 74210
rect 71324 74108 74030 74206
rect 80346 74204 80444 74212
rect 80514 74204 80648 74366
rect 81668 74204 81744 74208
rect 79042 74200 81744 74204
rect 76496 74190 76594 74198
rect 77818 74190 77894 74194
rect 75192 74186 77894 74190
rect 71324 74040 71378 74108
rect 72628 74106 72754 74108
rect 71324 73870 71338 74040
rect 71296 73868 71338 73870
rect 71372 73870 71378 74040
rect 71996 74040 72030 74056
rect 71372 73868 71388 73870
rect 42754 73732 45400 73768
rect 42754 73400 42904 73732
rect 45304 73400 45400 73732
rect 42754 73366 45400 73400
rect 46762 73730 49408 73766
rect 46762 73398 46912 73730
rect 49312 73398 49408 73730
rect 46762 73364 49408 73398
rect 50774 73730 53420 73766
rect 50774 73398 50924 73730
rect 53324 73398 53420 73730
rect 50774 73364 53420 73398
rect 54784 73730 57430 73766
rect 54784 73398 54934 73730
rect 57334 73398 57430 73730
rect 54784 73364 57430 73398
rect 71296 73274 71388 73868
rect 71968 73868 71996 73926
rect 72632 74040 72730 74106
rect 72632 73990 72654 74040
rect 72030 73868 72046 73926
rect 71968 73790 72046 73868
rect 72688 73990 72730 74040
rect 73276 74040 73400 74108
rect 73276 73994 73312 74040
rect 73286 73896 73312 73916
rect 72654 73852 72688 73868
rect 73262 73868 73312 73896
rect 73346 73994 73400 74040
rect 73954 74040 74030 74108
rect 73954 73964 73970 74040
rect 73346 73882 73364 73916
rect 73346 73868 73368 73882
rect 73262 73792 73368 73868
rect 74004 73964 74030 74040
rect 75188 74088 77894 74186
rect 75188 74020 75242 74088
rect 73970 73852 74004 73868
rect 75188 73850 75202 74020
rect 73148 73790 73368 73792
rect 71968 73714 73368 73790
rect 71968 73712 73164 73714
rect 71980 73710 73164 73712
rect 73288 73706 73368 73714
rect 75160 73848 75202 73850
rect 75236 73850 75242 74020
rect 75860 74020 75894 74036
rect 75236 73848 75252 73850
rect 73932 73282 74110 73292
rect 73924 73274 74110 73282
rect 45286 73244 45550 73258
rect 49294 73244 49558 73256
rect 53306 73244 53570 73256
rect 57316 73244 57580 73256
rect 42468 73228 57580 73244
rect 71292 73232 74110 73274
rect 75160 73254 75252 73848
rect 75832 73848 75860 73906
rect 76496 74020 76594 74088
rect 76496 73970 76518 74020
rect 75894 73848 75910 73906
rect 75832 73770 75910 73848
rect 76552 73970 76594 74020
rect 77176 74020 77210 74036
rect 77150 73876 77176 73896
rect 76518 73832 76552 73848
rect 77126 73848 77176 73876
rect 77818 74020 77894 74088
rect 77818 73944 77834 74020
rect 77210 73862 77228 73896
rect 77210 73848 77232 73862
rect 77126 73772 77232 73848
rect 77868 73944 77894 74020
rect 79038 74102 81744 74200
rect 79038 74034 79092 74102
rect 79038 73864 79052 74034
rect 77834 73832 77868 73848
rect 79010 73862 79052 73864
rect 79086 73864 79092 74034
rect 79710 74034 79744 74050
rect 79086 73862 79102 73864
rect 77012 73770 77232 73772
rect 75832 73694 77232 73770
rect 75832 73692 77028 73694
rect 75844 73690 77028 73692
rect 77152 73686 77232 73694
rect 77796 73262 77974 73272
rect 79010 73268 79102 73862
rect 79682 73862 79710 73920
rect 80346 74034 80444 74102
rect 80514 74096 80648 74102
rect 80346 73984 80368 74034
rect 79744 73862 79760 73920
rect 79682 73784 79760 73862
rect 80402 73984 80444 74034
rect 80996 74034 81090 74102
rect 80996 73976 81026 74034
rect 81000 73890 81026 73910
rect 80368 73846 80402 73862
rect 80976 73862 81026 73890
rect 81060 73976 81090 74034
rect 81668 74034 81744 74102
rect 81668 73958 81684 74034
rect 81060 73876 81078 73910
rect 81060 73862 81082 73876
rect 80976 73786 81082 73862
rect 81718 73958 81744 74034
rect 81684 73846 81718 73862
rect 80862 73784 81082 73786
rect 79682 73708 81082 73784
rect 79682 73706 80878 73708
rect 79694 73704 80878 73706
rect 81002 73700 81082 73708
rect 81646 73276 81824 73286
rect 81638 73268 81824 73276
rect 77788 73254 77974 73262
rect 42394 73194 42410 73228
rect 42582 73194 43104 73228
rect 43276 73194 43798 73228
rect 43970 73194 44492 73228
rect 44664 73194 45186 73228
rect 45358 73226 57580 73228
rect 45358 73194 46418 73226
rect 42468 73192 46418 73194
rect 46590 73192 47112 73226
rect 47284 73192 47806 73226
rect 47978 73192 48500 73226
rect 48672 73192 49194 73226
rect 49366 73192 50430 73226
rect 50602 73192 51124 73226
rect 51296 73192 51818 73226
rect 51990 73192 52512 73226
rect 52684 73192 53206 73226
rect 53378 73192 54440 73226
rect 54612 73192 55134 73226
rect 55306 73192 55828 73226
rect 56000 73192 56522 73226
rect 56694 73192 57216 73226
rect 57388 73192 57580 73226
rect 42484 73186 45550 73192
rect 45286 73182 45550 73186
rect 46492 73184 49558 73192
rect 50504 73184 53570 73192
rect 54514 73184 57580 73192
rect 42232 72582 42518 72596
rect 42232 72570 45368 72582
rect 42232 72536 42410 72570
rect 42582 72536 43104 72570
rect 43276 72536 43798 72570
rect 43970 72536 44492 72570
rect 44664 72536 45186 72570
rect 45358 72536 45374 72570
rect 42232 72528 45368 72536
rect 42232 72520 42518 72528
rect 42232 71274 42314 72520
rect 45472 71930 45526 73182
rect 49294 73180 49558 73184
rect 53306 73180 53570 73184
rect 57316 73180 57580 73184
rect 46240 72580 46526 72594
rect 46240 72568 49376 72580
rect 46240 72534 46418 72568
rect 46590 72534 47112 72568
rect 47284 72534 47806 72568
rect 47978 72534 48500 72568
rect 48672 72534 49194 72568
rect 49366 72534 49382 72568
rect 46240 72526 49376 72534
rect 46240 72518 46526 72526
rect 45322 71924 45586 71930
rect 42532 71912 45586 71924
rect 42394 71878 42410 71912
rect 42582 71878 43104 71912
rect 43276 71878 43798 71912
rect 43970 71878 44492 71912
rect 44664 71878 45186 71912
rect 45358 71878 45586 71912
rect 42532 71870 45586 71878
rect 45322 71854 45586 71870
rect 42228 71266 42548 71274
rect 42228 71254 45376 71266
rect 42228 71220 42410 71254
rect 42582 71220 43104 71254
rect 43276 71220 43798 71254
rect 43970 71220 44492 71254
rect 44664 71220 45186 71254
rect 45358 71220 45376 71254
rect 42228 71212 45376 71220
rect 42228 71198 42548 71212
rect 42232 69974 42314 71198
rect 45472 70616 45526 71854
rect 46240 71272 46322 72518
rect 49480 71928 49534 73180
rect 50252 72580 50538 72594
rect 50252 72568 53388 72580
rect 50252 72534 50430 72568
rect 50602 72534 51124 72568
rect 51296 72534 51818 72568
rect 51990 72534 52512 72568
rect 52684 72534 53206 72568
rect 53378 72534 53394 72568
rect 50252 72526 53388 72534
rect 50252 72518 50538 72526
rect 49330 71922 49594 71928
rect 46540 71910 49594 71922
rect 46402 71876 46418 71910
rect 46590 71876 47112 71910
rect 47284 71876 47806 71910
rect 47978 71876 48500 71910
rect 48672 71876 49194 71910
rect 49366 71876 49594 71910
rect 46540 71868 49594 71876
rect 49330 71852 49594 71868
rect 46236 71264 46556 71272
rect 46236 71252 49384 71264
rect 46236 71218 46418 71252
rect 46590 71218 47112 71252
rect 47284 71218 47806 71252
rect 47978 71218 48500 71252
rect 48672 71218 49194 71252
rect 49366 71218 49384 71252
rect 46236 71210 49384 71218
rect 46236 71196 46556 71210
rect 45292 70602 45556 70616
rect 42530 70596 45556 70602
rect 42394 70562 42410 70596
rect 42582 70562 43104 70596
rect 43276 70562 43798 70596
rect 43970 70562 44492 70596
rect 44664 70562 45186 70596
rect 45358 70562 45556 70596
rect 42530 70548 45556 70562
rect 45292 70540 45556 70548
rect 45472 70538 45526 70540
rect 42214 69968 42314 69974
rect 42214 69958 42528 69968
rect 46240 69966 46322 71196
rect 49480 70614 49534 71852
rect 50252 71272 50334 72518
rect 53492 71928 53546 73180
rect 54262 72580 54548 72594
rect 54262 72568 57398 72580
rect 54262 72534 54440 72568
rect 54612 72534 55134 72568
rect 55306 72534 55828 72568
rect 56000 72534 56522 72568
rect 56694 72534 57216 72568
rect 57388 72534 57404 72568
rect 54262 72526 57398 72534
rect 54262 72518 54548 72526
rect 53342 71922 53606 71928
rect 50552 71910 53606 71922
rect 50414 71876 50430 71910
rect 50602 71876 51124 71910
rect 51296 71876 51818 71910
rect 51990 71876 52512 71910
rect 52684 71876 53206 71910
rect 53378 71876 53606 71910
rect 50552 71868 53606 71876
rect 53342 71852 53606 71868
rect 50248 71264 50568 71272
rect 50248 71252 53396 71264
rect 50248 71218 50430 71252
rect 50602 71218 51124 71252
rect 51296 71218 51818 71252
rect 51990 71218 52512 71252
rect 52684 71218 53206 71252
rect 53378 71218 53396 71252
rect 50248 71210 53396 71218
rect 50248 71196 50568 71210
rect 49300 70600 49564 70614
rect 46538 70594 49564 70600
rect 46402 70560 46418 70594
rect 46590 70560 47112 70594
rect 47284 70560 47806 70594
rect 47978 70560 48500 70594
rect 48672 70560 49194 70594
rect 49366 70560 49564 70594
rect 46538 70546 49564 70560
rect 49300 70538 49564 70546
rect 49480 70536 49534 70538
rect 50252 69966 50334 71196
rect 53492 70614 53546 71852
rect 54262 71272 54344 72518
rect 57502 71928 57556 73180
rect 71296 73126 71352 73232
rect 71012 73066 71228 73126
rect 57352 71922 57616 71928
rect 54562 71910 57616 71922
rect 54424 71876 54440 71910
rect 54612 71876 55134 71910
rect 55306 71876 55828 71910
rect 56000 71876 56522 71910
rect 56694 71876 57216 71910
rect 57388 71876 57616 71910
rect 54562 71868 57616 71876
rect 57352 71852 57616 71868
rect 54258 71264 54578 71272
rect 54258 71252 57406 71264
rect 54258 71218 54440 71252
rect 54612 71218 55134 71252
rect 55306 71218 55828 71252
rect 56000 71218 56522 71252
rect 56694 71218 57216 71252
rect 57388 71218 57406 71252
rect 54258 71210 57406 71218
rect 54258 71196 54578 71210
rect 53312 70600 53576 70614
rect 50550 70594 53576 70600
rect 50414 70560 50430 70594
rect 50602 70560 51124 70594
rect 51296 70560 51818 70594
rect 51990 70560 52512 70594
rect 52684 70560 53206 70594
rect 53378 70560 53576 70594
rect 50550 70546 53576 70560
rect 53312 70538 53576 70546
rect 53492 70536 53546 70538
rect 54262 69966 54344 71196
rect 57502 70614 57556 71852
rect 57322 70600 57586 70614
rect 54560 70594 57586 70600
rect 54424 70560 54440 70594
rect 54612 70560 55134 70594
rect 55306 70560 55828 70594
rect 56000 70560 56522 70594
rect 56694 70560 57216 70594
rect 57388 70560 57586 70594
rect 54560 70546 57586 70560
rect 57322 70538 57586 70546
rect 46236 69958 46536 69966
rect 50248 69958 50548 69966
rect 54258 69958 54558 69966
rect 42214 69946 57274 69958
rect 42214 69938 57400 69946
rect 42214 69904 42410 69938
rect 42582 69904 43104 69938
rect 43276 69904 43798 69938
rect 43970 69904 44492 69938
rect 44664 69904 45186 69938
rect 45358 69936 57400 69938
rect 45358 69906 46418 69936
rect 45358 69904 45374 69906
rect 42214 69894 45370 69904
rect 46236 69902 46418 69906
rect 46590 69902 47112 69936
rect 47284 69902 47806 69936
rect 47978 69902 48500 69936
rect 48672 69902 49194 69936
rect 49366 69906 50430 69936
rect 49366 69902 49382 69906
rect 50248 69902 50430 69906
rect 50602 69902 51124 69936
rect 51296 69902 51818 69936
rect 51990 69902 52512 69936
rect 52684 69902 53206 69936
rect 53378 69906 54440 69936
rect 53378 69902 53394 69906
rect 54258 69902 54440 69906
rect 54612 69902 55134 69936
rect 55306 69902 55828 69936
rect 56000 69902 56522 69936
rect 56694 69902 57216 69936
rect 57388 69902 57404 69936
rect 42214 69892 42510 69894
rect 46236 69892 49378 69902
rect 50248 69892 53390 69902
rect 54258 69892 57400 69902
rect 42214 69890 42314 69892
rect 46236 69890 46518 69892
rect 50248 69890 50530 69892
rect 54258 69890 54540 69892
rect 42214 68398 42296 69890
rect 46240 69888 46322 69890
rect 50252 69888 50334 69890
rect 54262 69888 54344 69890
rect 57498 69648 57584 70538
rect 71012 70320 71042 73066
rect 71182 72724 71228 73066
rect 71296 72954 71310 73126
rect 71344 72954 71352 73126
rect 71968 73126 72002 73142
rect 71296 72724 71352 72954
rect 71182 72630 71352 72724
rect 71182 70320 71228 72630
rect 71012 70266 71228 70320
rect 71296 72432 71352 72630
rect 71296 72260 71310 72432
rect 71344 72260 71352 72432
rect 71296 71738 71352 72260
rect 71296 71566 71310 71738
rect 71344 71566 71352 71738
rect 71296 71044 71352 71566
rect 71296 70872 71310 71044
rect 71344 70872 71352 71044
rect 71296 70350 71352 70872
rect 71296 70302 71310 70350
rect 71284 70178 71310 70302
rect 71344 70278 71352 70350
rect 71958 72954 71968 73110
rect 72614 73126 72670 73232
rect 73924 73222 74110 73232
rect 72002 72954 72014 73110
rect 72614 73106 72626 73126
rect 71958 72432 72014 72954
rect 71958 72260 71968 72432
rect 72002 72260 72014 72432
rect 71958 71738 72014 72260
rect 71958 71566 71968 71738
rect 72002 71566 72014 71738
rect 71958 71044 72014 71566
rect 71958 70872 71968 71044
rect 72002 70872 72014 71044
rect 71958 70350 72014 70872
rect 71958 70310 71968 70350
rect 71344 70178 71350 70278
rect 57692 69722 57870 69752
rect 57692 69648 57710 69722
rect 42746 69534 45392 69570
rect 42746 69202 42896 69534
rect 45296 69202 45392 69534
rect 42746 69168 45392 69202
rect 46740 69534 49386 69570
rect 46740 69202 46890 69534
rect 49290 69202 49386 69534
rect 46740 69168 49386 69202
rect 50762 69534 53408 69570
rect 50762 69202 50912 69534
rect 53312 69202 53408 69534
rect 50762 69168 53408 69202
rect 54784 69534 57430 69570
rect 54784 69202 54934 69534
rect 57334 69202 57430 69534
rect 54784 69168 57430 69202
rect 57498 69514 57710 69648
rect 57498 69060 57584 69514
rect 57692 69438 57710 69514
rect 57854 69438 57870 69722
rect 71284 69498 71350 70178
rect 71948 70178 71968 70310
rect 72002 70266 72014 70350
rect 72612 72954 72626 73106
rect 72660 73074 72670 73126
rect 73284 73126 73318 73142
rect 72660 72954 72668 73074
rect 72612 72432 72668 72954
rect 72612 72260 72626 72432
rect 72660 72260 72668 72432
rect 72612 71738 72668 72260
rect 72612 71566 72626 71738
rect 72660 71566 72668 71738
rect 72612 71044 72668 71566
rect 72612 70872 72626 71044
rect 72660 70872 72668 71044
rect 72612 70350 72668 70872
rect 72002 70178 72008 70266
rect 72612 70262 72626 70350
rect 71948 70068 72008 70178
rect 72660 70262 72668 70350
rect 73272 72954 73284 73064
rect 73924 73126 74000 73222
rect 75156 73212 77974 73254
rect 79006 73226 81824 73268
rect 73318 72954 73328 73064
rect 73924 73044 73942 73126
rect 73272 72432 73328 72954
rect 73272 72260 73284 72432
rect 73318 72260 73328 72432
rect 73272 71738 73328 72260
rect 73272 71566 73284 71738
rect 73318 71566 73328 71738
rect 73272 71044 73328 71566
rect 73272 70872 73284 71044
rect 73318 70872 73328 71044
rect 73272 70350 73328 70872
rect 73272 70220 73284 70350
rect 72626 70162 72660 70178
rect 73276 70178 73284 70220
rect 73318 70308 73328 70350
rect 73926 72954 73942 73044
rect 73976 73044 74000 73126
rect 75160 73106 75216 73212
rect 74876 73046 75092 73106
rect 73976 72954 73982 73044
rect 73926 72432 73982 72954
rect 73926 72260 73942 72432
rect 73976 72260 73982 72432
rect 73926 71738 73982 72260
rect 73926 71566 73942 71738
rect 73976 71566 73982 71738
rect 73926 71044 73982 71566
rect 73926 70872 73942 71044
rect 73976 70872 73982 71044
rect 73926 70350 73982 70872
rect 73318 70178 73336 70308
rect 73926 70224 73942 70350
rect 73276 70072 73336 70178
rect 73976 70224 73982 70350
rect 74876 70300 74906 73046
rect 75046 70300 75092 73046
rect 74876 70246 75092 70300
rect 75160 72934 75174 73106
rect 75208 72934 75216 73106
rect 75832 73106 75866 73122
rect 75160 72412 75216 72934
rect 75160 72240 75174 72412
rect 75208 72240 75216 72412
rect 75160 71718 75216 72240
rect 75160 71546 75174 71718
rect 75208 71546 75216 71718
rect 75160 71024 75216 71546
rect 75160 70852 75174 71024
rect 75208 70852 75216 71024
rect 75160 70330 75216 70852
rect 75160 70282 75174 70330
rect 73942 70162 73976 70178
rect 75148 70158 75174 70282
rect 75208 70258 75216 70330
rect 75822 72934 75832 73090
rect 76478 73106 76534 73212
rect 77788 73202 77974 73212
rect 75866 72934 75878 73090
rect 76478 73086 76490 73106
rect 75822 72412 75878 72934
rect 75822 72240 75832 72412
rect 75866 72240 75878 72412
rect 75822 71718 75878 72240
rect 75822 71546 75832 71718
rect 75866 71546 75878 71718
rect 75822 71024 75878 71546
rect 75822 70852 75832 71024
rect 75866 70852 75878 71024
rect 75822 70330 75878 70852
rect 75822 70290 75832 70330
rect 75208 70158 75214 70258
rect 73276 70068 73434 70072
rect 71948 70006 73434 70068
rect 71948 70000 72008 70006
rect 73258 70002 73336 70006
rect 73276 69998 73336 70002
rect 73928 69506 74106 69516
rect 73920 69498 74106 69506
rect 71284 69456 74106 69498
rect 71284 69440 71350 69456
rect 57692 69408 57870 69438
rect 71292 69350 71348 69440
rect 45278 69042 45542 69060
rect 49272 69042 49536 69060
rect 53294 69042 53558 69060
rect 57316 69042 57584 69060
rect 42476 69030 57584 69042
rect 42386 68996 42402 69030
rect 42574 68996 43096 69030
rect 43268 68996 43790 69030
rect 43962 68996 44484 69030
rect 44656 68996 45178 69030
rect 45350 68996 46396 69030
rect 46568 68996 47090 69030
rect 47262 68996 47784 69030
rect 47956 68996 48478 69030
rect 48650 68996 49172 69030
rect 49344 68996 50418 69030
rect 50590 68996 51112 69030
rect 51284 68996 51806 69030
rect 51978 68996 52500 69030
rect 52672 68996 53194 69030
rect 53366 68996 54440 69030
rect 54612 68996 55134 69030
rect 55306 68996 55828 69030
rect 56000 68996 56522 69030
rect 56694 68996 57216 69030
rect 57388 68996 57584 69030
rect 42476 68992 57584 68996
rect 71008 69290 71224 69350
rect 42476 68990 57580 68992
rect 42476 68988 45542 68990
rect 46470 68988 49536 68990
rect 50492 68988 53558 68990
rect 54514 68988 57580 68990
rect 45278 68984 45542 68988
rect 49272 68984 49536 68988
rect 53294 68984 53558 68988
rect 57316 68984 57580 68988
rect 42214 68384 42510 68398
rect 42214 68372 45360 68384
rect 42214 68338 42402 68372
rect 42574 68338 43096 68372
rect 43268 68338 43790 68372
rect 43962 68338 44484 68372
rect 44656 68338 45178 68372
rect 45350 68338 45366 68372
rect 42214 68330 45360 68338
rect 42214 68322 42510 68330
rect 42214 68222 42306 68322
rect 42224 67076 42306 68222
rect 45464 67732 45518 68984
rect 46218 68384 46504 68398
rect 46218 68372 49354 68384
rect 46218 68338 46396 68372
rect 46568 68338 47090 68372
rect 47262 68338 47784 68372
rect 47956 68338 48478 68372
rect 48650 68338 49172 68372
rect 49344 68338 49360 68372
rect 46218 68330 49354 68338
rect 46218 68322 46504 68330
rect 45314 67726 45578 67732
rect 42524 67714 45578 67726
rect 42386 67680 42402 67714
rect 42574 67680 43096 67714
rect 43268 67680 43790 67714
rect 43962 67680 44484 67714
rect 44656 67680 45178 67714
rect 45350 67680 45578 67714
rect 42524 67672 45578 67680
rect 45314 67656 45578 67672
rect 42220 67068 42540 67076
rect 42220 67056 45368 67068
rect 42220 67022 42402 67056
rect 42574 67022 43096 67056
rect 43268 67022 43790 67056
rect 43962 67022 44484 67056
rect 44656 67022 45178 67056
rect 45350 67022 45368 67056
rect 42220 67014 45368 67022
rect 42220 67000 42540 67014
rect 19392 65970 20628 65994
rect 972 65928 2604 65962
rect 972 65786 1028 65928
rect 2542 65786 2604 65928
rect 972 65758 2604 65786
rect 3640 65924 5272 65958
rect 3640 65782 3696 65924
rect 5210 65782 5272 65924
rect 3640 65754 5272 65782
rect 6314 65930 7946 65964
rect 6314 65788 6370 65930
rect 7884 65788 7946 65930
rect 6314 65760 7946 65788
rect 8960 65930 10592 65964
rect 8960 65788 9016 65930
rect 10530 65788 10592 65930
rect 8960 65760 10592 65788
rect 11614 65924 13246 65958
rect 11614 65782 11670 65924
rect 13184 65782 13246 65924
rect 11614 65754 13246 65782
rect 14268 65930 15900 65964
rect 14268 65788 14324 65930
rect 15838 65788 15900 65930
rect 14268 65760 15900 65788
rect 16894 65934 18526 65968
rect 16894 65792 16950 65934
rect 18464 65792 18526 65934
rect 16894 65764 18526 65792
rect 19392 65776 19500 65970
rect 20566 65776 20628 65970
rect 19392 65724 20628 65776
rect 42224 65770 42306 67000
rect 45464 66418 45518 67656
rect 46218 67076 46300 68322
rect 49458 67732 49512 68984
rect 50240 68384 50526 68398
rect 50240 68372 53376 68384
rect 50240 68338 50418 68372
rect 50590 68338 51112 68372
rect 51284 68338 51806 68372
rect 51978 68338 52500 68372
rect 52672 68338 53194 68372
rect 53366 68338 53382 68372
rect 50240 68330 53376 68338
rect 50240 68322 50526 68330
rect 49308 67726 49572 67732
rect 46518 67714 49572 67726
rect 46380 67680 46396 67714
rect 46568 67680 47090 67714
rect 47262 67680 47784 67714
rect 47956 67680 48478 67714
rect 48650 67680 49172 67714
rect 49344 67680 49572 67714
rect 46518 67672 49572 67680
rect 49308 67656 49572 67672
rect 46214 67068 46534 67076
rect 46214 67056 49362 67068
rect 46214 67022 46396 67056
rect 46568 67022 47090 67056
rect 47262 67022 47784 67056
rect 47956 67022 48478 67056
rect 48650 67022 49172 67056
rect 49344 67022 49362 67056
rect 46214 67014 49362 67022
rect 46214 67000 46534 67014
rect 45284 66404 45548 66418
rect 42522 66398 45548 66404
rect 42386 66364 42402 66398
rect 42574 66364 43096 66398
rect 43268 66364 43790 66398
rect 43962 66364 44484 66398
rect 44656 66364 45178 66398
rect 45350 66364 45548 66398
rect 42522 66350 45548 66364
rect 45284 66342 45548 66350
rect 45464 66340 45518 66342
rect 46218 65770 46300 67000
rect 49458 66418 49512 67656
rect 50240 67076 50322 68322
rect 53480 67732 53534 68984
rect 57462 68842 57556 68984
rect 54262 68384 54548 68398
rect 54262 68372 57398 68384
rect 54262 68338 54440 68372
rect 54612 68338 55134 68372
rect 55306 68338 55828 68372
rect 56000 68338 56522 68372
rect 56694 68338 57216 68372
rect 57388 68338 57404 68372
rect 54262 68330 57398 68338
rect 54262 68322 54548 68330
rect 53330 67726 53594 67732
rect 50540 67714 53594 67726
rect 50402 67680 50418 67714
rect 50590 67680 51112 67714
rect 51284 67680 51806 67714
rect 51978 67680 52500 67714
rect 52672 67680 53194 67714
rect 53366 67680 53594 67714
rect 50540 67672 53594 67680
rect 53330 67656 53594 67672
rect 50236 67068 50556 67076
rect 50236 67056 53384 67068
rect 50236 67022 50418 67056
rect 50590 67022 51112 67056
rect 51284 67022 51806 67056
rect 51978 67022 52500 67056
rect 52672 67022 53194 67056
rect 53366 67022 53384 67056
rect 50236 67014 53384 67022
rect 50236 67000 50556 67014
rect 49278 66404 49542 66418
rect 46516 66398 49542 66404
rect 46380 66364 46396 66398
rect 46568 66364 47090 66398
rect 47262 66364 47784 66398
rect 47956 66364 48478 66398
rect 48650 66364 49172 66398
rect 49344 66364 49542 66398
rect 46516 66350 49542 66364
rect 49278 66342 49542 66350
rect 49458 66340 49512 66342
rect 50240 65770 50322 67000
rect 53480 66418 53534 67656
rect 54262 67076 54344 68322
rect 57502 67732 57556 68842
rect 57352 67726 57616 67732
rect 54562 67714 57616 67726
rect 54424 67680 54440 67714
rect 54612 67680 55134 67714
rect 55306 67680 55828 67714
rect 56000 67680 56522 67714
rect 56694 67680 57216 67714
rect 57388 67680 57616 67714
rect 54562 67672 57616 67680
rect 57352 67656 57616 67672
rect 54258 67068 54578 67076
rect 54258 67056 57406 67068
rect 54258 67022 54440 67056
rect 54612 67022 55134 67056
rect 55306 67022 55828 67056
rect 56000 67022 56522 67056
rect 56694 67022 57216 67056
rect 57388 67022 57406 67056
rect 54258 67014 57406 67022
rect 54258 67000 54578 67014
rect 53300 66404 53564 66418
rect 50538 66398 53564 66404
rect 50402 66364 50418 66398
rect 50590 66364 51112 66398
rect 51284 66364 51806 66398
rect 51978 66364 52500 66398
rect 52672 66364 53194 66398
rect 53366 66364 53564 66398
rect 50538 66350 53564 66364
rect 53300 66342 53564 66350
rect 53480 66340 53534 66342
rect 54262 65770 54344 67000
rect 57502 66418 57556 67656
rect 71008 66544 71038 69290
rect 71178 66544 71224 69290
rect 71292 69178 71306 69350
rect 71340 69178 71348 69350
rect 71964 69350 71998 69366
rect 71292 68656 71348 69178
rect 71292 68484 71306 68656
rect 71340 68484 71348 68656
rect 71292 67962 71348 68484
rect 71292 67790 71306 67962
rect 71340 67790 71348 67962
rect 71292 67268 71348 67790
rect 71292 67096 71306 67268
rect 71340 67096 71348 67268
rect 71292 66574 71348 67096
rect 71292 66562 71306 66574
rect 71008 66490 71224 66544
rect 57322 66408 57586 66418
rect 57322 66404 57604 66408
rect 54560 66398 57604 66404
rect 54424 66364 54440 66398
rect 54612 66364 55134 66398
rect 55306 66364 55828 66398
rect 56000 66364 56522 66398
rect 56694 66364 57216 66398
rect 57388 66364 57604 66398
rect 54560 66350 57604 66364
rect 57322 66342 57604 66350
rect 42220 65758 42520 65770
rect 46214 65758 46514 65770
rect 50236 65758 50536 65770
rect 54258 65758 54558 65770
rect 57450 65766 57604 66342
rect 71276 66402 71306 66562
rect 71340 66562 71348 66574
rect 71954 69178 71964 69334
rect 72610 69350 72666 69456
rect 73920 69446 74106 69456
rect 75148 69478 75214 70158
rect 75812 70158 75832 70290
rect 75866 70246 75878 70330
rect 76476 72934 76490 73086
rect 76524 73054 76534 73106
rect 77148 73106 77182 73122
rect 76524 72934 76532 73054
rect 76476 72412 76532 72934
rect 76476 72240 76490 72412
rect 76524 72240 76532 72412
rect 76476 71718 76532 72240
rect 76476 71546 76490 71718
rect 76524 71546 76532 71718
rect 76476 71024 76532 71546
rect 76476 70852 76490 71024
rect 76524 70852 76532 71024
rect 76476 70330 76532 70852
rect 75866 70158 75872 70246
rect 76476 70242 76490 70330
rect 75812 70048 75872 70158
rect 76524 70242 76532 70330
rect 77136 72934 77148 73044
rect 77788 73106 77864 73202
rect 79010 73120 79066 73226
rect 77182 72934 77192 73044
rect 77788 73024 77806 73106
rect 77136 72412 77192 72934
rect 77136 72240 77148 72412
rect 77182 72240 77192 72412
rect 77136 71718 77192 72240
rect 77136 71546 77148 71718
rect 77182 71546 77192 71718
rect 77136 71024 77192 71546
rect 77136 70852 77148 71024
rect 77182 70852 77192 71024
rect 77136 70330 77192 70852
rect 77136 70200 77148 70330
rect 76490 70142 76524 70158
rect 77140 70158 77148 70200
rect 77182 70288 77192 70330
rect 77790 72934 77806 73024
rect 77840 73024 77864 73106
rect 78726 73060 78942 73120
rect 77840 72934 77846 73024
rect 77790 72412 77846 72934
rect 77790 72240 77806 72412
rect 77840 72240 77846 72412
rect 77790 71718 77846 72240
rect 77790 71546 77806 71718
rect 77840 71546 77846 71718
rect 77790 71024 77846 71546
rect 77790 70852 77806 71024
rect 77840 70852 77846 71024
rect 77790 70330 77846 70852
rect 77182 70158 77200 70288
rect 77790 70204 77806 70330
rect 77140 70052 77200 70158
rect 77840 70204 77846 70330
rect 78726 70314 78756 73060
rect 78896 72856 78942 73060
rect 79010 72948 79024 73120
rect 79058 72948 79066 73120
rect 79682 73120 79716 73136
rect 79010 72856 79066 72948
rect 78896 72780 79066 72856
rect 78896 70314 78942 72780
rect 78726 70260 78942 70314
rect 79010 72426 79066 72780
rect 79010 72254 79024 72426
rect 79058 72254 79066 72426
rect 79010 71732 79066 72254
rect 79010 71560 79024 71732
rect 79058 71560 79066 71732
rect 79010 71038 79066 71560
rect 79010 70866 79024 71038
rect 79058 70866 79066 71038
rect 79010 70344 79066 70866
rect 79010 70296 79024 70344
rect 77806 70142 77840 70158
rect 78998 70172 79024 70296
rect 79058 70272 79066 70344
rect 79672 72948 79682 73104
rect 80328 73120 80384 73226
rect 81638 73216 81824 73226
rect 79716 72948 79728 73104
rect 80328 73100 80340 73120
rect 79672 72426 79728 72948
rect 79672 72254 79682 72426
rect 79716 72254 79728 72426
rect 79672 71732 79728 72254
rect 79672 71560 79682 71732
rect 79716 71560 79728 71732
rect 79672 71038 79728 71560
rect 79672 70866 79682 71038
rect 79716 70866 79728 71038
rect 79672 70344 79728 70866
rect 79672 70304 79682 70344
rect 79058 70172 79064 70272
rect 77140 70048 77298 70052
rect 75812 69986 77298 70048
rect 75812 69980 75872 69986
rect 77122 69982 77200 69986
rect 77140 69978 77200 69982
rect 77792 69486 77970 69496
rect 77784 69478 77970 69486
rect 71998 69178 72010 69334
rect 72610 69330 72622 69350
rect 71954 68656 72010 69178
rect 71954 68484 71964 68656
rect 71998 68484 72010 68656
rect 71954 67962 72010 68484
rect 71954 67790 71964 67962
rect 71998 67790 72010 67962
rect 71954 67268 72010 67790
rect 71954 67096 71964 67268
rect 71998 67096 72010 67268
rect 71954 66574 72010 67096
rect 71340 66402 71358 66562
rect 71954 66534 71964 66574
rect 57160 65758 57656 65766
rect 42220 65740 57656 65758
rect 20400 65682 20522 65724
rect 42220 65706 42402 65740
rect 42574 65706 43096 65740
rect 43268 65706 43790 65740
rect 43962 65706 44484 65740
rect 44656 65706 45178 65740
rect 45350 65706 46396 65740
rect 46568 65706 47090 65740
rect 47262 65706 47784 65740
rect 47956 65706 48478 65740
rect 48650 65706 49172 65740
rect 49344 65706 50418 65740
rect 50590 65706 51112 65740
rect 51284 65706 51806 65740
rect 51978 65706 52500 65740
rect 52672 65706 53194 65740
rect 53366 65706 54440 65740
rect 54612 65706 55134 65740
rect 55306 65706 55828 65740
rect 56000 65706 56522 65740
rect 56694 65706 57216 65740
rect 57388 65706 57656 65740
rect 42220 65696 45362 65706
rect 46214 65696 49356 65706
rect 50236 65696 53378 65706
rect 54258 65696 57656 65706
rect 71276 65728 71358 66402
rect 71944 66402 71964 66534
rect 71998 66490 72010 66574
rect 72608 69178 72622 69330
rect 72656 69298 72666 69350
rect 73280 69350 73314 69366
rect 72656 69178 72664 69298
rect 72608 68656 72664 69178
rect 72608 68484 72622 68656
rect 72656 68484 72664 68656
rect 72608 67962 72664 68484
rect 72608 67790 72622 67962
rect 72656 67790 72664 67962
rect 72608 67268 72664 67790
rect 72608 67096 72622 67268
rect 72656 67096 72664 67268
rect 72608 66574 72664 67096
rect 71998 66402 72004 66490
rect 72608 66486 72622 66574
rect 71944 66292 72004 66402
rect 72656 66486 72664 66574
rect 73268 69178 73280 69288
rect 73920 69350 73996 69446
rect 75148 69436 77970 69478
rect 75148 69420 75214 69436
rect 73314 69178 73324 69288
rect 73920 69268 73938 69350
rect 73268 68656 73324 69178
rect 73268 68484 73280 68656
rect 73314 68484 73324 68656
rect 73268 67962 73324 68484
rect 73268 67790 73280 67962
rect 73314 67790 73324 67962
rect 73268 67268 73324 67790
rect 73268 67096 73280 67268
rect 73314 67096 73324 67268
rect 73268 66574 73324 67096
rect 73268 66444 73280 66574
rect 72622 66386 72656 66402
rect 73272 66402 73280 66444
rect 73314 66532 73324 66574
rect 73922 69178 73938 69268
rect 73972 69268 73996 69350
rect 75156 69330 75212 69420
rect 74872 69270 75088 69330
rect 73972 69178 73978 69268
rect 73922 68656 73978 69178
rect 73922 68484 73938 68656
rect 73972 68484 73978 68656
rect 73922 67962 73978 68484
rect 73922 67790 73938 67962
rect 73972 67790 73978 67962
rect 73922 67268 73978 67790
rect 73922 67096 73938 67268
rect 73972 67096 73978 67268
rect 73922 66574 73978 67096
rect 73314 66402 73332 66532
rect 73922 66448 73938 66574
rect 73272 66296 73332 66402
rect 73972 66448 73978 66574
rect 74872 66524 74902 69270
rect 75042 66524 75088 69270
rect 75156 69158 75170 69330
rect 75204 69158 75212 69330
rect 75828 69330 75862 69346
rect 75156 68636 75212 69158
rect 75156 68464 75170 68636
rect 75204 68464 75212 68636
rect 75156 67942 75212 68464
rect 75156 67770 75170 67942
rect 75204 67770 75212 67942
rect 75156 67248 75212 67770
rect 75156 67076 75170 67248
rect 75204 67076 75212 67248
rect 75156 66554 75212 67076
rect 75156 66542 75170 66554
rect 74872 66470 75088 66524
rect 73938 66386 73972 66402
rect 75140 66382 75170 66542
rect 75204 66542 75212 66554
rect 75818 69158 75828 69314
rect 76474 69330 76530 69436
rect 77784 69426 77970 69436
rect 78998 69492 79064 70172
rect 79662 70172 79682 70304
rect 79716 70260 79728 70344
rect 80326 72948 80340 73100
rect 80374 73068 80384 73120
rect 80998 73120 81032 73136
rect 80374 72948 80382 73068
rect 80326 72426 80382 72948
rect 80326 72254 80340 72426
rect 80374 72254 80382 72426
rect 80326 71732 80382 72254
rect 80326 71560 80340 71732
rect 80374 71560 80382 71732
rect 80326 71038 80382 71560
rect 80326 70866 80340 71038
rect 80374 70866 80382 71038
rect 80326 70344 80382 70866
rect 79716 70172 79722 70260
rect 80326 70256 80340 70344
rect 79662 70062 79722 70172
rect 80374 70256 80382 70344
rect 80986 72948 80998 73058
rect 81638 73120 81714 73216
rect 81032 72948 81042 73058
rect 81638 73038 81656 73120
rect 80986 72426 81042 72948
rect 80986 72254 80998 72426
rect 81032 72254 81042 72426
rect 80986 71732 81042 72254
rect 80986 71560 80998 71732
rect 81032 71560 81042 71732
rect 80986 71038 81042 71560
rect 80986 70866 80998 71038
rect 81032 70866 81042 71038
rect 80986 70344 81042 70866
rect 80986 70214 80998 70344
rect 80340 70156 80374 70172
rect 80990 70172 80998 70214
rect 81032 70302 81042 70344
rect 81640 72948 81656 73038
rect 81690 73038 81714 73120
rect 81690 72948 81696 73038
rect 81640 72426 81696 72948
rect 81640 72254 81656 72426
rect 81690 72254 81696 72426
rect 81640 71732 81696 72254
rect 81640 71560 81656 71732
rect 81690 71560 81696 71732
rect 81640 71038 81696 71560
rect 81640 70866 81656 71038
rect 81690 70866 81696 71038
rect 81640 70344 81696 70866
rect 81032 70172 81050 70302
rect 81640 70218 81656 70344
rect 80990 70066 81050 70172
rect 81690 70218 81696 70344
rect 81656 70156 81690 70172
rect 80990 70062 81148 70066
rect 79662 70000 81148 70062
rect 79662 69994 79722 70000
rect 80972 69996 81050 70000
rect 80990 69992 81050 69996
rect 81642 69500 81820 69510
rect 81634 69492 81820 69500
rect 78998 69450 81820 69492
rect 78998 69434 79064 69450
rect 75862 69158 75874 69314
rect 76474 69310 76486 69330
rect 75818 68636 75874 69158
rect 75818 68464 75828 68636
rect 75862 68464 75874 68636
rect 75818 67942 75874 68464
rect 75818 67770 75828 67942
rect 75862 67770 75874 67942
rect 75818 67248 75874 67770
rect 75818 67076 75828 67248
rect 75862 67076 75874 67248
rect 75818 66554 75874 67076
rect 75204 66382 75222 66542
rect 75818 66514 75828 66554
rect 73272 66292 73430 66296
rect 71944 66230 73430 66292
rect 71944 66224 72004 66230
rect 73272 66222 73332 66230
rect 73928 65736 74106 65746
rect 73920 65728 74106 65736
rect 71276 65696 74106 65728
rect 42220 65694 42502 65696
rect 46214 65694 46496 65696
rect 50236 65694 50518 65696
rect 54258 65694 54540 65696
rect 42224 65692 42306 65694
rect 46218 65692 46300 65694
rect 50240 65692 50322 65694
rect 54262 65692 54344 65694
rect 2388 65640 20556 65682
rect 57160 65642 57656 65696
rect 71288 65686 74106 65696
rect 2388 65632 20580 65640
rect 2388 65620 20588 65632
rect 2388 65588 19572 65620
rect 936 65586 19572 65588
rect 19744 65586 20266 65620
rect 20438 65586 20588 65620
rect 936 65576 20588 65586
rect 936 65572 16888 65576
rect 936 65570 6308 65572
rect 936 65536 966 65570
rect 1138 65536 1660 65570
rect 1832 65536 2354 65570
rect 2526 65566 6308 65570
rect 2526 65536 3634 65566
rect 936 65532 3634 65536
rect 3806 65532 4328 65566
rect 4500 65532 5022 65566
rect 5194 65538 6308 65566
rect 6480 65538 7002 65572
rect 7174 65538 7696 65572
rect 7868 65538 8954 65572
rect 9126 65538 9648 65572
rect 9820 65538 10342 65572
rect 10514 65566 14262 65572
rect 10514 65538 11608 65566
rect 5194 65532 11608 65538
rect 11780 65532 12302 65566
rect 12474 65532 12996 65566
rect 13168 65538 14262 65566
rect 14434 65538 14956 65572
rect 15128 65538 15650 65572
rect 15822 65542 16888 65572
rect 17060 65542 17582 65576
rect 17754 65542 18276 65576
rect 18448 65542 20588 65576
rect 15822 65538 20588 65542
rect 13168 65532 20588 65538
rect 936 65524 20588 65532
rect 2388 65512 20588 65524
rect 774 64924 1094 64946
rect 774 64922 2502 64924
rect 756 64912 2502 64922
rect 756 64878 966 64912
rect 1138 64878 1660 64912
rect 1832 64878 2354 64912
rect 2526 64878 2542 64912
rect 756 64872 2502 64878
rect 756 64824 1094 64872
rect 756 63624 848 64824
rect 2638 64262 2706 65512
rect 3442 64920 3762 64942
rect 3442 64918 5170 64920
rect 984 64254 2706 64262
rect 950 64220 966 64254
rect 1138 64220 1660 64254
rect 1832 64220 2354 64254
rect 2526 64220 2706 64254
rect 984 64210 2706 64220
rect 2418 64208 2706 64210
rect 756 63602 1080 63624
rect 756 63596 2506 63602
rect 756 63562 966 63596
rect 1138 63562 1660 63596
rect 1832 63562 2354 63596
rect 2526 63562 2542 63596
rect 756 63550 2506 63562
rect 756 63502 1080 63550
rect 756 62310 848 63502
rect 2638 62950 2706 64208
rect 2430 62948 2706 62950
rect 998 62938 2706 62948
rect 950 62904 966 62938
rect 1138 62904 1660 62938
rect 1832 62904 2354 62938
rect 2526 62904 2706 62938
rect 998 62896 2706 62904
rect 750 62288 1070 62310
rect 750 62280 2516 62288
rect 750 62246 966 62280
rect 1138 62246 1660 62280
rect 1832 62246 2354 62280
rect 2526 62246 2542 62280
rect 750 62236 2516 62246
rect 750 62188 1070 62236
rect 756 61022 848 62188
rect 2638 61632 2706 62896
rect 3424 64908 5170 64918
rect 3424 64874 3634 64908
rect 3806 64874 4328 64908
rect 4500 64874 5022 64908
rect 5194 64874 5210 64908
rect 3424 64868 5170 64874
rect 3424 64820 3762 64868
rect 3424 63620 3516 64820
rect 5306 64258 5374 65512
rect 6116 64926 6436 64948
rect 6116 64924 7844 64926
rect 3652 64250 5374 64258
rect 3618 64216 3634 64250
rect 3806 64216 4328 64250
rect 4500 64216 5022 64250
rect 5194 64216 5374 64250
rect 3652 64206 5374 64216
rect 5086 64204 5374 64206
rect 3424 63598 3748 63620
rect 3424 63592 5174 63598
rect 3424 63558 3634 63592
rect 3806 63558 4328 63592
rect 4500 63558 5022 63592
rect 5194 63558 5210 63592
rect 3424 63546 5174 63558
rect 3424 63498 3748 63546
rect 3424 62306 3516 63498
rect 5306 62946 5374 64204
rect 5098 62944 5374 62946
rect 3666 62934 5374 62944
rect 3618 62900 3634 62934
rect 3806 62900 4328 62934
rect 4500 62900 5022 62934
rect 5194 62900 5374 62934
rect 3666 62892 5374 62900
rect 3418 62284 3738 62306
rect 3418 62276 5184 62284
rect 3418 62242 3634 62276
rect 3806 62242 4328 62276
rect 4500 62242 5022 62276
rect 5194 62242 5210 62276
rect 3418 62232 5184 62242
rect 3418 62184 3738 62232
rect 2420 61630 2706 61632
rect 1022 61622 2706 61630
rect 950 61588 966 61622
rect 1138 61588 1660 61622
rect 1832 61588 2354 61622
rect 2526 61588 2706 61622
rect 1022 61578 2706 61588
rect 740 60974 1060 61022
rect 740 60964 2564 60974
rect 740 60930 966 60964
rect 1138 60930 1660 60964
rect 1832 60930 2354 60964
rect 2526 60930 2564 60964
rect 2638 60946 2706 61578
rect 740 60922 2564 60930
rect 740 60900 1060 60922
rect 2628 60904 2706 60946
rect 2628 60320 2702 60904
rect 3424 61018 3516 62184
rect 5306 61628 5374 62892
rect 6098 64914 7844 64924
rect 6098 64880 6308 64914
rect 6480 64880 7002 64914
rect 7174 64880 7696 64914
rect 7868 64880 7884 64914
rect 6098 64874 7844 64880
rect 6098 64826 6436 64874
rect 6098 63626 6190 64826
rect 7980 64264 8048 65512
rect 8762 64926 9082 64948
rect 8762 64924 10490 64926
rect 6326 64256 8048 64264
rect 6292 64222 6308 64256
rect 6480 64222 7002 64256
rect 7174 64222 7696 64256
rect 7868 64222 8048 64256
rect 6326 64212 8048 64222
rect 7760 64210 8048 64212
rect 6098 63604 6422 63626
rect 6098 63598 7848 63604
rect 6098 63564 6308 63598
rect 6480 63564 7002 63598
rect 7174 63564 7696 63598
rect 7868 63564 7884 63598
rect 6098 63552 7848 63564
rect 6098 63504 6422 63552
rect 6098 62312 6190 63504
rect 7980 62952 8048 64210
rect 7772 62950 8048 62952
rect 6340 62940 8048 62950
rect 6292 62906 6308 62940
rect 6480 62906 7002 62940
rect 7174 62906 7696 62940
rect 7868 62906 8048 62940
rect 6340 62898 8048 62906
rect 6092 62290 6412 62312
rect 6092 62282 7858 62290
rect 6092 62248 6308 62282
rect 6480 62248 7002 62282
rect 7174 62248 7696 62282
rect 7868 62248 7884 62282
rect 6092 62238 7858 62248
rect 6092 62190 6412 62238
rect 5088 61626 5374 61628
rect 3690 61618 5374 61626
rect 3618 61584 3634 61618
rect 3806 61584 4328 61618
rect 4500 61584 5022 61618
rect 5194 61584 5374 61618
rect 3690 61574 5374 61584
rect 3408 61010 3728 61018
rect 3304 60970 3728 61010
rect 3304 60960 5232 60970
rect 3304 60926 3634 60960
rect 3806 60926 4328 60960
rect 4500 60926 5022 60960
rect 5194 60926 5232 60960
rect 5306 60942 5374 61574
rect 3304 60918 5232 60926
rect 3304 60896 3728 60918
rect 5296 60900 5374 60942
rect 3304 60868 3532 60896
rect 2484 60314 2706 60320
rect 5296 60316 5370 60900
rect 6098 61024 6190 62190
rect 7980 61634 8048 62898
rect 8744 64914 10490 64924
rect 8744 64880 8954 64914
rect 9126 64880 9648 64914
rect 9820 64880 10342 64914
rect 10514 64880 10530 64914
rect 8744 64874 10490 64880
rect 8744 64826 9082 64874
rect 8744 63626 8836 64826
rect 10626 64264 10694 65512
rect 11416 64920 11736 64942
rect 11416 64918 13144 64920
rect 8972 64256 10694 64264
rect 8938 64222 8954 64256
rect 9126 64222 9648 64256
rect 9820 64222 10342 64256
rect 10514 64222 10694 64256
rect 8972 64212 10694 64222
rect 10406 64210 10694 64212
rect 8744 63604 9068 63626
rect 8744 63598 10494 63604
rect 8744 63564 8954 63598
rect 9126 63564 9648 63598
rect 9820 63564 10342 63598
rect 10514 63564 10530 63598
rect 8744 63552 10494 63564
rect 8744 63504 9068 63552
rect 8744 62312 8836 63504
rect 10626 62952 10694 64210
rect 10418 62950 10694 62952
rect 8986 62940 10694 62950
rect 8938 62906 8954 62940
rect 9126 62906 9648 62940
rect 9820 62906 10342 62940
rect 10514 62906 10694 62940
rect 8986 62898 10694 62906
rect 8738 62290 9058 62312
rect 8738 62282 10504 62290
rect 8738 62248 8954 62282
rect 9126 62248 9648 62282
rect 9820 62248 10342 62282
rect 10514 62248 10530 62282
rect 8738 62238 10504 62248
rect 8738 62190 9058 62238
rect 7762 61632 8048 61634
rect 6364 61624 8048 61632
rect 6292 61590 6308 61624
rect 6480 61590 7002 61624
rect 7174 61590 7696 61624
rect 7868 61590 8048 61624
rect 6364 61580 8048 61590
rect 6082 61020 6402 61024
rect 5956 60976 6402 61020
rect 5956 60966 7906 60976
rect 5956 60932 6308 60966
rect 6480 60932 7002 60966
rect 7174 60932 7696 60966
rect 7868 60932 7906 60966
rect 7980 60948 8048 61580
rect 5956 60924 7906 60932
rect 5956 60910 6402 60924
rect 6082 60902 6402 60910
rect 7970 60906 8048 60948
rect 7970 60322 8044 60906
rect 8744 61036 8836 62190
rect 10626 61634 10694 62898
rect 11398 64908 13144 64918
rect 11398 64874 11608 64908
rect 11780 64874 12302 64908
rect 12474 64874 12996 64908
rect 13168 64874 13184 64908
rect 11398 64868 13144 64874
rect 11398 64820 11736 64868
rect 11398 63620 11490 64820
rect 13280 64258 13348 65512
rect 14070 64926 14390 64948
rect 14070 64924 15798 64926
rect 11626 64250 13348 64258
rect 11592 64216 11608 64250
rect 11780 64216 12302 64250
rect 12474 64216 12996 64250
rect 13168 64216 13348 64250
rect 11626 64206 13348 64216
rect 13060 64204 13348 64206
rect 11398 63598 11722 63620
rect 11398 63592 13148 63598
rect 11398 63558 11608 63592
rect 11780 63558 12302 63592
rect 12474 63558 12996 63592
rect 13168 63558 13184 63592
rect 11398 63546 13148 63558
rect 11398 63498 11722 63546
rect 11398 62306 11490 63498
rect 13280 62946 13348 64204
rect 13072 62944 13348 62946
rect 11640 62934 13348 62944
rect 11592 62900 11608 62934
rect 11780 62900 12302 62934
rect 12474 62900 12996 62934
rect 13168 62900 13348 62934
rect 11640 62892 13348 62900
rect 11392 62284 11712 62306
rect 11392 62276 13158 62284
rect 11392 62242 11608 62276
rect 11780 62242 12302 62276
rect 12474 62242 12996 62276
rect 13168 62242 13184 62276
rect 11392 62232 13158 62242
rect 11392 62184 11712 62232
rect 10408 61632 10694 61634
rect 9010 61624 10694 61632
rect 8938 61590 8954 61624
rect 9126 61590 9648 61624
rect 9820 61590 10342 61624
rect 10514 61590 10694 61624
rect 9010 61580 10694 61590
rect 8582 61024 8850 61036
rect 8582 60976 9048 61024
rect 8582 60966 10552 60976
rect 8582 60932 8954 60966
rect 9126 60932 9648 60966
rect 9820 60932 10342 60966
rect 10514 60932 10552 60966
rect 10626 60948 10694 61580
rect 8582 60924 10552 60932
rect 8582 60910 9048 60924
rect 8728 60902 9048 60910
rect 10616 60906 10694 60948
rect 10616 60322 10690 60906
rect 11398 61028 11490 62184
rect 13280 61628 13348 62892
rect 14052 64914 15798 64924
rect 14052 64880 14262 64914
rect 14434 64880 14956 64914
rect 15128 64880 15650 64914
rect 15822 64880 15838 64914
rect 14052 64874 15798 64880
rect 14052 64826 14390 64874
rect 14052 63626 14144 64826
rect 15934 64264 16002 65512
rect 16696 64930 17016 64952
rect 16696 64928 18424 64930
rect 14280 64256 16002 64264
rect 14246 64222 14262 64256
rect 14434 64222 14956 64256
rect 15128 64222 15650 64256
rect 15822 64222 16002 64256
rect 14280 64212 16002 64222
rect 15714 64210 16002 64212
rect 14052 63604 14376 63626
rect 14052 63598 15802 63604
rect 14052 63564 14262 63598
rect 14434 63564 14956 63598
rect 15128 63564 15650 63598
rect 15822 63564 15838 63598
rect 14052 63552 15802 63564
rect 14052 63504 14376 63552
rect 14052 62312 14144 63504
rect 15934 62952 16002 64210
rect 15726 62950 16002 62952
rect 14294 62940 16002 62950
rect 14246 62906 14262 62940
rect 14434 62906 14956 62940
rect 15128 62906 15650 62940
rect 15822 62906 16002 62940
rect 14294 62898 16002 62906
rect 14046 62290 14366 62312
rect 14046 62282 15812 62290
rect 14046 62248 14262 62282
rect 14434 62248 14956 62282
rect 15128 62248 15650 62282
rect 15822 62248 15838 62282
rect 14046 62238 15812 62248
rect 14046 62190 14366 62238
rect 13062 61626 13348 61628
rect 11664 61618 13348 61626
rect 11592 61584 11608 61618
rect 11780 61584 12302 61618
rect 12474 61584 12996 61618
rect 13168 61584 13348 61618
rect 11664 61574 13348 61584
rect 11274 60970 11948 61028
rect 11274 60960 13206 60970
rect 11274 60926 11608 60960
rect 11780 60926 12302 60960
rect 12474 60926 12996 60960
rect 13168 60926 13206 60960
rect 13280 60942 13348 61574
rect 11274 60918 13206 60926
rect 11274 60910 11948 60918
rect 11382 60896 11702 60910
rect 13270 60900 13348 60942
rect 7826 60316 8048 60322
rect 10472 60316 10694 60322
rect 13270 60316 13344 60900
rect 14052 61024 14144 62190
rect 15934 61634 16002 62898
rect 16678 64918 18424 64928
rect 16678 64884 16888 64918
rect 17060 64884 17582 64918
rect 17754 64884 18276 64918
rect 18448 64884 18464 64918
rect 16678 64878 18424 64884
rect 16678 64830 17016 64878
rect 16678 63630 16770 64830
rect 18560 64268 18628 65512
rect 19364 64978 19646 64988
rect 19364 64966 20442 64978
rect 20506 64966 20588 65512
rect 42734 65060 45380 65096
rect 53154 65094 53744 65134
rect 57160 65094 57326 65642
rect 71292 65580 71348 65686
rect 71008 65520 71224 65580
rect 19364 64962 20646 64966
rect 19364 64928 19572 64962
rect 19744 64928 20266 64962
rect 20438 64928 20646 64962
rect 19364 64920 20646 64928
rect 19364 64892 19646 64920
rect 20396 64916 20646 64920
rect 16906 64260 18628 64268
rect 16872 64226 16888 64260
rect 17060 64226 17582 64260
rect 17754 64226 18276 64260
rect 18448 64226 18628 64260
rect 16906 64216 18628 64226
rect 18340 64214 18628 64216
rect 16678 63608 17002 63630
rect 16678 63602 18428 63608
rect 16678 63568 16888 63602
rect 17060 63568 17582 63602
rect 17754 63568 18276 63602
rect 18448 63568 18464 63602
rect 16678 63556 18428 63568
rect 16678 63508 17002 63556
rect 16678 62316 16770 63508
rect 18560 62956 18628 64214
rect 18352 62954 18628 62956
rect 16920 62944 18628 62954
rect 16872 62910 16888 62944
rect 17060 62910 17582 62944
rect 17754 62910 18276 62944
rect 18448 62910 18628 62944
rect 16920 62902 18628 62910
rect 16672 62294 16992 62316
rect 16672 62286 18438 62294
rect 16672 62252 16888 62286
rect 17060 62252 17582 62286
rect 17754 62252 18276 62286
rect 18448 62252 18464 62286
rect 16672 62242 18438 62252
rect 16672 62194 16992 62242
rect 15716 61632 16002 61634
rect 14318 61624 16002 61632
rect 14246 61590 14262 61624
rect 14434 61590 14956 61624
rect 15128 61590 15650 61624
rect 15822 61590 16002 61624
rect 14318 61580 16002 61590
rect 14036 61002 14356 61024
rect 13874 60976 14488 61002
rect 13874 60966 15860 60976
rect 13874 60932 14262 60966
rect 14434 60932 14956 60966
rect 15128 60932 15650 60966
rect 15822 60932 15860 60966
rect 15934 60948 16002 61580
rect 13874 60924 15860 60932
rect 13874 60884 14488 60924
rect 15924 60906 16002 60948
rect 15924 60322 15998 60906
rect 16678 61036 16770 62194
rect 18560 61638 18628 62902
rect 19380 63672 19448 64892
rect 19640 64308 20442 64314
rect 20506 64308 20588 64916
rect 42734 64728 42884 65060
rect 45284 64728 45380 65060
rect 42734 64694 45380 64728
rect 46742 65058 49388 65094
rect 46742 64726 46892 65058
rect 49292 64726 49388 65058
rect 46742 64692 49388 64726
rect 50754 65058 53744 65094
rect 50754 64726 50904 65058
rect 53304 64726 53744 65058
rect 50754 64710 53744 64726
rect 54764 65058 57410 65094
rect 54764 64726 54914 65058
rect 57314 64726 57410 65058
rect 50754 64692 53400 64710
rect 54764 64692 57410 64726
rect 45266 64572 45530 64586
rect 49274 64572 49538 64584
rect 53286 64572 53550 64584
rect 56852 64572 56966 64692
rect 57296 64576 57560 64584
rect 57296 64572 57956 64576
rect 42448 64556 57956 64572
rect 42374 64522 42390 64556
rect 42562 64522 43084 64556
rect 43256 64522 43778 64556
rect 43950 64522 44472 64556
rect 44644 64522 45166 64556
rect 45338 64554 57956 64556
rect 45338 64522 46398 64554
rect 42448 64520 46398 64522
rect 46570 64520 47092 64554
rect 47264 64520 47786 64554
rect 47958 64520 48480 64554
rect 48652 64520 49174 64554
rect 49346 64520 50410 64554
rect 50582 64520 51104 64554
rect 51276 64520 51798 64554
rect 51970 64520 52492 64554
rect 52664 64520 53186 64554
rect 53358 64520 54420 64554
rect 54592 64520 55114 64554
rect 55286 64520 55808 64554
rect 55980 64520 56502 64554
rect 56674 64520 57196 64554
rect 57368 64520 57956 64554
rect 42464 64514 45530 64520
rect 45266 64510 45530 64514
rect 46472 64512 49538 64520
rect 50484 64512 53550 64520
rect 54494 64512 57956 64520
rect 19640 64304 20588 64308
rect 19556 64270 19572 64304
rect 19744 64270 20266 64304
rect 20438 64270 20588 64304
rect 19640 64256 20588 64270
rect 20332 64238 20588 64256
rect 20506 64120 20588 64238
rect 41772 64334 42106 64372
rect 20692 64128 20810 64144
rect 20692 64120 20714 64128
rect 20506 64070 20714 64120
rect 19380 63662 19666 63672
rect 19380 63646 20450 63662
rect 19380 63612 19572 63646
rect 19744 63612 20266 63646
rect 20438 63612 20454 63646
rect 19380 63604 20450 63612
rect 19380 63576 19666 63604
rect 19380 62344 19448 63576
rect 19652 62990 20454 62994
rect 20506 62990 20588 64070
rect 20692 64054 20714 64070
rect 20798 64054 20810 64128
rect 41772 64098 41814 64334
rect 42072 64098 42106 64334
rect 41772 64076 42106 64098
rect 20692 64032 20810 64054
rect 42212 63910 42498 63924
rect 42212 63898 45348 63910
rect 42212 63864 42390 63898
rect 42562 63864 43084 63898
rect 43256 63864 43778 63898
rect 43950 63864 44472 63898
rect 44644 63864 45166 63898
rect 45338 63864 45354 63898
rect 42212 63856 45348 63864
rect 42212 63848 42498 63856
rect 19652 62988 20606 62990
rect 19556 62954 19572 62988
rect 19744 62954 20266 62988
rect 20438 62954 20606 62988
rect 19652 62936 20606 62954
rect 20362 62920 20606 62936
rect 19376 62330 20438 62344
rect 19376 62296 19572 62330
rect 19744 62296 20266 62330
rect 20438 62296 20454 62330
rect 19376 62286 20438 62296
rect 19376 62248 19658 62286
rect 18342 61636 18628 61638
rect 16944 61628 18628 61636
rect 16872 61594 16888 61628
rect 17060 61594 17582 61628
rect 17754 61594 18276 61628
rect 18448 61594 18628 61628
rect 16944 61584 18628 61594
rect 16576 60980 17062 61036
rect 16576 60970 18486 60980
rect 16576 60936 16888 60970
rect 17060 60936 17582 60970
rect 17754 60936 18276 60970
rect 18448 60936 18486 60970
rect 18560 60952 18628 61584
rect 16576 60928 18486 60936
rect 16576 60878 17062 60928
rect 18550 60910 18628 60952
rect 18550 60326 18624 60910
rect 19380 61112 19448 62248
rect 20506 61686 20588 62920
rect 42212 62602 42294 63848
rect 45452 63258 45506 64510
rect 49274 64508 49538 64512
rect 53286 64508 53550 64512
rect 46220 63908 46506 63922
rect 46220 63896 49356 63908
rect 46220 63862 46398 63896
rect 46570 63862 47092 63896
rect 47264 63862 47786 63896
rect 47958 63862 48480 63896
rect 48652 63862 49174 63896
rect 49346 63862 49362 63896
rect 46220 63854 49356 63862
rect 46220 63846 46506 63854
rect 45302 63252 45566 63258
rect 42512 63240 45566 63252
rect 42374 63206 42390 63240
rect 42562 63206 43084 63240
rect 43256 63206 43778 63240
rect 43950 63206 44472 63240
rect 44644 63206 45166 63240
rect 45338 63206 45566 63240
rect 42512 63198 45566 63206
rect 45302 63182 45566 63198
rect 42208 62594 42528 62602
rect 42208 62582 45356 62594
rect 42208 62548 42390 62582
rect 42562 62548 43084 62582
rect 43256 62548 43778 62582
rect 43950 62548 44472 62582
rect 44644 62548 45166 62582
rect 45338 62548 45356 62582
rect 42208 62540 45356 62548
rect 42208 62526 42528 62540
rect 20344 61674 20588 61686
rect 19636 61672 20588 61674
rect 19556 61638 19572 61672
rect 19744 61638 20266 61672
rect 20438 61638 20588 61672
rect 19636 61616 20588 61638
rect 19082 61034 19448 61112
rect 19082 61024 19662 61034
rect 19082 61014 20422 61024
rect 19082 60980 19572 61014
rect 19744 60980 20266 61014
rect 20438 60980 20454 61014
rect 19082 60966 20422 60980
rect 19082 60944 19662 60966
rect 19380 60938 19662 60944
rect 20506 60380 20588 61616
rect 42212 61302 42294 62526
rect 45452 61944 45506 63182
rect 46220 62600 46302 63846
rect 49460 63256 49514 64508
rect 50232 63908 50518 63922
rect 50232 63896 53368 63908
rect 50232 63862 50410 63896
rect 50582 63862 51104 63896
rect 51276 63862 51798 63896
rect 51970 63862 52492 63896
rect 52664 63862 53186 63896
rect 53358 63862 53374 63896
rect 50232 63854 53368 63862
rect 50232 63846 50518 63854
rect 49310 63250 49574 63256
rect 46520 63238 49574 63250
rect 46382 63204 46398 63238
rect 46570 63204 47092 63238
rect 47264 63204 47786 63238
rect 47958 63204 48480 63238
rect 48652 63204 49174 63238
rect 49346 63204 49574 63238
rect 46520 63196 49574 63204
rect 49310 63180 49574 63196
rect 46216 62592 46536 62600
rect 46216 62580 49364 62592
rect 46216 62546 46398 62580
rect 46570 62546 47092 62580
rect 47264 62546 47786 62580
rect 47958 62546 48480 62580
rect 48652 62546 49174 62580
rect 49346 62546 49364 62580
rect 46216 62538 49364 62546
rect 46216 62524 46536 62538
rect 45272 61930 45536 61944
rect 42510 61924 45536 61930
rect 42374 61890 42390 61924
rect 42562 61890 43084 61924
rect 43256 61890 43778 61924
rect 43950 61890 44472 61924
rect 44644 61890 45166 61924
rect 45338 61890 45536 61924
rect 42510 61876 45536 61890
rect 45272 61868 45536 61876
rect 45452 61866 45506 61868
rect 20344 60368 20588 60380
rect 19620 60356 20588 60368
rect 15780 60316 16002 60322
rect 18406 60320 18628 60326
rect 19556 60322 19572 60356
rect 19744 60322 20266 60356
rect 20438 60322 20588 60356
rect 1058 60306 2706 60314
rect 5152 60310 5374 60316
rect 950 60272 966 60306
rect 1138 60272 1660 60306
rect 1832 60272 2354 60306
rect 2526 60272 2706 60306
rect 3726 60302 5374 60310
rect 6400 60308 8048 60316
rect 9046 60308 10694 60316
rect 13126 60310 13348 60316
rect 1058 60262 2706 60272
rect 3618 60268 3634 60302
rect 3806 60268 4328 60302
rect 4500 60268 5022 60302
rect 5194 60268 5374 60302
rect 6292 60274 6308 60308
rect 6480 60274 7002 60308
rect 7174 60274 7696 60308
rect 7868 60274 8048 60308
rect 8938 60274 8954 60308
rect 9126 60274 9648 60308
rect 9820 60274 10342 60308
rect 10514 60274 10694 60308
rect 11700 60302 13348 60310
rect 14354 60308 16002 60316
rect 16980 60312 18628 60320
rect 2484 60250 2706 60262
rect 3726 60258 5374 60268
rect 6400 60264 8048 60274
rect 9046 60264 10694 60274
rect 11592 60268 11608 60302
rect 11780 60268 12302 60302
rect 12474 60268 12996 60302
rect 13168 60268 13348 60302
rect 14246 60274 14262 60308
rect 14434 60274 14956 60308
rect 15128 60274 15650 60308
rect 15822 60274 16002 60308
rect 16872 60278 16888 60312
rect 17060 60278 17582 60312
rect 17754 60278 18276 60312
rect 18448 60278 18628 60312
rect 19620 60310 20588 60322
rect 20506 60304 20588 60310
rect 42194 61296 42294 61302
rect 42194 61286 42508 61296
rect 46220 61294 46302 62524
rect 49460 61942 49514 63180
rect 50232 62600 50314 63846
rect 53472 63256 53526 64508
rect 56852 64504 56966 64512
rect 57296 64508 57956 64512
rect 57408 64420 57956 64508
rect 54242 63908 54528 63922
rect 54242 63896 57378 63908
rect 54242 63862 54420 63896
rect 54592 63862 55114 63896
rect 55286 63862 55808 63896
rect 55980 63862 56502 63896
rect 56674 63862 57196 63896
rect 57368 63862 57384 63896
rect 54242 63854 57378 63862
rect 54242 63846 54528 63854
rect 53322 63250 53586 63256
rect 50532 63238 53586 63250
rect 50394 63204 50410 63238
rect 50582 63204 51104 63238
rect 51276 63204 51798 63238
rect 51970 63204 52492 63238
rect 52664 63204 53186 63238
rect 53358 63204 53586 63238
rect 50532 63196 53586 63204
rect 53322 63180 53586 63196
rect 50228 62592 50548 62600
rect 50228 62580 53376 62592
rect 50228 62546 50410 62580
rect 50582 62546 51104 62580
rect 51276 62546 51798 62580
rect 51970 62546 52492 62580
rect 52664 62546 53186 62580
rect 53358 62546 53376 62580
rect 50228 62538 53376 62546
rect 50228 62524 50548 62538
rect 49280 61928 49544 61942
rect 46518 61922 49544 61928
rect 46382 61888 46398 61922
rect 46570 61888 47092 61922
rect 47264 61888 47786 61922
rect 47958 61888 48480 61922
rect 48652 61888 49174 61922
rect 49346 61888 49544 61922
rect 46518 61874 49544 61888
rect 49280 61866 49544 61874
rect 49460 61864 49514 61866
rect 50232 61294 50314 62524
rect 53472 61942 53526 63180
rect 54242 62600 54324 63846
rect 57482 63256 57536 64420
rect 57332 63250 57596 63256
rect 54542 63238 57596 63250
rect 54404 63204 54420 63238
rect 54592 63204 55114 63238
rect 55286 63204 55808 63238
rect 55980 63204 56502 63238
rect 56674 63204 57196 63238
rect 57368 63204 57596 63238
rect 54542 63196 57596 63204
rect 57332 63180 57596 63196
rect 54238 62592 54558 62600
rect 54238 62580 57386 62592
rect 54238 62546 54420 62580
rect 54592 62546 55114 62580
rect 55286 62546 55808 62580
rect 55980 62546 56502 62580
rect 56674 62546 57196 62580
rect 57368 62546 57386 62580
rect 54238 62538 57386 62546
rect 54238 62524 54558 62538
rect 53292 61928 53556 61942
rect 50530 61922 53556 61928
rect 50394 61888 50410 61922
rect 50582 61888 51104 61922
rect 51276 61888 51798 61922
rect 51970 61888 52492 61922
rect 52664 61888 53186 61922
rect 53358 61888 53556 61922
rect 50530 61874 53556 61888
rect 53292 61866 53556 61874
rect 53472 61864 53526 61866
rect 54242 61294 54324 62524
rect 57482 61942 57536 63180
rect 71008 62774 71038 65520
rect 71178 62774 71224 65520
rect 71292 65408 71306 65580
rect 71340 65408 71348 65580
rect 71964 65580 71998 65596
rect 71292 64886 71348 65408
rect 71292 64714 71306 64886
rect 71340 64714 71348 64886
rect 71292 64192 71348 64714
rect 71292 64020 71306 64192
rect 71340 64020 71348 64192
rect 71292 63498 71348 64020
rect 71292 63326 71306 63498
rect 71340 63326 71348 63498
rect 71292 62838 71348 63326
rect 71008 62720 71224 62774
rect 71288 62804 71348 62838
rect 71288 62632 71306 62804
rect 71340 62632 71348 62804
rect 71954 65408 71964 65564
rect 72610 65580 72666 65686
rect 73920 65676 74106 65686
rect 75140 65708 75222 66382
rect 75808 66382 75828 66514
rect 75862 66470 75874 66554
rect 76472 69158 76486 69310
rect 76520 69278 76530 69330
rect 77144 69330 77178 69346
rect 76520 69158 76528 69278
rect 76472 68636 76528 69158
rect 76472 68464 76486 68636
rect 76520 68464 76528 68636
rect 76472 67942 76528 68464
rect 76472 67770 76486 67942
rect 76520 67770 76528 67942
rect 76472 67248 76528 67770
rect 76472 67076 76486 67248
rect 76520 67076 76528 67248
rect 76472 66554 76528 67076
rect 75862 66382 75868 66470
rect 76472 66466 76486 66554
rect 75808 66272 75868 66382
rect 76520 66466 76528 66554
rect 77132 69158 77144 69268
rect 77784 69330 77860 69426
rect 79006 69344 79062 69434
rect 77178 69158 77188 69268
rect 77784 69248 77802 69330
rect 77132 68636 77188 69158
rect 77132 68464 77144 68636
rect 77178 68464 77188 68636
rect 77132 67942 77188 68464
rect 77132 67770 77144 67942
rect 77178 67770 77188 67942
rect 77132 67248 77188 67770
rect 77132 67076 77144 67248
rect 77178 67076 77188 67248
rect 77132 66554 77188 67076
rect 77132 66424 77144 66554
rect 76486 66366 76520 66382
rect 77136 66382 77144 66424
rect 77178 66512 77188 66554
rect 77786 69158 77802 69248
rect 77836 69248 77860 69330
rect 78722 69284 78938 69344
rect 77836 69158 77842 69248
rect 77786 68636 77842 69158
rect 77786 68464 77802 68636
rect 77836 68464 77842 68636
rect 77786 67942 77842 68464
rect 77786 67770 77802 67942
rect 77836 67770 77842 67942
rect 77786 67248 77842 67770
rect 77786 67076 77802 67248
rect 77836 67076 77842 67248
rect 77786 66554 77842 67076
rect 77178 66382 77196 66512
rect 77786 66428 77802 66554
rect 77136 66276 77196 66382
rect 77836 66428 77842 66554
rect 78722 66538 78752 69284
rect 78892 66538 78938 69284
rect 79006 69172 79020 69344
rect 79054 69172 79062 69344
rect 79678 69344 79712 69360
rect 79006 68650 79062 69172
rect 79006 68478 79020 68650
rect 79054 68478 79062 68650
rect 79006 67956 79062 68478
rect 79006 67784 79020 67956
rect 79054 67784 79062 67956
rect 79006 67262 79062 67784
rect 79006 67090 79020 67262
rect 79054 67090 79062 67262
rect 79006 66568 79062 67090
rect 79006 66556 79020 66568
rect 78722 66484 78938 66538
rect 77802 66366 77836 66382
rect 78990 66396 79020 66556
rect 79054 66556 79062 66568
rect 79668 69172 79678 69328
rect 80324 69344 80380 69450
rect 81634 69440 81820 69450
rect 79712 69172 79724 69328
rect 80324 69324 80336 69344
rect 79668 68650 79724 69172
rect 79668 68478 79678 68650
rect 79712 68478 79724 68650
rect 79668 67956 79724 68478
rect 79668 67784 79678 67956
rect 79712 67784 79724 67956
rect 79668 67262 79724 67784
rect 79668 67090 79678 67262
rect 79712 67090 79724 67262
rect 79668 66568 79724 67090
rect 79054 66396 79072 66556
rect 79668 66528 79678 66568
rect 77136 66272 77294 66276
rect 75808 66210 77294 66272
rect 75808 66204 75868 66210
rect 77136 66202 77196 66210
rect 77792 65716 77970 65726
rect 77784 65708 77970 65716
rect 75140 65676 77970 65708
rect 78990 65722 79072 66396
rect 79658 66396 79678 66528
rect 79712 66484 79724 66568
rect 80322 69172 80336 69324
rect 80370 69292 80380 69344
rect 80994 69344 81028 69360
rect 80370 69172 80378 69292
rect 80322 68650 80378 69172
rect 80322 68478 80336 68650
rect 80370 68478 80378 68650
rect 80322 67956 80378 68478
rect 80322 67784 80336 67956
rect 80370 67784 80378 67956
rect 80322 67262 80378 67784
rect 80322 67090 80336 67262
rect 80370 67090 80378 67262
rect 80322 66568 80378 67090
rect 79712 66396 79718 66484
rect 80322 66480 80336 66568
rect 79658 66286 79718 66396
rect 80370 66480 80378 66568
rect 80982 69172 80994 69282
rect 81634 69344 81710 69440
rect 81028 69172 81038 69282
rect 81634 69262 81652 69344
rect 80982 68650 81038 69172
rect 80982 68478 80994 68650
rect 81028 68478 81038 68650
rect 80982 67956 81038 68478
rect 80982 67784 80994 67956
rect 81028 67784 81038 67956
rect 80982 67262 81038 67784
rect 80982 67090 80994 67262
rect 81028 67090 81038 67262
rect 80982 66568 81038 67090
rect 80982 66438 80994 66568
rect 80336 66380 80370 66396
rect 80986 66396 80994 66438
rect 81028 66526 81038 66568
rect 81636 69172 81652 69262
rect 81686 69262 81710 69344
rect 81686 69172 81692 69262
rect 81636 68650 81692 69172
rect 81636 68478 81652 68650
rect 81686 68478 81692 68650
rect 81636 67956 81692 68478
rect 81636 67784 81652 67956
rect 81686 67784 81692 67956
rect 81636 67262 81692 67784
rect 81636 67090 81652 67262
rect 81686 67090 81692 67262
rect 81636 66568 81692 67090
rect 81028 66396 81046 66526
rect 81636 66442 81652 66568
rect 80986 66290 81046 66396
rect 81686 66442 81692 66568
rect 81652 66380 81686 66396
rect 80986 66286 81144 66290
rect 79658 66224 81144 66286
rect 79658 66218 79718 66224
rect 80986 66216 81046 66224
rect 81642 65730 81820 65740
rect 81634 65722 81820 65730
rect 78990 65690 81820 65722
rect 79002 65680 81820 65690
rect 71998 65408 72010 65564
rect 72610 65560 72622 65580
rect 71954 64886 72010 65408
rect 71954 64714 71964 64886
rect 71998 64714 72010 64886
rect 71954 64192 72010 64714
rect 71954 64020 71964 64192
rect 71998 64020 72010 64192
rect 71954 63498 72010 64020
rect 71954 63326 71964 63498
rect 71998 63326 72010 63498
rect 71954 62804 72010 63326
rect 71954 62764 71964 62804
rect 71288 61964 71348 62632
rect 71944 62632 71964 62764
rect 71998 62720 72010 62804
rect 72608 65408 72622 65560
rect 72656 65528 72666 65580
rect 73280 65580 73314 65596
rect 72656 65408 72664 65528
rect 72608 64886 72664 65408
rect 72608 64714 72622 64886
rect 72656 64714 72664 64886
rect 72608 64192 72664 64714
rect 72608 64020 72622 64192
rect 72656 64020 72664 64192
rect 72608 63498 72664 64020
rect 72608 63326 72622 63498
rect 72656 63326 72664 63498
rect 72608 62804 72664 63326
rect 71998 62632 72004 62720
rect 72608 62716 72622 62804
rect 71944 62522 72004 62632
rect 72656 62716 72664 62804
rect 73268 65408 73280 65518
rect 73920 65580 73996 65676
rect 75152 65666 77970 65676
rect 73314 65408 73324 65518
rect 73920 65498 73938 65580
rect 73268 64886 73324 65408
rect 73268 64714 73280 64886
rect 73314 64714 73324 64886
rect 73268 64192 73324 64714
rect 73268 64020 73280 64192
rect 73314 64020 73324 64192
rect 73268 63498 73324 64020
rect 73268 63326 73280 63498
rect 73314 63326 73324 63498
rect 73268 62804 73324 63326
rect 73268 62674 73280 62804
rect 72622 62616 72656 62632
rect 73272 62632 73280 62674
rect 73314 62762 73324 62804
rect 73922 65408 73938 65498
rect 73972 65498 73996 65580
rect 75156 65560 75212 65666
rect 74872 65500 75088 65560
rect 73972 65408 73978 65498
rect 73922 64886 73978 65408
rect 73922 64714 73938 64886
rect 73972 64714 73978 64886
rect 73922 64192 73978 64714
rect 73922 64020 73938 64192
rect 73972 64020 73978 64192
rect 73922 63498 73978 64020
rect 73922 63326 73938 63498
rect 73972 63326 73978 63498
rect 73922 62804 73978 63326
rect 73314 62632 73332 62762
rect 73922 62678 73938 62804
rect 73272 62526 73332 62632
rect 73972 62678 73978 62804
rect 74872 62754 74902 65500
rect 75042 62754 75088 65500
rect 75156 65388 75170 65560
rect 75204 65388 75212 65560
rect 75828 65560 75862 65576
rect 75156 64866 75212 65388
rect 75156 64694 75170 64866
rect 75204 64694 75212 64866
rect 75156 64172 75212 64694
rect 75156 64000 75170 64172
rect 75204 64000 75212 64172
rect 75156 63478 75212 64000
rect 75156 63306 75170 63478
rect 75204 63306 75212 63478
rect 75156 62818 75212 63306
rect 74872 62700 75088 62754
rect 75152 62784 75212 62818
rect 73938 62616 73972 62632
rect 75152 62612 75170 62784
rect 75204 62612 75212 62784
rect 75818 65388 75828 65544
rect 76474 65560 76530 65666
rect 77784 65656 77970 65666
rect 75862 65388 75874 65544
rect 76474 65540 76486 65560
rect 75818 64866 75874 65388
rect 75818 64694 75828 64866
rect 75862 64694 75874 64866
rect 75818 64172 75874 64694
rect 75818 64000 75828 64172
rect 75862 64000 75874 64172
rect 75818 63478 75874 64000
rect 75818 63306 75828 63478
rect 75862 63306 75874 63478
rect 75818 62784 75874 63306
rect 75818 62744 75828 62784
rect 73272 62522 73430 62526
rect 71944 62460 73430 62522
rect 71944 62454 72004 62460
rect 73272 62452 73332 62460
rect 73928 61972 74106 61982
rect 73920 61964 74106 61972
rect 57302 61928 57566 61942
rect 54540 61922 57566 61928
rect 71288 61922 74106 61964
rect 54404 61888 54420 61922
rect 54592 61888 55114 61922
rect 55286 61888 55808 61922
rect 55980 61888 56502 61922
rect 56674 61888 57196 61922
rect 57368 61888 57566 61922
rect 54540 61874 57566 61888
rect 57302 61866 57566 61874
rect 46216 61286 46516 61294
rect 50228 61286 50528 61294
rect 54238 61286 54538 61294
rect 42194 61274 57254 61286
rect 42194 61266 57380 61274
rect 42194 61232 42390 61266
rect 42562 61232 43084 61266
rect 43256 61232 43778 61266
rect 43950 61232 44472 61266
rect 44644 61232 45166 61266
rect 45338 61264 57380 61266
rect 45338 61234 46398 61264
rect 45338 61232 45354 61234
rect 42194 61222 45350 61232
rect 46216 61230 46398 61234
rect 46570 61230 47092 61264
rect 47264 61230 47786 61264
rect 47958 61230 48480 61264
rect 48652 61230 49174 61264
rect 49346 61234 50410 61264
rect 49346 61230 49362 61234
rect 50228 61230 50410 61234
rect 50582 61230 51104 61264
rect 51276 61230 51798 61264
rect 51970 61230 52492 61264
rect 52664 61230 53186 61264
rect 53358 61234 54420 61264
rect 53358 61230 53374 61234
rect 54238 61230 54420 61234
rect 54592 61230 55114 61264
rect 55286 61230 55808 61264
rect 55980 61230 56502 61264
rect 56674 61230 57196 61264
rect 57368 61230 57384 61264
rect 42194 61220 42490 61222
rect 46216 61220 49358 61230
rect 50228 61220 53370 61230
rect 54238 61220 57380 61230
rect 42194 61218 42294 61220
rect 46216 61218 46498 61220
rect 50228 61218 50510 61220
rect 54238 61218 54520 61220
rect 5152 60246 5374 60258
rect 7826 60252 8048 60264
rect 10472 60252 10694 60264
rect 11700 60258 13348 60268
rect 14354 60264 16002 60274
rect 16980 60268 18628 60278
rect 13126 60246 13348 60258
rect 15780 60252 16002 60264
rect 18406 60256 18628 60268
rect 18240 59700 18680 59802
rect 42194 59726 42276 61218
rect 46220 61216 46302 61218
rect 50232 61216 50314 61218
rect 54242 61216 54324 61218
rect 42726 60862 45372 60898
rect 42726 60530 42876 60862
rect 45276 60530 45372 60862
rect 42726 60496 45372 60530
rect 46720 60862 49366 60898
rect 46720 60530 46870 60862
rect 49270 60530 49366 60862
rect 46720 60496 49366 60530
rect 50742 60862 53388 60898
rect 50742 60530 50892 60862
rect 53292 60530 53388 60862
rect 50742 60496 53388 60530
rect 54764 60862 57410 60898
rect 54764 60530 54914 60862
rect 57314 60530 57410 60862
rect 54764 60496 57410 60530
rect 57478 60388 57564 61866
rect 71292 61816 71348 61922
rect 71008 61756 71224 61816
rect 57706 61190 58040 61298
rect 57706 60506 57780 61190
rect 57972 60506 58040 61190
rect 57706 60396 58040 60506
rect 45258 60370 45522 60388
rect 49252 60370 49516 60388
rect 53274 60370 53538 60388
rect 57296 60370 57564 60388
rect 42456 60358 57564 60370
rect 42366 60324 42382 60358
rect 42554 60324 43076 60358
rect 43248 60324 43770 60358
rect 43942 60324 44464 60358
rect 44636 60324 45158 60358
rect 45330 60324 46376 60358
rect 46548 60324 47070 60358
rect 47242 60324 47764 60358
rect 47936 60324 48458 60358
rect 48630 60324 49152 60358
rect 49324 60324 50398 60358
rect 50570 60324 51092 60358
rect 51264 60324 51786 60358
rect 51958 60324 52480 60358
rect 52652 60324 53174 60358
rect 53346 60324 54420 60358
rect 54592 60324 55114 60358
rect 55286 60324 55808 60358
rect 55980 60324 56502 60358
rect 56674 60324 57196 60358
rect 57368 60324 57564 60358
rect 42456 60320 57564 60324
rect 42456 60318 57560 60320
rect 42456 60316 45522 60318
rect 46450 60316 49516 60318
rect 50472 60316 53538 60318
rect 54494 60316 57560 60318
rect 45258 60312 45522 60316
rect 49252 60312 49516 60316
rect 53274 60312 53538 60316
rect 57296 60312 57560 60316
rect 944 59660 2576 59694
rect 944 59518 1000 59660
rect 2514 59518 2576 59660
rect 944 59490 2576 59518
rect 3612 59656 5244 59690
rect 3612 59514 3668 59656
rect 5182 59514 5244 59656
rect 3612 59486 5244 59514
rect 6286 59662 7918 59696
rect 6286 59520 6342 59662
rect 7856 59520 7918 59662
rect 6286 59492 7918 59520
rect 8932 59662 10564 59696
rect 8932 59520 8988 59662
rect 10502 59520 10564 59662
rect 8932 59492 10564 59520
rect 11586 59656 13218 59690
rect 11586 59514 11642 59656
rect 13156 59514 13218 59656
rect 11586 59486 13218 59514
rect 14240 59662 15872 59696
rect 14240 59520 14296 59662
rect 15810 59520 15872 59662
rect 14240 59492 15872 59520
rect 16866 59666 18680 59700
rect 16866 59524 16922 59666
rect 18436 59542 18680 59666
rect 19364 59702 20600 59726
rect 18436 59524 18498 59542
rect 16866 59496 18498 59524
rect 19364 59508 19472 59702
rect 20538 59508 20600 59702
rect 42194 59712 42490 59726
rect 42194 59700 45340 59712
rect 42194 59666 42382 59700
rect 42554 59666 43076 59700
rect 43248 59666 43770 59700
rect 43942 59666 44464 59700
rect 44636 59666 45158 59700
rect 45330 59666 45346 59700
rect 42194 59658 45340 59666
rect 42194 59650 42490 59658
rect 42194 59550 42286 59650
rect 19364 59456 20600 59508
rect 2360 59384 20528 59414
rect 2360 59352 20840 59384
rect 2360 59320 19544 59352
rect 908 59318 19544 59320
rect 19716 59318 20238 59352
rect 20410 59318 20840 59352
rect 908 59308 20840 59318
rect 908 59304 16860 59308
rect 908 59302 6280 59304
rect 908 59268 938 59302
rect 1110 59268 1632 59302
rect 1804 59268 2326 59302
rect 2498 59298 6280 59302
rect 2498 59268 3606 59298
rect 908 59264 3606 59268
rect 3778 59264 4300 59298
rect 4472 59264 4994 59298
rect 5166 59270 6280 59298
rect 6452 59270 6974 59304
rect 7146 59270 7668 59304
rect 7840 59270 8926 59304
rect 9098 59270 9620 59304
rect 9792 59270 10314 59304
rect 10486 59298 14234 59304
rect 10486 59270 11580 59298
rect 5166 59264 11580 59270
rect 11752 59264 12274 59298
rect 12446 59264 12968 59298
rect 13140 59270 14234 59298
rect 14406 59270 14928 59304
rect 15100 59270 15622 59304
rect 15794 59274 16860 59304
rect 17032 59274 17554 59308
rect 17726 59274 18248 59308
rect 18420 59274 20840 59308
rect 15794 59270 20840 59274
rect 13140 59264 20840 59270
rect 908 59256 20840 59264
rect 2360 59244 20840 59256
rect 746 58656 1066 58678
rect 746 58654 2474 58656
rect 728 58644 2474 58654
rect 728 58610 938 58644
rect 1110 58610 1632 58644
rect 1804 58610 2326 58644
rect 2498 58610 2514 58644
rect 728 58604 2474 58610
rect 728 58556 1066 58604
rect 222 57816 554 57874
rect 222 56666 280 57816
rect 496 57298 554 57816
rect 728 57356 820 58556
rect 2610 57994 2678 59244
rect 3414 58652 3734 58674
rect 3414 58650 5142 58652
rect 956 57986 2678 57994
rect 922 57952 938 57986
rect 1110 57952 1632 57986
rect 1804 57952 2326 57986
rect 2498 57952 2678 57986
rect 956 57942 2678 57952
rect 2390 57940 2678 57942
rect 728 57334 1052 57356
rect 728 57328 2478 57334
rect 728 57298 938 57328
rect 496 57294 938 57298
rect 1110 57294 1632 57328
rect 1804 57294 2326 57328
rect 2498 57294 2514 57328
rect 496 57282 2478 57294
rect 496 57234 1052 57282
rect 496 57184 854 57234
rect 496 56666 554 57184
rect 222 56552 554 56666
rect 728 56042 820 57184
rect 2610 56682 2678 57940
rect 2402 56680 2678 56682
rect 970 56670 2678 56680
rect 922 56636 938 56670
rect 1110 56636 1632 56670
rect 1804 56636 2326 56670
rect 2498 56636 2678 56670
rect 970 56628 2678 56636
rect 722 56020 1042 56042
rect 722 56012 2488 56020
rect 722 55978 938 56012
rect 1110 55978 1632 56012
rect 1804 55978 2326 56012
rect 2498 55978 2514 56012
rect 722 55968 2488 55978
rect 722 55920 1042 55968
rect 728 54754 820 55920
rect 2610 55364 2678 56628
rect 3396 58640 5142 58650
rect 3396 58606 3606 58640
rect 3778 58606 4300 58640
rect 4472 58606 4994 58640
rect 5166 58606 5182 58640
rect 3396 58600 5142 58606
rect 3396 58552 3734 58600
rect 3396 57352 3488 58552
rect 5278 57990 5346 59244
rect 6088 58658 6408 58680
rect 6088 58656 7816 58658
rect 3624 57982 5346 57990
rect 3590 57948 3606 57982
rect 3778 57948 4300 57982
rect 4472 57948 4994 57982
rect 5166 57948 5346 57982
rect 3624 57938 5346 57948
rect 5058 57936 5346 57938
rect 3396 57330 3720 57352
rect 3396 57324 5146 57330
rect 3396 57290 3606 57324
rect 3778 57290 4300 57324
rect 4472 57290 4994 57324
rect 5166 57290 5182 57324
rect 3396 57278 5146 57290
rect 3396 57230 3720 57278
rect 3396 56038 3488 57230
rect 5278 56678 5346 57936
rect 5070 56676 5346 56678
rect 3638 56666 5346 56676
rect 3590 56632 3606 56666
rect 3778 56632 4300 56666
rect 4472 56632 4994 56666
rect 5166 56632 5346 56666
rect 3638 56624 5346 56632
rect 3390 56016 3710 56038
rect 3390 56008 5156 56016
rect 3390 55974 3606 56008
rect 3778 55974 4300 56008
rect 4472 55974 4994 56008
rect 5166 55974 5182 56008
rect 3390 55964 5156 55974
rect 3390 55916 3710 55964
rect 2392 55362 2678 55364
rect 994 55354 2678 55362
rect 922 55320 938 55354
rect 1110 55320 1632 55354
rect 1804 55320 2326 55354
rect 2498 55320 2678 55354
rect 994 55310 2678 55320
rect 712 54706 1032 54754
rect 712 54696 2536 54706
rect 712 54662 938 54696
rect 1110 54662 1632 54696
rect 1804 54662 2326 54696
rect 2498 54662 2536 54696
rect 2610 54678 2678 55310
rect 712 54654 2536 54662
rect 712 54632 1032 54654
rect 2600 54636 2678 54678
rect 2600 54052 2674 54636
rect 3396 54750 3488 55916
rect 5278 55360 5346 56624
rect 6070 58646 7816 58656
rect 6070 58612 6280 58646
rect 6452 58612 6974 58646
rect 7146 58612 7668 58646
rect 7840 58612 7856 58646
rect 6070 58606 7816 58612
rect 6070 58558 6408 58606
rect 6070 57358 6162 58558
rect 7952 57996 8020 59244
rect 8734 58658 9054 58680
rect 8734 58656 10462 58658
rect 6298 57988 8020 57996
rect 6264 57954 6280 57988
rect 6452 57954 6974 57988
rect 7146 57954 7668 57988
rect 7840 57954 8020 57988
rect 6298 57944 8020 57954
rect 7732 57942 8020 57944
rect 6070 57336 6394 57358
rect 6070 57330 7820 57336
rect 6070 57296 6280 57330
rect 6452 57296 6974 57330
rect 7146 57296 7668 57330
rect 7840 57296 7856 57330
rect 6070 57284 7820 57296
rect 6070 57236 6394 57284
rect 6070 56044 6162 57236
rect 7952 56684 8020 57942
rect 7744 56682 8020 56684
rect 6312 56672 8020 56682
rect 6264 56638 6280 56672
rect 6452 56638 6974 56672
rect 7146 56638 7668 56672
rect 7840 56638 8020 56672
rect 6312 56630 8020 56638
rect 6064 56022 6384 56044
rect 6064 56014 7830 56022
rect 6064 55980 6280 56014
rect 6452 55980 6974 56014
rect 7146 55980 7668 56014
rect 7840 55980 7856 56014
rect 6064 55970 7830 55980
rect 6064 55922 6384 55970
rect 5060 55358 5346 55360
rect 3662 55350 5346 55358
rect 3590 55316 3606 55350
rect 3778 55316 4300 55350
rect 4472 55316 4994 55350
rect 5166 55316 5346 55350
rect 3662 55306 5346 55316
rect 3380 54742 3700 54750
rect 3276 54702 3700 54742
rect 3276 54692 5204 54702
rect 3276 54658 3606 54692
rect 3778 54658 4300 54692
rect 4472 54658 4994 54692
rect 5166 54658 5204 54692
rect 5278 54674 5346 55306
rect 3276 54650 5204 54658
rect 3276 54628 3700 54650
rect 5268 54632 5346 54674
rect 3276 54600 3504 54628
rect 2456 54046 2678 54052
rect 5268 54048 5342 54632
rect 6070 54756 6162 55922
rect 7952 55366 8020 56630
rect 8716 58646 10462 58656
rect 8716 58612 8926 58646
rect 9098 58612 9620 58646
rect 9792 58612 10314 58646
rect 10486 58612 10502 58646
rect 8716 58606 10462 58612
rect 8716 58558 9054 58606
rect 8716 57358 8808 58558
rect 10598 57996 10666 59244
rect 11388 58652 11708 58674
rect 11388 58650 13116 58652
rect 8944 57988 10666 57996
rect 8910 57954 8926 57988
rect 9098 57954 9620 57988
rect 9792 57954 10314 57988
rect 10486 57954 10666 57988
rect 8944 57944 10666 57954
rect 10378 57942 10666 57944
rect 8716 57336 9040 57358
rect 8716 57330 10466 57336
rect 8716 57296 8926 57330
rect 9098 57296 9620 57330
rect 9792 57296 10314 57330
rect 10486 57296 10502 57330
rect 8716 57284 10466 57296
rect 8716 57236 9040 57284
rect 8716 56044 8808 57236
rect 10598 56684 10666 57942
rect 10390 56682 10666 56684
rect 8958 56672 10666 56682
rect 8910 56638 8926 56672
rect 9098 56638 9620 56672
rect 9792 56638 10314 56672
rect 10486 56638 10666 56672
rect 8958 56630 10666 56638
rect 8710 56022 9030 56044
rect 8710 56014 10476 56022
rect 8710 55980 8926 56014
rect 9098 55980 9620 56014
rect 9792 55980 10314 56014
rect 10486 55980 10502 56014
rect 8710 55970 10476 55980
rect 8710 55922 9030 55970
rect 7734 55364 8020 55366
rect 6336 55356 8020 55364
rect 6264 55322 6280 55356
rect 6452 55322 6974 55356
rect 7146 55322 7668 55356
rect 7840 55322 8020 55356
rect 6336 55312 8020 55322
rect 6054 54752 6374 54756
rect 5928 54708 6374 54752
rect 5928 54698 7878 54708
rect 5928 54664 6280 54698
rect 6452 54664 6974 54698
rect 7146 54664 7668 54698
rect 7840 54664 7878 54698
rect 7952 54680 8020 55312
rect 5928 54656 7878 54664
rect 5928 54642 6374 54656
rect 6054 54634 6374 54642
rect 7942 54638 8020 54680
rect 7942 54054 8016 54638
rect 8716 54768 8808 55922
rect 10598 55366 10666 56630
rect 11370 58640 13116 58650
rect 11370 58606 11580 58640
rect 11752 58606 12274 58640
rect 12446 58606 12968 58640
rect 13140 58606 13156 58640
rect 11370 58600 13116 58606
rect 11370 58552 11708 58600
rect 11370 57352 11462 58552
rect 13252 57990 13320 59244
rect 14042 58658 14362 58680
rect 14042 58656 15770 58658
rect 11598 57982 13320 57990
rect 11564 57948 11580 57982
rect 11752 57948 12274 57982
rect 12446 57948 12968 57982
rect 13140 57948 13320 57982
rect 11598 57938 13320 57948
rect 13032 57936 13320 57938
rect 11370 57330 11694 57352
rect 11370 57324 13120 57330
rect 11370 57290 11580 57324
rect 11752 57290 12274 57324
rect 12446 57290 12968 57324
rect 13140 57290 13156 57324
rect 11370 57278 13120 57290
rect 11370 57230 11694 57278
rect 11370 56038 11462 57230
rect 13252 56678 13320 57936
rect 13044 56676 13320 56678
rect 11612 56666 13320 56676
rect 11564 56632 11580 56666
rect 11752 56632 12274 56666
rect 12446 56632 12968 56666
rect 13140 56632 13320 56666
rect 11612 56624 13320 56632
rect 11364 56016 11684 56038
rect 11364 56008 13130 56016
rect 11364 55974 11580 56008
rect 11752 55974 12274 56008
rect 12446 55974 12968 56008
rect 13140 55974 13156 56008
rect 11364 55964 13130 55974
rect 11364 55916 11684 55964
rect 10380 55364 10666 55366
rect 8982 55356 10666 55364
rect 8910 55322 8926 55356
rect 9098 55322 9620 55356
rect 9792 55322 10314 55356
rect 10486 55322 10666 55356
rect 8982 55312 10666 55322
rect 8554 54756 8822 54768
rect 8554 54708 9020 54756
rect 8554 54698 10524 54708
rect 8554 54664 8926 54698
rect 9098 54664 9620 54698
rect 9792 54664 10314 54698
rect 10486 54664 10524 54698
rect 10598 54680 10666 55312
rect 8554 54656 10524 54664
rect 8554 54642 9020 54656
rect 8700 54634 9020 54642
rect 10588 54638 10666 54680
rect 10588 54054 10662 54638
rect 11370 54760 11462 55916
rect 13252 55360 13320 56624
rect 14024 58646 15770 58656
rect 14024 58612 14234 58646
rect 14406 58612 14928 58646
rect 15100 58612 15622 58646
rect 15794 58612 15810 58646
rect 14024 58606 15770 58612
rect 14024 58558 14362 58606
rect 14024 57358 14116 58558
rect 15906 57996 15974 59244
rect 16668 58662 16988 58684
rect 16668 58660 18396 58662
rect 14252 57988 15974 57996
rect 14218 57954 14234 57988
rect 14406 57954 14928 57988
rect 15100 57954 15622 57988
rect 15794 57954 15974 57988
rect 14252 57944 15974 57954
rect 15686 57942 15974 57944
rect 14024 57336 14348 57358
rect 14024 57330 15774 57336
rect 14024 57296 14234 57330
rect 14406 57296 14928 57330
rect 15100 57296 15622 57330
rect 15794 57296 15810 57330
rect 14024 57284 15774 57296
rect 14024 57236 14348 57284
rect 14024 56044 14116 57236
rect 15906 56684 15974 57942
rect 15698 56682 15974 56684
rect 14266 56672 15974 56682
rect 14218 56638 14234 56672
rect 14406 56638 14928 56672
rect 15100 56638 15622 56672
rect 15794 56638 15974 56672
rect 14266 56630 15974 56638
rect 14018 56022 14338 56044
rect 14018 56014 15784 56022
rect 14018 55980 14234 56014
rect 14406 55980 14928 56014
rect 15100 55980 15622 56014
rect 15794 55980 15810 56014
rect 14018 55970 15784 55980
rect 14018 55922 14338 55970
rect 13034 55358 13320 55360
rect 11636 55350 13320 55358
rect 11564 55316 11580 55350
rect 11752 55316 12274 55350
rect 12446 55316 12968 55350
rect 13140 55316 13320 55350
rect 11636 55306 13320 55316
rect 11246 54702 11920 54760
rect 11246 54692 13178 54702
rect 11246 54658 11580 54692
rect 11752 54658 12274 54692
rect 12446 54658 12968 54692
rect 13140 54658 13178 54692
rect 13252 54674 13320 55306
rect 11246 54650 13178 54658
rect 11246 54642 11920 54650
rect 11354 54628 11674 54642
rect 13242 54632 13320 54674
rect 7798 54048 8020 54054
rect 10444 54048 10666 54054
rect 13242 54048 13316 54632
rect 14024 54756 14116 55922
rect 15906 55366 15974 56630
rect 16650 58650 18396 58660
rect 16650 58616 16860 58650
rect 17032 58616 17554 58650
rect 17726 58616 18248 58650
rect 18420 58616 18436 58650
rect 16650 58610 18396 58616
rect 16650 58562 16988 58610
rect 16650 57362 16742 58562
rect 18532 58000 18600 59244
rect 20430 59236 20840 59244
rect 19336 58710 19618 58720
rect 19336 58694 20414 58710
rect 19336 58660 19544 58694
rect 19716 58660 20238 58694
rect 20410 58660 20426 58694
rect 19336 58652 20414 58660
rect 19336 58624 19618 58652
rect 16878 57992 18600 58000
rect 16844 57958 16860 57992
rect 17032 57958 17554 57992
rect 17726 57958 18248 57992
rect 18420 57958 18600 57992
rect 16878 57948 18600 57958
rect 18312 57946 18600 57948
rect 16650 57340 16974 57362
rect 16650 57334 18400 57340
rect 16650 57300 16860 57334
rect 17032 57300 17554 57334
rect 17726 57300 18248 57334
rect 18420 57300 18436 57334
rect 16650 57288 18400 57300
rect 16650 57240 16974 57288
rect 16650 56048 16742 57240
rect 18532 56688 18600 57946
rect 18324 56686 18600 56688
rect 16892 56676 18600 56686
rect 16844 56642 16860 56676
rect 17032 56642 17554 56676
rect 17726 56642 18248 56676
rect 18420 56642 18600 56676
rect 16892 56634 18600 56642
rect 16644 56026 16964 56048
rect 16644 56018 18410 56026
rect 16644 55984 16860 56018
rect 17032 55984 17554 56018
rect 17726 55984 18248 56018
rect 18420 55984 18436 56018
rect 16644 55974 18410 55984
rect 16644 55926 16964 55974
rect 15688 55364 15974 55366
rect 14290 55356 15974 55364
rect 14218 55322 14234 55356
rect 14406 55322 14928 55356
rect 15100 55322 15622 55356
rect 15794 55322 15974 55356
rect 14290 55312 15974 55322
rect 14008 54734 14328 54756
rect 13846 54708 14460 54734
rect 13846 54698 15832 54708
rect 13846 54664 14234 54698
rect 14406 54664 14928 54698
rect 15100 54664 15622 54698
rect 15794 54664 15832 54698
rect 15906 54680 15974 55312
rect 13846 54656 15832 54664
rect 13846 54616 14460 54656
rect 15896 54638 15974 54680
rect 15896 54054 15970 54638
rect 16650 54768 16742 55926
rect 18532 55370 18600 56634
rect 19352 57404 19420 58624
rect 19612 58040 20414 58046
rect 20478 58040 20560 59236
rect 42204 58404 42286 59550
rect 45444 59060 45498 60312
rect 46198 59712 46484 59726
rect 46198 59700 49334 59712
rect 46198 59666 46376 59700
rect 46548 59666 47070 59700
rect 47242 59666 47764 59700
rect 47936 59666 48458 59700
rect 48630 59666 49152 59700
rect 49324 59666 49340 59700
rect 46198 59658 49334 59666
rect 46198 59650 46484 59658
rect 45294 59054 45558 59060
rect 42504 59042 45558 59054
rect 42366 59008 42382 59042
rect 42554 59008 43076 59042
rect 43248 59008 43770 59042
rect 43942 59008 44464 59042
rect 44636 59008 45158 59042
rect 45330 59008 45558 59042
rect 42504 59000 45558 59008
rect 45294 58984 45558 59000
rect 42200 58396 42520 58404
rect 42200 58384 45348 58396
rect 42200 58350 42382 58384
rect 42554 58350 43076 58384
rect 43248 58350 43770 58384
rect 43942 58350 44464 58384
rect 44636 58350 45158 58384
rect 45330 58350 45348 58384
rect 42200 58342 45348 58350
rect 42200 58328 42520 58342
rect 19612 58036 20560 58040
rect 19528 58002 19544 58036
rect 19716 58002 20238 58036
rect 20410 58002 20560 58036
rect 19612 57988 20560 58002
rect 20304 57970 20560 57988
rect 19352 57394 19638 57404
rect 19352 57378 20422 57394
rect 19352 57344 19544 57378
rect 19716 57344 20238 57378
rect 20410 57344 20426 57378
rect 19352 57336 20422 57344
rect 19352 57308 19638 57336
rect 19352 56076 19420 57308
rect 19624 56722 20426 56726
rect 20478 56722 20560 57970
rect 30150 57488 30206 57492
rect 30022 57486 30208 57488
rect 23726 57480 30208 57486
rect 23618 57446 23634 57480
rect 23806 57446 24328 57480
rect 24500 57446 25022 57480
rect 25194 57446 25716 57480
rect 25888 57446 26410 57480
rect 26582 57446 27104 57480
rect 27276 57446 27798 57480
rect 27970 57446 28492 57480
rect 28664 57446 29186 57480
rect 29358 57446 29880 57480
rect 30052 57446 30208 57480
rect 23726 57432 30208 57446
rect 23726 57424 30040 57432
rect 30150 56832 30206 57432
rect 42204 57098 42286 58328
rect 45444 57746 45498 58984
rect 46198 58404 46280 59650
rect 49438 59060 49492 60312
rect 50220 59712 50506 59726
rect 50220 59700 53356 59712
rect 50220 59666 50398 59700
rect 50570 59666 51092 59700
rect 51264 59666 51786 59700
rect 51958 59666 52480 59700
rect 52652 59666 53174 59700
rect 53346 59666 53362 59700
rect 50220 59658 53356 59666
rect 50220 59650 50506 59658
rect 49288 59054 49552 59060
rect 46498 59042 49552 59054
rect 46360 59008 46376 59042
rect 46548 59008 47070 59042
rect 47242 59008 47764 59042
rect 47936 59008 48458 59042
rect 48630 59008 49152 59042
rect 49324 59008 49552 59042
rect 46498 59000 49552 59008
rect 49288 58984 49552 59000
rect 46194 58396 46514 58404
rect 46194 58384 49342 58396
rect 46194 58350 46376 58384
rect 46548 58350 47070 58384
rect 47242 58350 47764 58384
rect 47936 58350 48458 58384
rect 48630 58350 49152 58384
rect 49324 58350 49342 58384
rect 46194 58342 49342 58350
rect 46194 58328 46514 58342
rect 45264 57732 45528 57746
rect 42502 57726 45528 57732
rect 42366 57692 42382 57726
rect 42554 57692 43076 57726
rect 43248 57692 43770 57726
rect 43942 57692 44464 57726
rect 44636 57692 45158 57726
rect 45330 57692 45528 57726
rect 42502 57678 45528 57692
rect 45264 57670 45528 57678
rect 45444 57668 45498 57670
rect 46198 57098 46280 58328
rect 49438 57746 49492 58984
rect 50220 58404 50302 59650
rect 53460 59060 53514 60312
rect 57442 60170 57536 60312
rect 54242 59712 54528 59726
rect 54242 59700 57378 59712
rect 54242 59666 54420 59700
rect 54592 59666 55114 59700
rect 55286 59666 55808 59700
rect 55980 59666 56502 59700
rect 56674 59666 57196 59700
rect 57368 59666 57384 59700
rect 54242 59658 57378 59666
rect 54242 59650 54528 59658
rect 53310 59054 53574 59060
rect 50520 59042 53574 59054
rect 50382 59008 50398 59042
rect 50570 59008 51092 59042
rect 51264 59008 51786 59042
rect 51958 59008 52480 59042
rect 52652 59008 53174 59042
rect 53346 59008 53574 59042
rect 50520 59000 53574 59008
rect 53310 58984 53574 59000
rect 50216 58396 50536 58404
rect 50216 58384 53364 58396
rect 50216 58350 50398 58384
rect 50570 58350 51092 58384
rect 51264 58350 51786 58384
rect 51958 58350 52480 58384
rect 52652 58350 53174 58384
rect 53346 58350 53364 58384
rect 50216 58342 53364 58350
rect 50216 58328 50536 58342
rect 49258 57732 49522 57746
rect 46496 57726 49522 57732
rect 46360 57692 46376 57726
rect 46548 57692 47070 57726
rect 47242 57692 47764 57726
rect 47936 57692 48458 57726
rect 48630 57692 49152 57726
rect 49324 57692 49522 57726
rect 46496 57678 49522 57692
rect 49258 57670 49522 57678
rect 49438 57668 49492 57670
rect 50220 57098 50302 58328
rect 53460 57746 53514 58984
rect 54242 58404 54324 59650
rect 57482 59060 57536 60170
rect 57332 59054 57596 59060
rect 54542 59042 57596 59054
rect 54404 59008 54420 59042
rect 54592 59008 55114 59042
rect 55286 59008 55808 59042
rect 55980 59008 56502 59042
rect 56674 59008 57196 59042
rect 57368 59008 57596 59042
rect 54542 59000 57596 59008
rect 57332 58984 57596 59000
rect 71008 59010 71038 61756
rect 71178 59010 71224 61756
rect 71292 61644 71306 61816
rect 71340 61644 71348 61816
rect 71964 61816 71998 61832
rect 71292 61122 71348 61644
rect 71292 60950 71306 61122
rect 71340 60950 71348 61122
rect 71292 60428 71348 60950
rect 71292 60256 71306 60428
rect 71340 60256 71348 60428
rect 71292 59734 71348 60256
rect 71292 59562 71306 59734
rect 71340 59562 71348 59734
rect 71292 59156 71348 59562
rect 71954 61644 71964 61800
rect 72610 61816 72666 61922
rect 73920 61912 74106 61922
rect 75152 61944 75212 62612
rect 75808 62612 75828 62744
rect 75862 62700 75874 62784
rect 76472 65388 76486 65540
rect 76520 65508 76530 65560
rect 77144 65560 77178 65576
rect 76520 65388 76528 65508
rect 76472 64866 76528 65388
rect 76472 64694 76486 64866
rect 76520 64694 76528 64866
rect 76472 64172 76528 64694
rect 76472 64000 76486 64172
rect 76520 64000 76528 64172
rect 76472 63478 76528 64000
rect 76472 63306 76486 63478
rect 76520 63306 76528 63478
rect 76472 62784 76528 63306
rect 75862 62612 75868 62700
rect 76472 62696 76486 62784
rect 75808 62502 75868 62612
rect 76520 62696 76528 62784
rect 77132 65388 77144 65498
rect 77784 65560 77860 65656
rect 79006 65574 79062 65680
rect 77178 65388 77188 65498
rect 77784 65478 77802 65560
rect 77132 64866 77188 65388
rect 77132 64694 77144 64866
rect 77178 64694 77188 64866
rect 77132 64172 77188 64694
rect 77132 64000 77144 64172
rect 77178 64000 77188 64172
rect 77132 63478 77188 64000
rect 77132 63306 77144 63478
rect 77178 63306 77188 63478
rect 77132 62784 77188 63306
rect 77132 62654 77144 62784
rect 76486 62596 76520 62612
rect 77136 62612 77144 62654
rect 77178 62742 77188 62784
rect 77786 65388 77802 65478
rect 77836 65478 77860 65560
rect 78722 65514 78938 65574
rect 77836 65388 77842 65478
rect 77786 64866 77842 65388
rect 77786 64694 77802 64866
rect 77836 64694 77842 64866
rect 77786 64172 77842 64694
rect 77786 64000 77802 64172
rect 77836 64000 77842 64172
rect 77786 63478 77842 64000
rect 77786 63306 77802 63478
rect 77836 63306 77842 63478
rect 77786 62784 77842 63306
rect 77178 62612 77196 62742
rect 77786 62658 77802 62784
rect 77136 62506 77196 62612
rect 77836 62658 77842 62784
rect 78722 62768 78752 65514
rect 78892 62768 78938 65514
rect 79006 65402 79020 65574
rect 79054 65402 79062 65574
rect 79678 65574 79712 65590
rect 79006 64880 79062 65402
rect 79006 64708 79020 64880
rect 79054 64708 79062 64880
rect 79006 64186 79062 64708
rect 79006 64014 79020 64186
rect 79054 64014 79062 64186
rect 79006 63492 79062 64014
rect 79006 63320 79020 63492
rect 79054 63320 79062 63492
rect 79006 62832 79062 63320
rect 78722 62714 78938 62768
rect 79002 62798 79062 62832
rect 77802 62596 77836 62612
rect 79002 62626 79020 62798
rect 79054 62626 79062 62798
rect 79668 65402 79678 65558
rect 80324 65574 80380 65680
rect 81634 65670 81820 65680
rect 79712 65402 79724 65558
rect 80324 65554 80336 65574
rect 79668 64880 79724 65402
rect 79668 64708 79678 64880
rect 79712 64708 79724 64880
rect 79668 64186 79724 64708
rect 79668 64014 79678 64186
rect 79712 64014 79724 64186
rect 79668 63492 79724 64014
rect 79668 63320 79678 63492
rect 79712 63320 79724 63492
rect 79668 62798 79724 63320
rect 79668 62758 79678 62798
rect 77136 62502 77294 62506
rect 75808 62440 77294 62502
rect 75808 62434 75868 62440
rect 77136 62432 77196 62440
rect 77792 61952 77970 61962
rect 77784 61944 77970 61952
rect 71998 61644 72010 61800
rect 72610 61796 72622 61816
rect 71954 61122 72010 61644
rect 71954 60950 71964 61122
rect 71998 60950 72010 61122
rect 71954 60428 72010 60950
rect 71954 60256 71964 60428
rect 71998 60256 72010 60428
rect 71954 59734 72010 60256
rect 71954 59562 71964 59734
rect 71998 59562 72010 59734
rect 54238 58396 54558 58404
rect 54238 58384 57386 58396
rect 54238 58350 54420 58384
rect 54592 58350 55114 58384
rect 55286 58350 55808 58384
rect 55980 58350 56502 58384
rect 56674 58350 57196 58384
rect 57368 58350 57386 58384
rect 54238 58342 57386 58350
rect 54238 58328 54558 58342
rect 53280 57732 53544 57746
rect 50518 57726 53544 57732
rect 50382 57692 50398 57726
rect 50570 57692 51092 57726
rect 51264 57692 51786 57726
rect 51958 57692 52480 57726
rect 52652 57692 53174 57726
rect 53346 57692 53544 57726
rect 50518 57678 53544 57692
rect 53280 57670 53544 57678
rect 53460 57668 53514 57670
rect 54242 57098 54324 58328
rect 57482 57746 57536 58984
rect 71008 58956 71224 59010
rect 71288 59040 71364 59156
rect 71288 58868 71306 59040
rect 71340 58868 71364 59040
rect 71954 59040 72010 59562
rect 71954 59000 71964 59040
rect 71288 58188 71364 58868
rect 71944 58868 71964 59000
rect 71998 58956 72010 59040
rect 72608 61644 72622 61796
rect 72656 61764 72666 61816
rect 73280 61816 73314 61832
rect 72656 61644 72664 61764
rect 72608 61122 72664 61644
rect 72608 60950 72622 61122
rect 72656 60950 72664 61122
rect 72608 60428 72664 60950
rect 72608 60256 72622 60428
rect 72656 60256 72664 60428
rect 72608 59734 72664 60256
rect 72608 59562 72622 59734
rect 72656 59562 72664 59734
rect 72608 59040 72664 59562
rect 71998 58868 72004 58956
rect 72608 58952 72622 59040
rect 71944 58758 72004 58868
rect 72656 58952 72664 59040
rect 73268 61644 73280 61754
rect 73920 61816 73996 61912
rect 75152 61902 77970 61944
rect 79002 61958 79062 62626
rect 79658 62626 79678 62758
rect 79712 62714 79724 62798
rect 80322 65402 80336 65554
rect 80370 65522 80380 65574
rect 80994 65574 81028 65590
rect 80370 65402 80378 65522
rect 80322 64880 80378 65402
rect 80322 64708 80336 64880
rect 80370 64708 80378 64880
rect 80322 64186 80378 64708
rect 80322 64014 80336 64186
rect 80370 64014 80378 64186
rect 80322 63492 80378 64014
rect 80322 63320 80336 63492
rect 80370 63320 80378 63492
rect 80322 62798 80378 63320
rect 79712 62626 79718 62714
rect 80322 62710 80336 62798
rect 79658 62516 79718 62626
rect 80370 62710 80378 62798
rect 80982 65402 80994 65512
rect 81634 65574 81710 65670
rect 81028 65402 81038 65512
rect 81634 65492 81652 65574
rect 80982 64880 81038 65402
rect 80982 64708 80994 64880
rect 81028 64708 81038 64880
rect 80982 64186 81038 64708
rect 80982 64014 80994 64186
rect 81028 64014 81038 64186
rect 80982 63492 81038 64014
rect 80982 63320 80994 63492
rect 81028 63320 81038 63492
rect 80982 62798 81038 63320
rect 80982 62668 80994 62798
rect 80336 62610 80370 62626
rect 80986 62626 80994 62668
rect 81028 62756 81038 62798
rect 81636 65402 81652 65492
rect 81686 65492 81710 65574
rect 81686 65402 81692 65492
rect 81636 64880 81692 65402
rect 81636 64708 81652 64880
rect 81686 64708 81692 64880
rect 81636 64186 81692 64708
rect 81636 64014 81652 64186
rect 81686 64014 81692 64186
rect 81636 63492 81692 64014
rect 81636 63320 81652 63492
rect 81686 63320 81692 63492
rect 81636 62798 81692 63320
rect 81028 62626 81046 62756
rect 81636 62672 81652 62798
rect 80986 62520 81046 62626
rect 81686 62672 81692 62798
rect 81652 62610 81686 62626
rect 80986 62516 81144 62520
rect 79658 62454 81144 62516
rect 79658 62448 79718 62454
rect 80986 62446 81046 62454
rect 81642 61966 81820 61976
rect 81634 61958 81820 61966
rect 79002 61916 81820 61958
rect 73314 61644 73324 61754
rect 73920 61734 73938 61816
rect 73268 61122 73324 61644
rect 73268 60950 73280 61122
rect 73314 60950 73324 61122
rect 73268 60428 73324 60950
rect 73268 60256 73280 60428
rect 73314 60256 73324 60428
rect 73268 59734 73324 60256
rect 73268 59562 73280 59734
rect 73314 59562 73324 59734
rect 73268 59040 73324 59562
rect 73268 58910 73280 59040
rect 72622 58852 72656 58868
rect 73272 58868 73280 58910
rect 73314 58998 73324 59040
rect 73922 61644 73938 61734
rect 73972 61734 73996 61816
rect 75156 61796 75212 61902
rect 74872 61736 75088 61796
rect 73972 61644 73978 61734
rect 73922 61122 73978 61644
rect 73922 60950 73938 61122
rect 73972 60950 73978 61122
rect 73922 60428 73978 60950
rect 73922 60256 73938 60428
rect 73972 60256 73978 60428
rect 73922 59734 73978 60256
rect 73922 59562 73938 59734
rect 73972 59562 73978 59734
rect 73922 59040 73978 59562
rect 73314 58868 73332 58998
rect 73922 58914 73938 59040
rect 73272 58762 73332 58868
rect 73972 58914 73978 59040
rect 74872 58990 74902 61736
rect 75042 58990 75088 61736
rect 75156 61624 75170 61796
rect 75204 61624 75212 61796
rect 75828 61796 75862 61812
rect 75156 61102 75212 61624
rect 75156 60930 75170 61102
rect 75204 60930 75212 61102
rect 75156 60408 75212 60930
rect 75156 60236 75170 60408
rect 75204 60236 75212 60408
rect 75156 59714 75212 60236
rect 75156 59542 75170 59714
rect 75204 59542 75212 59714
rect 75156 59136 75212 59542
rect 75818 61624 75828 61780
rect 76474 61796 76530 61902
rect 77784 61892 77970 61902
rect 75862 61624 75874 61780
rect 76474 61776 76486 61796
rect 75818 61102 75874 61624
rect 75818 60930 75828 61102
rect 75862 60930 75874 61102
rect 75818 60408 75874 60930
rect 75818 60236 75828 60408
rect 75862 60236 75874 60408
rect 75818 59714 75874 60236
rect 75818 59542 75828 59714
rect 75862 59542 75874 59714
rect 74872 58936 75088 58990
rect 75152 59020 75228 59136
rect 73938 58852 73972 58868
rect 75152 58848 75170 59020
rect 75204 58848 75228 59020
rect 75818 59020 75874 59542
rect 75818 58980 75828 59020
rect 73272 58758 73430 58762
rect 71944 58696 73430 58758
rect 71944 58690 72004 58696
rect 73272 58688 73332 58696
rect 73928 58196 74106 58206
rect 73920 58188 74106 58196
rect 71288 58146 74106 58188
rect 71288 58088 71364 58146
rect 71292 58040 71348 58088
rect 71008 57980 71224 58040
rect 57302 57732 57566 57746
rect 54540 57726 57566 57732
rect 54404 57692 54420 57726
rect 54592 57692 55114 57726
rect 55286 57692 55808 57726
rect 55980 57692 56502 57726
rect 56674 57692 57196 57726
rect 57368 57692 57566 57726
rect 54540 57678 57566 57692
rect 57302 57670 57566 57678
rect 57482 57668 57536 57670
rect 57190 57112 58092 57124
rect 42200 57086 42500 57098
rect 46194 57086 46494 57098
rect 50216 57086 50516 57098
rect 54238 57086 54538 57098
rect 57190 57086 58868 57112
rect 42200 57068 58868 57086
rect 42200 57034 42382 57068
rect 42554 57034 43076 57068
rect 43248 57034 43770 57068
rect 43942 57034 44464 57068
rect 44636 57034 45158 57068
rect 45330 57034 46376 57068
rect 46548 57034 47070 57068
rect 47242 57034 47764 57068
rect 47936 57034 48458 57068
rect 48630 57034 49152 57068
rect 49324 57034 50398 57068
rect 50570 57034 51092 57068
rect 51264 57034 51786 57068
rect 51958 57034 52480 57068
rect 52652 57034 53174 57068
rect 53346 57034 54420 57068
rect 54592 57034 55114 57068
rect 55286 57034 55808 57068
rect 55980 57034 56502 57068
rect 56674 57034 57196 57068
rect 57368 57034 58868 57068
rect 42200 57024 45342 57034
rect 46194 57024 49336 57034
rect 50216 57024 53358 57034
rect 54238 57024 58868 57034
rect 42200 57022 42482 57024
rect 46194 57022 46476 57024
rect 50216 57022 50498 57024
rect 54238 57022 54520 57024
rect 42204 57020 42286 57022
rect 46198 57020 46280 57022
rect 50220 57020 50302 57022
rect 54242 57020 54324 57022
rect 57190 56922 58868 57024
rect 57190 56896 58092 56922
rect 30322 56854 30416 56870
rect 30322 56832 30340 56854
rect 23482 56830 23760 56832
rect 30150 56830 30340 56832
rect 23482 56822 30340 56830
rect 23482 56788 23634 56822
rect 23806 56788 24328 56822
rect 24500 56788 25022 56822
rect 25194 56788 25716 56822
rect 25888 56788 26410 56822
rect 26582 56788 27104 56822
rect 27276 56788 27798 56822
rect 27970 56788 28492 56822
rect 28664 56788 29186 56822
rect 29358 56788 29880 56822
rect 30052 56790 30340 56822
rect 30052 56788 30230 56790
rect 23482 56768 30042 56788
rect 23482 56764 23760 56768
rect 19624 56720 20578 56722
rect 19528 56686 19544 56720
rect 19716 56686 20238 56720
rect 20410 56686 20578 56720
rect 19624 56668 20578 56686
rect 20334 56652 20578 56668
rect 19348 56062 20410 56076
rect 19348 56028 19544 56062
rect 19716 56028 20238 56062
rect 20410 56028 20426 56062
rect 19348 56018 20410 56028
rect 19348 55980 19630 56018
rect 18314 55368 18600 55370
rect 16916 55360 18600 55368
rect 16844 55326 16860 55360
rect 17032 55326 17554 55360
rect 17726 55326 18248 55360
rect 18420 55326 18600 55360
rect 16916 55316 18600 55326
rect 16548 54712 17034 54768
rect 16548 54702 18458 54712
rect 16548 54668 16860 54702
rect 17032 54668 17554 54702
rect 17726 54668 18248 54702
rect 18420 54668 18458 54702
rect 18532 54684 18600 55316
rect 16548 54660 18458 54668
rect 16548 54610 17034 54660
rect 18522 54642 18600 54684
rect 18522 54058 18596 54642
rect 19352 54844 19420 55980
rect 20478 55614 20560 56652
rect 30150 56180 30206 56788
rect 30322 56768 30340 56790
rect 30394 56768 30416 56854
rect 30322 56750 30416 56768
rect 29994 56176 30206 56180
rect 23706 56164 30206 56176
rect 23618 56130 23634 56164
rect 23806 56130 24328 56164
rect 24500 56130 25022 56164
rect 25194 56130 25716 56164
rect 25888 56130 26410 56164
rect 26582 56130 27104 56164
rect 27276 56130 27798 56164
rect 27970 56130 28492 56164
rect 28664 56130 29186 56164
rect 29358 56130 29880 56164
rect 30052 56130 30206 56164
rect 23706 56120 30206 56130
rect 42678 56472 45324 56508
rect 42678 56140 42828 56472
rect 45228 56140 45324 56472
rect 23706 56118 30202 56120
rect 23706 56114 30020 56118
rect 29406 55990 29534 56114
rect 42678 56106 45324 56140
rect 46686 56470 49332 56506
rect 46686 56138 46836 56470
rect 49236 56138 49332 56470
rect 46686 56104 49332 56138
rect 50698 56470 53344 56506
rect 50698 56138 50848 56470
rect 53248 56138 53344 56470
rect 50698 56104 53344 56138
rect 54708 56470 57354 56506
rect 54708 56138 54858 56470
rect 57258 56138 57354 56470
rect 54708 56104 57354 56138
rect 28686 55970 29576 55990
rect 45210 55984 45474 55998
rect 49218 55984 49482 55996
rect 53230 55984 53494 55996
rect 57240 55984 57504 55996
rect 24274 55868 25162 55908
rect 24274 55766 24368 55868
rect 25098 55766 25162 55868
rect 28686 55872 28714 55970
rect 29532 55872 29576 55970
rect 42392 55968 57504 55984
rect 42318 55934 42334 55968
rect 42506 55934 43028 55968
rect 43200 55934 43722 55968
rect 43894 55934 44416 55968
rect 44588 55934 45110 55968
rect 45282 55966 57504 55968
rect 45282 55934 46342 55966
rect 42392 55932 46342 55934
rect 46514 55932 47036 55966
rect 47208 55932 47730 55966
rect 47902 55932 48424 55966
rect 48596 55932 49118 55966
rect 49290 55932 50354 55966
rect 50526 55932 51048 55966
rect 51220 55932 51742 55966
rect 51914 55932 52436 55966
rect 52608 55932 53130 55966
rect 53302 55932 54364 55966
rect 54536 55932 55058 55966
rect 55230 55932 55752 55966
rect 55924 55932 56446 55966
rect 56618 55932 57140 55966
rect 57312 55932 57504 55966
rect 42408 55926 45474 55932
rect 45210 55922 45474 55926
rect 46416 55924 49482 55932
rect 50428 55924 53494 55932
rect 54438 55924 57504 55932
rect 28686 55848 29576 55872
rect 24274 55732 25162 55766
rect 20464 55596 23774 55614
rect 30154 55598 30214 55652
rect 30028 55596 30214 55598
rect 20464 55590 30214 55596
rect 20464 55556 23640 55590
rect 23812 55556 24334 55590
rect 24506 55556 25028 55590
rect 25200 55556 25722 55590
rect 25894 55556 26416 55590
rect 26588 55556 27110 55590
rect 27282 55556 27804 55590
rect 27976 55556 28498 55590
rect 28670 55556 29192 55590
rect 29364 55556 29886 55590
rect 30058 55556 30214 55590
rect 20464 55542 30214 55556
rect 20464 55534 30046 55542
rect 20464 55532 23774 55534
rect 20478 55418 20560 55532
rect 20316 55406 20560 55418
rect 19608 55404 20560 55406
rect 19528 55370 19544 55404
rect 19716 55370 20238 55404
rect 20410 55370 20560 55404
rect 19608 55348 20560 55370
rect 19054 54766 19420 54844
rect 19054 54756 19634 54766
rect 19054 54746 20394 54756
rect 19054 54712 19544 54746
rect 19716 54712 20238 54746
rect 20410 54712 20426 54746
rect 19054 54698 20394 54712
rect 19054 54676 19634 54698
rect 19352 54670 19634 54676
rect 20478 54112 20560 55348
rect 22916 55346 23202 55376
rect 22916 54924 22980 55346
rect 23102 55070 23202 55346
rect 23102 54974 23484 55070
rect 23102 54942 23538 54974
rect 23102 54940 23766 54942
rect 23102 54932 30048 54940
rect 23102 54924 23640 54932
rect 22916 54898 23640 54924
rect 23812 54898 24334 54932
rect 24506 54898 25028 54932
rect 25200 54898 25722 54932
rect 25894 54898 26416 54932
rect 26588 54898 27110 54932
rect 27282 54898 27804 54932
rect 27976 54898 28498 54932
rect 28670 54898 29192 54932
rect 29364 54898 29886 54932
rect 30058 54898 30074 54932
rect 22916 54892 30048 54898
rect 22916 54860 23202 54892
rect 23316 54878 30048 54892
rect 23316 54874 23766 54878
rect 23316 54844 23538 54874
rect 23278 54734 23414 54780
rect 20658 54660 20824 54672
rect 20658 54424 20678 54660
rect 20792 54424 20824 54660
rect 20658 54392 20824 54424
rect 23278 54418 23294 54734
rect 23382 54418 23414 54734
rect 23278 54366 23414 54418
rect 30156 54290 30212 55542
rect 30000 54286 30212 54290
rect 23712 54274 30212 54286
rect 23624 54240 23640 54274
rect 23812 54240 24334 54274
rect 24506 54240 25028 54274
rect 25200 54240 25722 54274
rect 25894 54240 26416 54274
rect 26588 54240 27110 54274
rect 27282 54240 27804 54274
rect 27976 54240 28498 54274
rect 28670 54240 29192 54274
rect 29364 54240 29886 54274
rect 30058 54240 30212 54274
rect 23712 54230 30212 54240
rect 42156 55322 42442 55336
rect 42156 55310 45292 55322
rect 42156 55276 42334 55310
rect 42506 55276 43028 55310
rect 43200 55276 43722 55310
rect 43894 55276 44416 55310
rect 44588 55276 45110 55310
rect 45282 55276 45298 55310
rect 42156 55268 45292 55276
rect 42156 55260 42442 55268
rect 23712 54228 30208 54230
rect 23712 54224 30026 54228
rect 20316 54100 20560 54112
rect 19592 54088 20560 54100
rect 15752 54048 15974 54054
rect 18378 54052 18600 54058
rect 19528 54054 19544 54088
rect 19716 54054 20238 54088
rect 20410 54054 20560 54088
rect 1030 54038 2678 54046
rect 5124 54042 5346 54048
rect 922 54004 938 54038
rect 1110 54004 1632 54038
rect 1804 54004 2326 54038
rect 2498 54004 2678 54038
rect 3698 54034 5346 54042
rect 6372 54040 8020 54048
rect 9018 54040 10666 54048
rect 13098 54042 13320 54048
rect 1030 53994 2678 54004
rect 3590 54000 3606 54034
rect 3778 54000 4300 54034
rect 4472 54000 4994 54034
rect 5166 54000 5346 54034
rect 6264 54006 6280 54040
rect 6452 54006 6974 54040
rect 7146 54006 7668 54040
rect 7840 54006 8020 54040
rect 8910 54006 8926 54040
rect 9098 54006 9620 54040
rect 9792 54006 10314 54040
rect 10486 54006 10666 54040
rect 11672 54034 13320 54042
rect 14326 54040 15974 54048
rect 16952 54044 18600 54052
rect 2456 53982 2678 53994
rect 3698 53990 5346 54000
rect 6372 53996 8020 54006
rect 9018 53996 10666 54006
rect 11564 54000 11580 54034
rect 11752 54000 12274 54034
rect 12446 54000 12968 54034
rect 13140 54000 13320 54034
rect 14218 54006 14234 54040
rect 14406 54006 14928 54040
rect 15100 54006 15622 54040
rect 15794 54006 15974 54040
rect 16844 54010 16860 54044
rect 17032 54010 17554 54044
rect 17726 54010 18248 54044
rect 18420 54010 18600 54044
rect 19592 54042 20560 54054
rect 20478 54036 20560 54042
rect 28692 54094 29582 54100
rect 28692 54080 29852 54094
rect 5124 53978 5346 53990
rect 7798 53984 8020 53996
rect 10444 53984 10666 53996
rect 11672 53990 13320 54000
rect 14326 53996 15974 54006
rect 16952 54000 18600 54010
rect 13098 53978 13320 53990
rect 15752 53984 15974 53996
rect 18378 53988 18600 54000
rect 24280 53978 25168 54018
rect 24280 53876 24374 53978
rect 25104 53876 25168 53978
rect 28692 53982 28720 54080
rect 29538 53982 29852 54080
rect 42156 54014 42238 55260
rect 45396 54670 45450 55922
rect 49218 55920 49482 55924
rect 53230 55920 53494 55924
rect 57240 55920 57504 55924
rect 46164 55320 46450 55334
rect 46164 55308 49300 55320
rect 46164 55274 46342 55308
rect 46514 55274 47036 55308
rect 47208 55274 47730 55308
rect 47902 55274 48424 55308
rect 48596 55274 49118 55308
rect 49290 55274 49306 55308
rect 46164 55266 49300 55274
rect 46164 55258 46450 55266
rect 45246 54664 45510 54670
rect 42456 54652 45510 54664
rect 42318 54618 42334 54652
rect 42506 54618 43028 54652
rect 43200 54618 43722 54652
rect 43894 54618 44416 54652
rect 44588 54618 45110 54652
rect 45282 54618 45510 54652
rect 42456 54610 45510 54618
rect 45246 54594 45510 54610
rect 28692 53978 29852 53982
rect 42152 54006 42472 54014
rect 42152 53994 45300 54006
rect 28692 53958 29582 53978
rect 42152 53960 42334 53994
rect 42506 53960 43028 53994
rect 43200 53960 43722 53994
rect 43894 53960 44416 53994
rect 44588 53960 45110 53994
rect 45282 53960 45300 53994
rect 42152 53952 45300 53960
rect 42152 53938 42472 53952
rect 24280 53842 25168 53876
rect 30172 53656 30228 53660
rect 30044 53654 30230 53656
rect 23748 53648 30230 53654
rect 23640 53614 23656 53648
rect 23828 53614 24350 53648
rect 24522 53614 25044 53648
rect 25216 53614 25738 53648
rect 25910 53614 26432 53648
rect 26604 53614 27126 53648
rect 27298 53614 27820 53648
rect 27992 53614 28514 53648
rect 28686 53614 29208 53648
rect 29380 53614 29902 53648
rect 30074 53614 30230 53648
rect 23748 53600 30230 53614
rect 23748 53592 30062 53600
rect 19364 53336 20600 53360
rect 944 53294 2576 53328
rect 944 53152 1000 53294
rect 2514 53152 2576 53294
rect 944 53124 2576 53152
rect 3612 53290 5244 53324
rect 3612 53148 3668 53290
rect 5182 53148 5244 53290
rect 3612 53120 5244 53148
rect 6286 53296 7918 53330
rect 6286 53154 6342 53296
rect 7856 53154 7918 53296
rect 6286 53126 7918 53154
rect 8932 53296 10564 53330
rect 8932 53154 8988 53296
rect 10502 53154 10564 53296
rect 8932 53126 10564 53154
rect 11586 53290 13218 53324
rect 11586 53148 11642 53290
rect 13156 53148 13218 53290
rect 11586 53120 13218 53148
rect 14240 53296 15872 53330
rect 14240 53154 14296 53296
rect 15810 53154 15872 53296
rect 14240 53126 15872 53154
rect 16866 53300 18498 53334
rect 16866 53158 16922 53300
rect 18436 53158 18498 53300
rect 16866 53130 18498 53158
rect 19364 53142 19472 53336
rect 20538 53142 20600 53336
rect 19364 53090 20600 53142
rect 2360 53006 20528 53048
rect 2360 52998 20552 53006
rect 30172 53002 30228 53600
rect 30360 53076 30510 53106
rect 30360 53002 30374 53076
rect 23504 52998 23782 53000
rect 30034 52998 30374 53002
rect 2360 52986 20560 52998
rect 2360 52954 19544 52986
rect 908 52952 19544 52954
rect 19716 52952 20238 52986
rect 20410 52952 20560 52986
rect 908 52942 20560 52952
rect 908 52938 16860 52942
rect 908 52936 6280 52938
rect 908 52902 938 52936
rect 1110 52902 1632 52936
rect 1804 52902 2326 52936
rect 2498 52932 6280 52936
rect 2498 52902 3606 52932
rect 908 52898 3606 52902
rect 3778 52898 4300 52932
rect 4472 52898 4994 52932
rect 5166 52904 6280 52932
rect 6452 52904 6974 52938
rect 7146 52904 7668 52938
rect 7840 52904 8926 52938
rect 9098 52904 9620 52938
rect 9792 52904 10314 52938
rect 10486 52932 14234 52938
rect 10486 52904 11580 52932
rect 5166 52898 11580 52904
rect 11752 52898 12274 52932
rect 12446 52898 12968 52932
rect 13140 52904 14234 52932
rect 14406 52904 14928 52938
rect 15100 52904 15622 52938
rect 15794 52908 16860 52938
rect 17032 52908 17554 52942
rect 17726 52908 18248 52942
rect 18420 52908 20560 52942
rect 23504 52990 30374 52998
rect 23504 52956 23656 52990
rect 23828 52956 24350 52990
rect 24522 52956 25044 52990
rect 25216 52956 25738 52990
rect 25910 52956 26432 52990
rect 26604 52956 27126 52990
rect 27298 52956 27820 52990
rect 27992 52956 28514 52990
rect 28686 52956 29208 52990
rect 29380 52956 29902 52990
rect 30074 52956 30374 52990
rect 23504 52940 30374 52956
rect 23504 52936 30064 52940
rect 23504 52932 23782 52936
rect 15794 52904 20560 52908
rect 13140 52898 20560 52904
rect 908 52890 20560 52898
rect 2360 52878 20560 52890
rect 746 52290 1066 52312
rect 746 52288 2474 52290
rect 728 52278 2474 52288
rect 728 52244 938 52278
rect 1110 52244 1632 52278
rect 1804 52244 2326 52278
rect 2498 52244 2514 52278
rect 728 52238 2474 52244
rect 728 52190 1066 52238
rect 728 50990 820 52190
rect 2610 51628 2678 52878
rect 3414 52286 3734 52308
rect 3414 52284 5142 52286
rect 956 51620 2678 51628
rect 922 51586 938 51620
rect 1110 51586 1632 51620
rect 1804 51586 2326 51620
rect 2498 51586 2678 51620
rect 956 51576 2678 51586
rect 2390 51574 2678 51576
rect 728 50968 1052 50990
rect 728 50962 2478 50968
rect 728 50928 938 50962
rect 1110 50928 1632 50962
rect 1804 50928 2326 50962
rect 2498 50928 2514 50962
rect 728 50916 2478 50928
rect 728 50868 1052 50916
rect 728 49676 820 50868
rect 2610 50316 2678 51574
rect 2402 50314 2678 50316
rect 970 50304 2678 50314
rect 922 50270 938 50304
rect 1110 50270 1632 50304
rect 1804 50270 2326 50304
rect 2498 50270 2678 50304
rect 970 50262 2678 50270
rect 722 49654 1042 49676
rect 722 49646 2488 49654
rect 722 49612 938 49646
rect 1110 49612 1632 49646
rect 1804 49612 2326 49646
rect 2498 49612 2514 49646
rect 722 49602 2488 49612
rect 722 49554 1042 49602
rect 728 48388 820 49554
rect 2610 48998 2678 50262
rect 3396 52274 5142 52284
rect 3396 52240 3606 52274
rect 3778 52240 4300 52274
rect 4472 52240 4994 52274
rect 5166 52240 5182 52274
rect 3396 52234 5142 52240
rect 3396 52186 3734 52234
rect 3396 50986 3488 52186
rect 5278 51624 5346 52878
rect 6088 52292 6408 52314
rect 6088 52290 7816 52292
rect 3624 51616 5346 51624
rect 3590 51582 3606 51616
rect 3778 51582 4300 51616
rect 4472 51582 4994 51616
rect 5166 51582 5346 51616
rect 3624 51572 5346 51582
rect 5058 51570 5346 51572
rect 3396 50964 3720 50986
rect 3396 50958 5146 50964
rect 3396 50924 3606 50958
rect 3778 50924 4300 50958
rect 4472 50924 4994 50958
rect 5166 50924 5182 50958
rect 3396 50912 5146 50924
rect 3396 50864 3720 50912
rect 3396 49672 3488 50864
rect 5278 50312 5346 51570
rect 5070 50310 5346 50312
rect 3638 50300 5346 50310
rect 3590 50266 3606 50300
rect 3778 50266 4300 50300
rect 4472 50266 4994 50300
rect 5166 50266 5346 50300
rect 3638 50258 5346 50266
rect 3390 49650 3710 49672
rect 3390 49642 5156 49650
rect 3390 49608 3606 49642
rect 3778 49608 4300 49642
rect 4472 49608 4994 49642
rect 5166 49608 5182 49642
rect 3390 49598 5156 49608
rect 3390 49550 3710 49598
rect 2392 48996 2678 48998
rect 994 48988 2678 48996
rect 922 48954 938 48988
rect 1110 48954 1632 48988
rect 1804 48954 2326 48988
rect 2498 48954 2678 48988
rect 994 48944 2678 48954
rect 712 48340 1032 48388
rect 712 48330 2536 48340
rect 712 48296 938 48330
rect 1110 48296 1632 48330
rect 1804 48296 2326 48330
rect 2498 48296 2536 48330
rect 2610 48312 2678 48944
rect 712 48288 2536 48296
rect 712 48266 1032 48288
rect 2600 48270 2678 48312
rect 2600 47686 2674 48270
rect 3396 48384 3488 49550
rect 5278 48994 5346 50258
rect 6070 52280 7816 52290
rect 6070 52246 6280 52280
rect 6452 52246 6974 52280
rect 7146 52246 7668 52280
rect 7840 52246 7856 52280
rect 6070 52240 7816 52246
rect 6070 52192 6408 52240
rect 6070 50992 6162 52192
rect 7952 51630 8020 52878
rect 8734 52292 9054 52314
rect 8734 52290 10462 52292
rect 6298 51622 8020 51630
rect 6264 51588 6280 51622
rect 6452 51588 6974 51622
rect 7146 51588 7668 51622
rect 7840 51588 8020 51622
rect 6298 51578 8020 51588
rect 7732 51576 8020 51578
rect 6070 50970 6394 50992
rect 6070 50964 7820 50970
rect 6070 50930 6280 50964
rect 6452 50930 6974 50964
rect 7146 50930 7668 50964
rect 7840 50930 7856 50964
rect 6070 50918 7820 50930
rect 6070 50870 6394 50918
rect 6070 49678 6162 50870
rect 7952 50318 8020 51576
rect 7744 50316 8020 50318
rect 6312 50306 8020 50316
rect 6264 50272 6280 50306
rect 6452 50272 6974 50306
rect 7146 50272 7668 50306
rect 7840 50272 8020 50306
rect 6312 50264 8020 50272
rect 6064 49656 6384 49678
rect 6064 49648 7830 49656
rect 6064 49614 6280 49648
rect 6452 49614 6974 49648
rect 7146 49614 7668 49648
rect 7840 49614 7856 49648
rect 6064 49604 7830 49614
rect 6064 49556 6384 49604
rect 5060 48992 5346 48994
rect 3662 48984 5346 48992
rect 3590 48950 3606 48984
rect 3778 48950 4300 48984
rect 4472 48950 4994 48984
rect 5166 48950 5346 48984
rect 3662 48940 5346 48950
rect 3380 48376 3700 48384
rect 3276 48336 3700 48376
rect 3276 48326 5204 48336
rect 3276 48292 3606 48326
rect 3778 48292 4300 48326
rect 4472 48292 4994 48326
rect 5166 48292 5204 48326
rect 5278 48308 5346 48940
rect 3276 48284 5204 48292
rect 3276 48262 3700 48284
rect 5268 48266 5346 48308
rect 3276 48234 3504 48262
rect 2456 47680 2678 47686
rect 5268 47682 5342 48266
rect 6070 48390 6162 49556
rect 7952 49000 8020 50264
rect 8716 52280 10462 52290
rect 8716 52246 8926 52280
rect 9098 52246 9620 52280
rect 9792 52246 10314 52280
rect 10486 52246 10502 52280
rect 8716 52240 10462 52246
rect 8716 52192 9054 52240
rect 8716 50992 8808 52192
rect 10598 51630 10666 52878
rect 11388 52286 11708 52308
rect 11388 52284 13116 52286
rect 8944 51622 10666 51630
rect 8910 51588 8926 51622
rect 9098 51588 9620 51622
rect 9792 51588 10314 51622
rect 10486 51588 10666 51622
rect 8944 51578 10666 51588
rect 10378 51576 10666 51578
rect 8716 50970 9040 50992
rect 8716 50964 10466 50970
rect 8716 50930 8926 50964
rect 9098 50930 9620 50964
rect 9792 50930 10314 50964
rect 10486 50930 10502 50964
rect 8716 50918 10466 50930
rect 8716 50870 9040 50918
rect 8716 49678 8808 50870
rect 10598 50318 10666 51576
rect 10390 50316 10666 50318
rect 8958 50306 10666 50316
rect 8910 50272 8926 50306
rect 9098 50272 9620 50306
rect 9792 50272 10314 50306
rect 10486 50272 10666 50306
rect 8958 50264 10666 50272
rect 8710 49656 9030 49678
rect 8710 49648 10476 49656
rect 8710 49614 8926 49648
rect 9098 49614 9620 49648
rect 9792 49614 10314 49648
rect 10486 49614 10502 49648
rect 8710 49604 10476 49614
rect 8710 49556 9030 49604
rect 7734 48998 8020 49000
rect 6336 48990 8020 48998
rect 6264 48956 6280 48990
rect 6452 48956 6974 48990
rect 7146 48956 7668 48990
rect 7840 48956 8020 48990
rect 6336 48946 8020 48956
rect 6054 48386 6374 48390
rect 5928 48342 6374 48386
rect 5928 48332 7878 48342
rect 5928 48298 6280 48332
rect 6452 48298 6974 48332
rect 7146 48298 7668 48332
rect 7840 48298 7878 48332
rect 7952 48314 8020 48946
rect 5928 48290 7878 48298
rect 5928 48276 6374 48290
rect 6054 48268 6374 48276
rect 7942 48272 8020 48314
rect 7942 47688 8016 48272
rect 8716 48402 8808 49556
rect 10598 49000 10666 50264
rect 11370 52274 13116 52284
rect 11370 52240 11580 52274
rect 11752 52240 12274 52274
rect 12446 52240 12968 52274
rect 13140 52240 13156 52274
rect 11370 52234 13116 52240
rect 11370 52186 11708 52234
rect 11370 50986 11462 52186
rect 13252 51624 13320 52878
rect 14042 52292 14362 52314
rect 14042 52290 15770 52292
rect 11598 51616 13320 51624
rect 11564 51582 11580 51616
rect 11752 51582 12274 51616
rect 12446 51582 12968 51616
rect 13140 51582 13320 51616
rect 11598 51572 13320 51582
rect 13032 51570 13320 51572
rect 11370 50964 11694 50986
rect 11370 50958 13120 50964
rect 11370 50924 11580 50958
rect 11752 50924 12274 50958
rect 12446 50924 12968 50958
rect 13140 50924 13156 50958
rect 11370 50912 13120 50924
rect 11370 50864 11694 50912
rect 11370 49672 11462 50864
rect 13252 50312 13320 51570
rect 13044 50310 13320 50312
rect 11612 50300 13320 50310
rect 11564 50266 11580 50300
rect 11752 50266 12274 50300
rect 12446 50266 12968 50300
rect 13140 50266 13320 50300
rect 11612 50258 13320 50266
rect 11364 49650 11684 49672
rect 11364 49642 13130 49650
rect 11364 49608 11580 49642
rect 11752 49608 12274 49642
rect 12446 49608 12968 49642
rect 13140 49608 13156 49642
rect 11364 49598 13130 49608
rect 11364 49550 11684 49598
rect 10380 48998 10666 49000
rect 8982 48990 10666 48998
rect 8910 48956 8926 48990
rect 9098 48956 9620 48990
rect 9792 48956 10314 48990
rect 10486 48956 10666 48990
rect 8982 48946 10666 48956
rect 8554 48390 8822 48402
rect 8554 48342 9020 48390
rect 8554 48332 10524 48342
rect 8554 48298 8926 48332
rect 9098 48298 9620 48332
rect 9792 48298 10314 48332
rect 10486 48298 10524 48332
rect 10598 48314 10666 48946
rect 8554 48290 10524 48298
rect 8554 48276 9020 48290
rect 8700 48268 9020 48276
rect 10588 48272 10666 48314
rect 10588 47688 10662 48272
rect 11370 48394 11462 49550
rect 13252 48994 13320 50258
rect 14024 52280 15770 52290
rect 14024 52246 14234 52280
rect 14406 52246 14928 52280
rect 15100 52246 15622 52280
rect 15794 52246 15810 52280
rect 14024 52240 15770 52246
rect 14024 52192 14362 52240
rect 14024 50992 14116 52192
rect 15906 51630 15974 52878
rect 16668 52296 16988 52318
rect 16668 52294 18396 52296
rect 14252 51622 15974 51630
rect 14218 51588 14234 51622
rect 14406 51588 14928 51622
rect 15100 51588 15622 51622
rect 15794 51588 15974 51622
rect 14252 51578 15974 51588
rect 15686 51576 15974 51578
rect 14024 50970 14348 50992
rect 14024 50964 15774 50970
rect 14024 50930 14234 50964
rect 14406 50930 14928 50964
rect 15100 50930 15622 50964
rect 15794 50930 15810 50964
rect 14024 50918 15774 50930
rect 14024 50870 14348 50918
rect 14024 49678 14116 50870
rect 15906 50318 15974 51576
rect 15698 50316 15974 50318
rect 14266 50306 15974 50316
rect 14218 50272 14234 50306
rect 14406 50272 14928 50306
rect 15100 50272 15622 50306
rect 15794 50272 15974 50306
rect 14266 50264 15974 50272
rect 14018 49656 14338 49678
rect 14018 49648 15784 49656
rect 14018 49614 14234 49648
rect 14406 49614 14928 49648
rect 15100 49614 15622 49648
rect 15794 49614 15810 49648
rect 14018 49604 15784 49614
rect 14018 49556 14338 49604
rect 13034 48992 13320 48994
rect 11636 48984 13320 48992
rect 11564 48950 11580 48984
rect 11752 48950 12274 48984
rect 12446 48950 12968 48984
rect 13140 48950 13320 48984
rect 11636 48940 13320 48950
rect 11246 48336 11920 48394
rect 11246 48326 13178 48336
rect 11246 48292 11580 48326
rect 11752 48292 12274 48326
rect 12446 48292 12968 48326
rect 13140 48292 13178 48326
rect 13252 48308 13320 48940
rect 11246 48284 13178 48292
rect 11246 48276 11920 48284
rect 11354 48262 11674 48276
rect 13242 48266 13320 48308
rect 7798 47682 8020 47688
rect 10444 47682 10666 47688
rect 13242 47682 13316 48266
rect 14024 48390 14116 49556
rect 15906 49000 15974 50264
rect 16650 52284 18396 52294
rect 16650 52250 16860 52284
rect 17032 52250 17554 52284
rect 17726 52250 18248 52284
rect 18420 52250 18436 52284
rect 16650 52244 18396 52250
rect 16650 52196 16988 52244
rect 16650 50996 16742 52196
rect 18532 51634 18600 52878
rect 19336 52344 19618 52354
rect 19336 52328 20414 52344
rect 19336 52294 19544 52328
rect 19716 52294 20238 52328
rect 20410 52294 20426 52328
rect 19336 52286 20414 52294
rect 19336 52258 19618 52286
rect 16878 51626 18600 51634
rect 16844 51592 16860 51626
rect 17032 51592 17554 51626
rect 17726 51592 18248 51626
rect 18420 51592 18600 51626
rect 16878 51582 18600 51592
rect 18312 51580 18600 51582
rect 16650 50974 16974 50996
rect 16650 50968 18400 50974
rect 16650 50934 16860 50968
rect 17032 50934 17554 50968
rect 17726 50934 18248 50968
rect 18420 50934 18436 50968
rect 16650 50922 18400 50934
rect 16650 50874 16974 50922
rect 16650 49682 16742 50874
rect 18532 50322 18600 51580
rect 18324 50320 18600 50322
rect 16892 50310 18600 50320
rect 16844 50276 16860 50310
rect 17032 50276 17554 50310
rect 17726 50276 18248 50310
rect 18420 50276 18600 50310
rect 16892 50268 18600 50276
rect 16644 49660 16964 49682
rect 16644 49652 18410 49660
rect 16644 49618 16860 49652
rect 17032 49618 17554 49652
rect 17726 49618 18248 49652
rect 18420 49618 18436 49652
rect 16644 49608 18410 49618
rect 16644 49560 16964 49608
rect 15688 48998 15974 49000
rect 14290 48990 15974 48998
rect 14218 48956 14234 48990
rect 14406 48956 14928 48990
rect 15100 48956 15622 48990
rect 15794 48956 15974 48990
rect 14290 48946 15974 48956
rect 14008 48368 14328 48390
rect 13846 48342 14460 48368
rect 13846 48332 15832 48342
rect 13846 48298 14234 48332
rect 14406 48298 14928 48332
rect 15100 48298 15622 48332
rect 15794 48298 15832 48332
rect 15906 48314 15974 48946
rect 13846 48290 15832 48298
rect 13846 48250 14460 48290
rect 15896 48272 15974 48314
rect 15896 47688 15970 48272
rect 16650 48402 16742 49560
rect 18532 49004 18600 50268
rect 19352 51038 19420 52258
rect 19612 51674 20414 51680
rect 20478 51674 20560 52878
rect 30172 52348 30228 52940
rect 30360 52928 30374 52940
rect 30470 52928 30510 53076
rect 30360 52892 30510 52928
rect 42156 52714 42238 53938
rect 45396 53356 45450 54594
rect 46164 54012 46246 55258
rect 49404 54668 49458 55920
rect 50176 55320 50462 55334
rect 50176 55308 53312 55320
rect 50176 55274 50354 55308
rect 50526 55274 51048 55308
rect 51220 55274 51742 55308
rect 51914 55274 52436 55308
rect 52608 55274 53130 55308
rect 53302 55274 53318 55308
rect 50176 55266 53312 55274
rect 50176 55258 50462 55266
rect 49254 54662 49518 54668
rect 46464 54650 49518 54662
rect 46326 54616 46342 54650
rect 46514 54616 47036 54650
rect 47208 54616 47730 54650
rect 47902 54616 48424 54650
rect 48596 54616 49118 54650
rect 49290 54616 49518 54650
rect 46464 54608 49518 54616
rect 49254 54592 49518 54608
rect 46160 54004 46480 54012
rect 46160 53992 49308 54004
rect 46160 53958 46342 53992
rect 46514 53958 47036 53992
rect 47208 53958 47730 53992
rect 47902 53958 48424 53992
rect 48596 53958 49118 53992
rect 49290 53958 49308 53992
rect 46160 53950 49308 53958
rect 46160 53936 46480 53950
rect 45216 53342 45480 53356
rect 42454 53336 45480 53342
rect 42318 53302 42334 53336
rect 42506 53302 43028 53336
rect 43200 53302 43722 53336
rect 43894 53302 44416 53336
rect 44588 53302 45110 53336
rect 45282 53302 45480 53336
rect 42454 53288 45480 53302
rect 45216 53280 45480 53288
rect 45396 53278 45450 53280
rect 29484 52344 29558 52346
rect 30016 52344 30228 52348
rect 23728 52332 30228 52344
rect 23640 52298 23656 52332
rect 23828 52298 24350 52332
rect 24522 52298 25044 52332
rect 25216 52298 25738 52332
rect 25910 52298 26432 52332
rect 26604 52298 27126 52332
rect 27298 52298 27820 52332
rect 27992 52298 28514 52332
rect 28686 52298 29208 52332
rect 29380 52298 29902 52332
rect 30074 52298 30228 52332
rect 23728 52288 30228 52298
rect 42138 52708 42238 52714
rect 42138 52698 42452 52708
rect 46164 52706 46246 53936
rect 49404 53354 49458 54592
rect 50176 54012 50258 55258
rect 53416 54668 53470 55920
rect 54186 55320 54472 55334
rect 54186 55308 57322 55320
rect 54186 55274 54364 55308
rect 54536 55274 55058 55308
rect 55230 55274 55752 55308
rect 55924 55274 56446 55308
rect 56618 55274 57140 55308
rect 57312 55274 57328 55308
rect 54186 55266 57322 55274
rect 54186 55258 54472 55266
rect 53266 54662 53530 54668
rect 50476 54650 53530 54662
rect 50338 54616 50354 54650
rect 50526 54616 51048 54650
rect 51220 54616 51742 54650
rect 51914 54616 52436 54650
rect 52608 54616 53130 54650
rect 53302 54616 53530 54650
rect 50476 54608 53530 54616
rect 53266 54592 53530 54608
rect 50172 54004 50492 54012
rect 50172 53992 53320 54004
rect 50172 53958 50354 53992
rect 50526 53958 51048 53992
rect 51220 53958 51742 53992
rect 51914 53958 52436 53992
rect 52608 53958 53130 53992
rect 53302 53958 53320 53992
rect 50172 53950 53320 53958
rect 50172 53936 50492 53950
rect 49224 53340 49488 53354
rect 46462 53334 49488 53340
rect 46326 53300 46342 53334
rect 46514 53300 47036 53334
rect 47208 53300 47730 53334
rect 47902 53300 48424 53334
rect 48596 53300 49118 53334
rect 49290 53300 49488 53334
rect 46462 53286 49488 53300
rect 49224 53278 49488 53286
rect 49404 53276 49458 53278
rect 50176 52706 50258 53936
rect 53416 53354 53470 54592
rect 54186 54012 54268 55258
rect 57426 54668 57480 55920
rect 57276 54662 57540 54668
rect 54486 54650 57540 54662
rect 54348 54616 54364 54650
rect 54536 54616 55058 54650
rect 55230 54616 55752 54650
rect 55924 54616 56446 54650
rect 56618 54616 57140 54650
rect 57312 54616 57540 54650
rect 54486 54608 57540 54616
rect 57276 54592 57540 54608
rect 54182 54004 54502 54012
rect 54182 53992 57330 54004
rect 54182 53958 54364 53992
rect 54536 53958 55058 53992
rect 55230 53958 55752 53992
rect 55924 53958 56446 53992
rect 56618 53958 57140 53992
rect 57312 53958 57330 53992
rect 54182 53950 57330 53958
rect 54182 53936 54502 53950
rect 53236 53340 53500 53354
rect 50474 53334 53500 53340
rect 50338 53300 50354 53334
rect 50526 53300 51048 53334
rect 51220 53300 51742 53334
rect 51914 53300 52436 53334
rect 52608 53300 53130 53334
rect 53302 53300 53500 53334
rect 50474 53286 53500 53300
rect 53236 53278 53500 53286
rect 53416 53276 53470 53278
rect 54186 52706 54268 53936
rect 57426 53354 57480 54592
rect 57246 53340 57510 53354
rect 54484 53334 57510 53340
rect 54348 53300 54364 53334
rect 54536 53300 55058 53334
rect 55230 53300 55752 53334
rect 55924 53300 56446 53334
rect 56618 53300 57140 53334
rect 57312 53300 57510 53334
rect 54484 53286 57510 53300
rect 57246 53278 57510 53286
rect 46160 52698 46460 52706
rect 50172 52698 50472 52706
rect 54182 52698 54482 52706
rect 42138 52686 57198 52698
rect 42138 52678 57324 52686
rect 42138 52644 42334 52678
rect 42506 52644 43028 52678
rect 43200 52644 43722 52678
rect 43894 52644 44416 52678
rect 44588 52644 45110 52678
rect 45282 52676 57324 52678
rect 45282 52646 46342 52676
rect 45282 52644 45298 52646
rect 42138 52634 45294 52644
rect 46160 52642 46342 52646
rect 46514 52642 47036 52676
rect 47208 52642 47730 52676
rect 47902 52642 48424 52676
rect 48596 52642 49118 52676
rect 49290 52646 50354 52676
rect 49290 52642 49306 52646
rect 50172 52642 50354 52646
rect 50526 52642 51048 52676
rect 51220 52642 51742 52676
rect 51914 52642 52436 52676
rect 52608 52642 53130 52676
rect 53302 52646 54364 52676
rect 53302 52642 53318 52646
rect 54182 52642 54364 52646
rect 54536 52642 55058 52676
rect 55230 52642 55752 52676
rect 55924 52642 56446 52676
rect 56618 52642 57140 52676
rect 57312 52642 57328 52676
rect 42138 52632 42434 52634
rect 46160 52632 49302 52642
rect 50172 52632 53314 52642
rect 54182 52632 57324 52642
rect 42138 52630 42238 52632
rect 46160 52630 46442 52632
rect 50172 52630 50454 52632
rect 54182 52630 54464 52632
rect 23728 52286 30224 52288
rect 23728 52282 30042 52286
rect 29484 52158 29558 52282
rect 28708 52138 29598 52158
rect 24296 52036 25184 52076
rect 24296 51934 24390 52036
rect 25120 51934 25184 52036
rect 28708 52040 28736 52138
rect 29554 52040 29598 52138
rect 28708 52016 29598 52040
rect 24296 51900 25184 51934
rect 19612 51670 20560 51674
rect 19528 51636 19544 51670
rect 19716 51636 20238 51670
rect 20410 51636 20560 51670
rect 19612 51622 20560 51636
rect 20304 51604 20560 51622
rect 19352 51028 19638 51038
rect 19352 51012 20422 51028
rect 19352 50978 19544 51012
rect 19716 50978 20238 51012
rect 20410 50978 20426 51012
rect 19352 50970 20422 50978
rect 19352 50942 19638 50970
rect 19352 49710 19420 50942
rect 19624 50356 20426 50360
rect 20478 50356 20560 51604
rect 19624 50354 20578 50356
rect 19528 50320 19544 50354
rect 19716 50320 20238 50354
rect 20410 50320 20578 50354
rect 19624 50302 20578 50320
rect 20334 50286 20578 50302
rect 19348 49696 20410 49710
rect 19348 49662 19544 49696
rect 19716 49662 20238 49696
rect 20410 49662 20426 49696
rect 19348 49652 20410 49662
rect 19348 49614 19630 49652
rect 18314 49002 18600 49004
rect 16916 48994 18600 49002
rect 16844 48960 16860 48994
rect 17032 48960 17554 48994
rect 17726 48960 18248 48994
rect 18420 48960 18600 48994
rect 16916 48950 18600 48960
rect 16548 48346 17034 48402
rect 16548 48336 18458 48346
rect 16548 48302 16860 48336
rect 17032 48302 17554 48336
rect 17726 48302 18248 48336
rect 18420 48302 18458 48336
rect 18532 48318 18600 48950
rect 16548 48294 18458 48302
rect 16548 48244 17034 48294
rect 18522 48276 18600 48318
rect 18522 47692 18596 48276
rect 19352 48478 19420 49614
rect 20478 49052 20560 50286
rect 20316 49040 20560 49052
rect 19608 49038 20560 49040
rect 19528 49004 19544 49038
rect 19716 49004 20238 49038
rect 20410 49004 20560 49038
rect 19608 48982 20560 49004
rect 19054 48400 19420 48478
rect 20478 48738 20560 48982
rect 20654 48742 20766 48758
rect 20654 48738 20678 48742
rect 20478 48698 20678 48738
rect 19054 48390 19634 48400
rect 19054 48386 20394 48390
rect 20478 48386 20560 48698
rect 20654 48690 20678 48698
rect 20750 48690 20766 48742
rect 20654 48666 20766 48690
rect 19054 48380 20560 48386
rect 19054 48346 19544 48380
rect 19716 48346 20238 48380
rect 20410 48346 20560 48380
rect 19054 48332 20560 48346
rect 19054 48310 19634 48332
rect 20336 48318 20560 48332
rect 19352 48304 19634 48310
rect 20280 47746 20410 47766
rect 20478 47746 20560 48318
rect 20280 47734 20560 47746
rect 19592 47722 20560 47734
rect 15752 47682 15974 47688
rect 18378 47686 18600 47692
rect 19528 47688 19544 47722
rect 19716 47688 20238 47722
rect 20410 47688 20560 47722
rect 1030 47672 2678 47680
rect 5124 47676 5346 47682
rect 922 47638 938 47672
rect 1110 47638 1632 47672
rect 1804 47638 2326 47672
rect 2498 47638 2678 47672
rect 3698 47668 5346 47676
rect 6372 47674 8020 47682
rect 9018 47674 10666 47682
rect 13098 47676 13320 47682
rect 1030 47628 2678 47638
rect 3590 47634 3606 47668
rect 3778 47634 4300 47668
rect 4472 47634 4994 47668
rect 5166 47634 5346 47668
rect 6264 47640 6280 47674
rect 6452 47640 6974 47674
rect 7146 47640 7668 47674
rect 7840 47640 8020 47674
rect 8910 47640 8926 47674
rect 9098 47640 9620 47674
rect 9792 47640 10314 47674
rect 10486 47640 10666 47674
rect 11672 47668 13320 47676
rect 14326 47674 15974 47682
rect 16952 47678 18600 47686
rect 2456 47616 2678 47628
rect 3698 47624 5346 47634
rect 6372 47630 8020 47640
rect 9018 47630 10666 47640
rect 11564 47634 11580 47668
rect 11752 47634 12274 47668
rect 12446 47634 12968 47668
rect 13140 47634 13320 47668
rect 14218 47640 14234 47674
rect 14406 47640 14928 47674
rect 15100 47640 15622 47674
rect 15794 47640 15974 47674
rect 16844 47644 16860 47678
rect 17032 47644 17554 47678
rect 17726 47644 18248 47678
rect 18420 47644 18600 47678
rect 19592 47676 20560 47688
rect 5124 47612 5346 47624
rect 7798 47618 8020 47630
rect 10444 47618 10666 47630
rect 11672 47624 13320 47634
rect 14326 47630 15974 47640
rect 16952 47634 18600 47644
rect 13098 47612 13320 47624
rect 15752 47618 15974 47630
rect 18378 47622 18600 47634
rect 9038 47404 10634 47430
rect 2460 47370 4416 47400
rect 2460 47240 2592 47370
rect 4384 47240 4416 47370
rect 2460 47210 4416 47240
rect 9038 47244 9118 47404
rect 10578 47244 10634 47404
rect 9038 47202 10634 47244
rect 14164 47386 15696 47416
rect 14164 47226 14218 47386
rect 15628 47226 15696 47386
rect 14164 47188 15696 47226
rect 16962 47408 18414 47434
rect 20280 47412 20410 47676
rect 20478 47670 20560 47676
rect 16962 47262 17048 47408
rect 18368 47262 18414 47408
rect 16962 47206 18414 47262
rect 19406 47378 20524 47412
rect 19406 47222 19456 47378
rect 20474 47222 20524 47378
rect 19406 47190 20524 47222
rect 24498 45070 24856 51900
rect 42138 51138 42220 52630
rect 46164 52628 46246 52630
rect 50176 52628 50258 52630
rect 54186 52628 54268 52630
rect 42670 52274 45316 52310
rect 42670 51942 42820 52274
rect 45220 51942 45316 52274
rect 42670 51908 45316 51942
rect 46664 52274 49310 52310
rect 46664 51942 46814 52274
rect 49214 51942 49310 52274
rect 46664 51908 49310 51942
rect 50686 52274 53332 52310
rect 50686 51942 50836 52274
rect 53236 51942 53332 52274
rect 50686 51908 53332 51942
rect 54708 52274 57354 52310
rect 54708 51942 54858 52274
rect 57258 51942 57354 52274
rect 54708 51908 57354 51942
rect 57422 52304 57508 53278
rect 57610 52376 57800 52450
rect 57610 52304 57626 52376
rect 57422 52054 57626 52304
rect 57422 51800 57508 52054
rect 57610 51974 57626 52054
rect 57772 51974 57800 52376
rect 57610 51908 57800 51974
rect 45202 51782 45466 51800
rect 49196 51782 49460 51800
rect 53218 51782 53482 51800
rect 57240 51782 57508 51800
rect 42400 51770 57508 51782
rect 42310 51736 42326 51770
rect 42498 51736 43020 51770
rect 43192 51736 43714 51770
rect 43886 51736 44408 51770
rect 44580 51736 45102 51770
rect 45274 51736 46320 51770
rect 46492 51736 47014 51770
rect 47186 51736 47708 51770
rect 47880 51736 48402 51770
rect 48574 51736 49096 51770
rect 49268 51736 50342 51770
rect 50514 51736 51036 51770
rect 51208 51736 51730 51770
rect 51902 51736 52424 51770
rect 52596 51736 53118 51770
rect 53290 51736 54364 51770
rect 54536 51736 55058 51770
rect 55230 51736 55752 51770
rect 55924 51736 56446 51770
rect 56618 51736 57140 51770
rect 57312 51736 57508 51770
rect 42400 51732 57508 51736
rect 42400 51730 57504 51732
rect 42400 51728 45466 51730
rect 46394 51728 49460 51730
rect 50416 51728 53482 51730
rect 54438 51728 57504 51730
rect 45202 51724 45466 51728
rect 49196 51724 49460 51728
rect 53218 51724 53482 51728
rect 57240 51724 57504 51728
rect 42138 51124 42434 51138
rect 42138 51112 45284 51124
rect 42138 51078 42326 51112
rect 42498 51078 43020 51112
rect 43192 51078 43714 51112
rect 43886 51078 44408 51112
rect 44580 51078 45102 51112
rect 45274 51078 45290 51112
rect 42138 51070 45284 51078
rect 42138 51062 42434 51070
rect 42138 50962 42230 51062
rect 42148 49816 42230 50962
rect 45388 50472 45442 51724
rect 46142 51124 46428 51138
rect 46142 51112 49278 51124
rect 46142 51078 46320 51112
rect 46492 51078 47014 51112
rect 47186 51078 47708 51112
rect 47880 51078 48402 51112
rect 48574 51078 49096 51112
rect 49268 51078 49284 51112
rect 46142 51070 49278 51078
rect 46142 51062 46428 51070
rect 45238 50466 45502 50472
rect 42448 50454 45502 50466
rect 42310 50420 42326 50454
rect 42498 50420 43020 50454
rect 43192 50420 43714 50454
rect 43886 50420 44408 50454
rect 44580 50420 45102 50454
rect 45274 50420 45502 50454
rect 42448 50412 45502 50420
rect 45238 50396 45502 50412
rect 42144 49808 42464 49816
rect 42144 49796 45292 49808
rect 42144 49762 42326 49796
rect 42498 49762 43020 49796
rect 43192 49762 43714 49796
rect 43886 49762 44408 49796
rect 44580 49762 45102 49796
rect 45274 49762 45292 49796
rect 42144 49754 45292 49762
rect 42144 49740 42464 49754
rect 42148 48510 42230 49740
rect 45388 49158 45442 50396
rect 46142 49816 46224 51062
rect 49382 50472 49436 51724
rect 50164 51124 50450 51138
rect 50164 51112 53300 51124
rect 50164 51078 50342 51112
rect 50514 51078 51036 51112
rect 51208 51078 51730 51112
rect 51902 51078 52424 51112
rect 52596 51078 53118 51112
rect 53290 51078 53306 51112
rect 50164 51070 53300 51078
rect 50164 51062 50450 51070
rect 49232 50466 49496 50472
rect 46442 50454 49496 50466
rect 46304 50420 46320 50454
rect 46492 50420 47014 50454
rect 47186 50420 47708 50454
rect 47880 50420 48402 50454
rect 48574 50420 49096 50454
rect 49268 50420 49496 50454
rect 46442 50412 49496 50420
rect 49232 50396 49496 50412
rect 46138 49808 46458 49816
rect 46138 49796 49286 49808
rect 46138 49762 46320 49796
rect 46492 49762 47014 49796
rect 47186 49762 47708 49796
rect 47880 49762 48402 49796
rect 48574 49762 49096 49796
rect 49268 49762 49286 49796
rect 46138 49754 49286 49762
rect 46138 49740 46458 49754
rect 45208 49144 45472 49158
rect 42446 49138 45472 49144
rect 42310 49104 42326 49138
rect 42498 49104 43020 49138
rect 43192 49104 43714 49138
rect 43886 49104 44408 49138
rect 44580 49104 45102 49138
rect 45274 49104 45472 49138
rect 42446 49090 45472 49104
rect 45208 49082 45472 49090
rect 45388 49080 45442 49082
rect 46142 48510 46224 49740
rect 49382 49158 49436 50396
rect 50164 49816 50246 51062
rect 53404 50472 53458 51724
rect 57386 51582 57480 51724
rect 54186 51124 54472 51138
rect 54186 51112 57322 51124
rect 54186 51078 54364 51112
rect 54536 51078 55058 51112
rect 55230 51078 55752 51112
rect 55924 51078 56446 51112
rect 56618 51078 57140 51112
rect 57312 51078 57328 51112
rect 54186 51070 57322 51078
rect 54186 51062 54472 51070
rect 53254 50466 53518 50472
rect 50464 50454 53518 50466
rect 50326 50420 50342 50454
rect 50514 50420 51036 50454
rect 51208 50420 51730 50454
rect 51902 50420 52424 50454
rect 52596 50420 53118 50454
rect 53290 50420 53518 50454
rect 50464 50412 53518 50420
rect 53254 50396 53518 50412
rect 50160 49808 50480 49816
rect 50160 49796 53308 49808
rect 50160 49762 50342 49796
rect 50514 49762 51036 49796
rect 51208 49762 51730 49796
rect 51902 49762 52424 49796
rect 52596 49762 53118 49796
rect 53290 49762 53308 49796
rect 50160 49754 53308 49762
rect 50160 49740 50480 49754
rect 49202 49144 49466 49158
rect 46440 49138 49466 49144
rect 46304 49104 46320 49138
rect 46492 49104 47014 49138
rect 47186 49104 47708 49138
rect 47880 49104 48402 49138
rect 48574 49104 49096 49138
rect 49268 49104 49466 49138
rect 46440 49090 49466 49104
rect 49202 49082 49466 49090
rect 49382 49080 49436 49082
rect 50164 48510 50246 49740
rect 53404 49158 53458 50396
rect 54186 49816 54268 51062
rect 57426 50472 57480 51582
rect 57276 50466 57540 50472
rect 54486 50454 57540 50466
rect 54348 50420 54364 50454
rect 54536 50420 55058 50454
rect 55230 50420 55752 50454
rect 55924 50420 56446 50454
rect 56618 50420 57140 50454
rect 57312 50420 57540 50454
rect 54486 50412 57540 50420
rect 57276 50396 57540 50412
rect 54182 49808 54502 49816
rect 54182 49796 57330 49808
rect 54182 49762 54364 49796
rect 54536 49762 55058 49796
rect 55230 49762 55752 49796
rect 55924 49762 56446 49796
rect 56618 49762 57140 49796
rect 57312 49762 57330 49796
rect 54182 49754 57330 49762
rect 54182 49740 54502 49754
rect 53224 49144 53488 49158
rect 50462 49138 53488 49144
rect 50326 49104 50342 49138
rect 50514 49104 51036 49138
rect 51208 49104 51730 49138
rect 51902 49104 52424 49138
rect 52596 49104 53118 49138
rect 53290 49104 53488 49138
rect 50462 49090 53488 49104
rect 53224 49082 53488 49090
rect 53404 49080 53458 49082
rect 54186 48510 54268 49740
rect 57426 49184 57480 50396
rect 57366 49158 57502 49184
rect 57246 49144 57510 49158
rect 54484 49138 57510 49144
rect 54348 49104 54364 49138
rect 54536 49104 55058 49138
rect 55230 49104 55752 49138
rect 55924 49104 56446 49138
rect 56618 49104 57140 49138
rect 57312 49104 57510 49138
rect 54484 49090 57510 49104
rect 57246 49082 57510 49090
rect 57024 48512 57212 48522
rect 57366 48512 57502 49082
rect 42144 48498 42444 48510
rect 46138 48498 46438 48510
rect 50160 48498 50460 48510
rect 54182 48498 54482 48510
rect 57024 48498 57532 48512
rect 42144 48480 57532 48498
rect 42144 48446 42326 48480
rect 42498 48446 43020 48480
rect 43192 48446 43714 48480
rect 43886 48446 44408 48480
rect 44580 48446 45102 48480
rect 45274 48446 46320 48480
rect 46492 48446 47014 48480
rect 47186 48446 47708 48480
rect 47880 48446 48402 48480
rect 48574 48446 49096 48480
rect 49268 48446 50342 48480
rect 50514 48446 51036 48480
rect 51208 48446 51730 48480
rect 51902 48446 52424 48480
rect 52596 48446 53118 48480
rect 53290 48446 54364 48480
rect 54536 48446 55058 48480
rect 55230 48446 55752 48480
rect 55924 48446 56446 48480
rect 56618 48446 57140 48480
rect 57312 48446 57532 48480
rect 42144 48436 45286 48446
rect 46138 48436 49280 48446
rect 50160 48436 53302 48446
rect 54182 48436 57532 48446
rect 42144 48434 42426 48436
rect 46138 48434 46420 48436
rect 50160 48434 50442 48436
rect 54182 48434 54464 48436
rect 42148 48432 42230 48434
rect 46142 48432 46224 48434
rect 50164 48432 50246 48434
rect 54186 48432 54268 48434
rect 57024 48408 57532 48436
rect 42620 48166 44984 48258
rect 57024 48218 57212 48408
rect 42620 47902 42766 48166
rect 44904 47902 44984 48166
rect 42620 47836 44984 47902
rect 46528 48178 49418 48218
rect 46528 47914 46660 48178
rect 49352 47914 49418 48178
rect 46528 47862 49418 47914
rect 50606 48140 53444 48206
rect 50606 47914 50790 48140
rect 53312 47914 53444 48140
rect 50606 47848 53444 47914
rect 54354 48152 57272 48218
rect 54354 47928 54448 48152
rect 57206 47928 57272 48152
rect 54354 47862 57272 47928
rect 57024 47840 57212 47862
rect 58938 46504 59118 56840
rect 71008 55234 71038 57980
rect 71178 55234 71224 57980
rect 71008 55180 71224 55234
rect 71292 57868 71306 58040
rect 71340 57868 71348 58040
rect 71964 58040 71998 58056
rect 71292 57346 71348 57868
rect 71292 57174 71306 57346
rect 71340 57174 71348 57346
rect 71292 56652 71348 57174
rect 71292 56480 71306 56652
rect 71340 56480 71348 56652
rect 71292 55958 71348 56480
rect 71292 55786 71306 55958
rect 71340 55786 71348 55958
rect 71292 55368 71348 55786
rect 71954 57868 71964 58024
rect 72610 58040 72666 58146
rect 73920 58136 74106 58146
rect 75152 58168 75228 58848
rect 75808 58848 75828 58980
rect 75862 58936 75874 59020
rect 76472 61624 76486 61776
rect 76520 61744 76530 61796
rect 77144 61796 77178 61812
rect 76520 61624 76528 61744
rect 76472 61102 76528 61624
rect 76472 60930 76486 61102
rect 76520 60930 76528 61102
rect 76472 60408 76528 60930
rect 76472 60236 76486 60408
rect 76520 60236 76528 60408
rect 76472 59714 76528 60236
rect 76472 59542 76486 59714
rect 76520 59542 76528 59714
rect 76472 59020 76528 59542
rect 75862 58848 75868 58936
rect 76472 58932 76486 59020
rect 75808 58738 75868 58848
rect 76520 58932 76528 59020
rect 77132 61624 77144 61734
rect 77784 61796 77860 61892
rect 79006 61810 79062 61916
rect 77178 61624 77188 61734
rect 77784 61714 77802 61796
rect 77132 61102 77188 61624
rect 77132 60930 77144 61102
rect 77178 60930 77188 61102
rect 77132 60408 77188 60930
rect 77132 60236 77144 60408
rect 77178 60236 77188 60408
rect 77132 59714 77188 60236
rect 77132 59542 77144 59714
rect 77178 59542 77188 59714
rect 77132 59020 77188 59542
rect 77132 58890 77144 59020
rect 76486 58832 76520 58848
rect 77136 58848 77144 58890
rect 77178 58978 77188 59020
rect 77786 61624 77802 61714
rect 77836 61714 77860 61796
rect 78722 61750 78938 61810
rect 77836 61624 77842 61714
rect 77786 61102 77842 61624
rect 77786 60930 77802 61102
rect 77836 60930 77842 61102
rect 77786 60408 77842 60930
rect 77786 60236 77802 60408
rect 77836 60236 77842 60408
rect 77786 59714 77842 60236
rect 77786 59542 77802 59714
rect 77836 59542 77842 59714
rect 77786 59020 77842 59542
rect 77178 58848 77196 58978
rect 77786 58894 77802 59020
rect 77136 58742 77196 58848
rect 77836 58894 77842 59020
rect 78722 59004 78752 61750
rect 78892 59004 78938 61750
rect 79006 61638 79020 61810
rect 79054 61638 79062 61810
rect 79678 61810 79712 61826
rect 79006 61116 79062 61638
rect 79006 60944 79020 61116
rect 79054 60944 79062 61116
rect 79006 60422 79062 60944
rect 79006 60250 79020 60422
rect 79054 60250 79062 60422
rect 79006 59728 79062 60250
rect 79006 59556 79020 59728
rect 79054 59556 79062 59728
rect 79006 59150 79062 59556
rect 79668 61638 79678 61794
rect 80324 61810 80380 61916
rect 81634 61906 81820 61916
rect 79712 61638 79724 61794
rect 80324 61790 80336 61810
rect 79668 61116 79724 61638
rect 79668 60944 79678 61116
rect 79712 60944 79724 61116
rect 79668 60422 79724 60944
rect 79668 60250 79678 60422
rect 79712 60250 79724 60422
rect 79668 59728 79724 60250
rect 79668 59556 79678 59728
rect 79712 59556 79724 59728
rect 78722 58950 78938 59004
rect 79002 59034 79078 59150
rect 77802 58832 77836 58848
rect 79002 58862 79020 59034
rect 79054 58862 79078 59034
rect 79668 59034 79724 59556
rect 79668 58994 79678 59034
rect 77136 58738 77294 58742
rect 75808 58676 77294 58738
rect 75808 58670 75868 58676
rect 77136 58668 77196 58676
rect 77792 58176 77970 58186
rect 77784 58168 77970 58176
rect 71998 57868 72010 58024
rect 72610 58020 72622 58040
rect 71954 57346 72010 57868
rect 71954 57174 71964 57346
rect 71998 57174 72010 57346
rect 71954 56652 72010 57174
rect 71954 56480 71964 56652
rect 71998 56480 72010 56652
rect 71954 55958 72010 56480
rect 71954 55786 71964 55958
rect 71998 55786 72010 55958
rect 71292 55264 71372 55368
rect 71292 55192 71306 55264
rect 71296 55092 71306 55192
rect 71340 55092 71372 55264
rect 71954 55264 72010 55786
rect 71954 55224 71964 55264
rect 71296 54416 71372 55092
rect 71944 55092 71964 55224
rect 71998 55180 72010 55264
rect 72608 57868 72622 58020
rect 72656 57988 72666 58040
rect 73280 58040 73314 58056
rect 72656 57868 72664 57988
rect 72608 57346 72664 57868
rect 72608 57174 72622 57346
rect 72656 57174 72664 57346
rect 72608 56652 72664 57174
rect 72608 56480 72622 56652
rect 72656 56480 72664 56652
rect 72608 55958 72664 56480
rect 72608 55786 72622 55958
rect 72656 55786 72664 55958
rect 72608 55264 72664 55786
rect 71998 55092 72004 55180
rect 72608 55176 72622 55264
rect 71944 54982 72004 55092
rect 72656 55176 72664 55264
rect 73268 57868 73280 57978
rect 73920 58040 73996 58136
rect 75152 58126 77970 58168
rect 75152 58068 75228 58126
rect 73314 57868 73324 57978
rect 73920 57958 73938 58040
rect 73268 57346 73324 57868
rect 73268 57174 73280 57346
rect 73314 57174 73324 57346
rect 73268 56652 73324 57174
rect 73268 56480 73280 56652
rect 73314 56480 73324 56652
rect 73268 55958 73324 56480
rect 73268 55786 73280 55958
rect 73314 55786 73324 55958
rect 73268 55264 73324 55786
rect 73268 55134 73280 55264
rect 72622 55076 72656 55092
rect 73272 55092 73280 55134
rect 73314 55222 73324 55264
rect 73922 57868 73938 57958
rect 73972 57958 73996 58040
rect 75156 58020 75212 58068
rect 74872 57960 75088 58020
rect 73972 57868 73978 57958
rect 73922 57346 73978 57868
rect 73922 57174 73938 57346
rect 73972 57174 73978 57346
rect 73922 56652 73978 57174
rect 73922 56480 73938 56652
rect 73972 56480 73978 56652
rect 73922 55958 73978 56480
rect 73922 55786 73938 55958
rect 73972 55786 73978 55958
rect 73922 55264 73978 55786
rect 73314 55092 73332 55222
rect 73922 55138 73938 55264
rect 73272 54986 73332 55092
rect 73972 55138 73978 55264
rect 74872 55214 74902 57960
rect 75042 55214 75088 57960
rect 74872 55160 75088 55214
rect 75156 57848 75170 58020
rect 75204 57848 75212 58020
rect 75828 58020 75862 58036
rect 75156 57326 75212 57848
rect 75156 57154 75170 57326
rect 75204 57154 75212 57326
rect 75156 56632 75212 57154
rect 75156 56460 75170 56632
rect 75204 56460 75212 56632
rect 75156 55938 75212 56460
rect 75156 55766 75170 55938
rect 75204 55766 75212 55938
rect 75156 55348 75212 55766
rect 75818 57848 75828 58004
rect 76474 58020 76530 58126
rect 77784 58116 77970 58126
rect 79002 58182 79078 58862
rect 79658 58862 79678 58994
rect 79712 58950 79724 59034
rect 80322 61638 80336 61790
rect 80370 61758 80380 61810
rect 80994 61810 81028 61826
rect 80370 61638 80378 61758
rect 80322 61116 80378 61638
rect 80322 60944 80336 61116
rect 80370 60944 80378 61116
rect 80322 60422 80378 60944
rect 80322 60250 80336 60422
rect 80370 60250 80378 60422
rect 80322 59728 80378 60250
rect 80322 59556 80336 59728
rect 80370 59556 80378 59728
rect 80322 59034 80378 59556
rect 79712 58862 79718 58950
rect 80322 58946 80336 59034
rect 79658 58752 79718 58862
rect 80370 58946 80378 59034
rect 80982 61638 80994 61748
rect 81634 61810 81710 61906
rect 81028 61638 81038 61748
rect 81634 61728 81652 61810
rect 80982 61116 81038 61638
rect 80982 60944 80994 61116
rect 81028 60944 81038 61116
rect 80982 60422 81038 60944
rect 80982 60250 80994 60422
rect 81028 60250 81038 60422
rect 80982 59728 81038 60250
rect 80982 59556 80994 59728
rect 81028 59556 81038 59728
rect 80982 59034 81038 59556
rect 80982 58904 80994 59034
rect 80336 58846 80370 58862
rect 80986 58862 80994 58904
rect 81028 58992 81038 59034
rect 81636 61638 81652 61728
rect 81686 61728 81710 61810
rect 81686 61638 81692 61728
rect 81636 61116 81692 61638
rect 81636 60944 81652 61116
rect 81686 60944 81692 61116
rect 81636 60422 81692 60944
rect 81636 60250 81652 60422
rect 81686 60250 81692 60422
rect 81636 59728 81692 60250
rect 81636 59556 81652 59728
rect 81686 59556 81692 59728
rect 81636 59034 81692 59556
rect 81028 58862 81046 58992
rect 81636 58908 81652 59034
rect 80986 58756 81046 58862
rect 81686 58908 81692 59034
rect 81652 58846 81686 58862
rect 80986 58752 81144 58756
rect 79658 58690 81144 58752
rect 79658 58684 79718 58690
rect 80986 58682 81046 58690
rect 81642 58190 81820 58200
rect 81634 58182 81820 58190
rect 79002 58140 81820 58182
rect 75862 57848 75874 58004
rect 76474 58000 76486 58020
rect 75818 57326 75874 57848
rect 75818 57154 75828 57326
rect 75862 57154 75874 57326
rect 75818 56632 75874 57154
rect 75818 56460 75828 56632
rect 75862 56460 75874 56632
rect 75818 55938 75874 56460
rect 75818 55766 75828 55938
rect 75862 55766 75874 55938
rect 75156 55244 75236 55348
rect 75156 55172 75170 55244
rect 73938 55076 73972 55092
rect 75160 55072 75170 55172
rect 75204 55072 75236 55244
rect 75818 55244 75874 55766
rect 75818 55204 75828 55244
rect 73272 54982 73430 54986
rect 71944 54920 73430 54982
rect 71944 54914 72004 54920
rect 73272 54912 73332 54920
rect 73932 54424 74110 54434
rect 73924 54416 74110 54424
rect 71292 54374 74110 54416
rect 75160 54396 75236 55072
rect 75808 55072 75828 55204
rect 75862 55160 75874 55244
rect 76472 57848 76486 58000
rect 76520 57968 76530 58020
rect 77144 58020 77178 58036
rect 76520 57848 76528 57968
rect 76472 57326 76528 57848
rect 76472 57154 76486 57326
rect 76520 57154 76528 57326
rect 76472 56632 76528 57154
rect 76472 56460 76486 56632
rect 76520 56460 76528 56632
rect 76472 55938 76528 56460
rect 76472 55766 76486 55938
rect 76520 55766 76528 55938
rect 76472 55244 76528 55766
rect 75862 55072 75868 55160
rect 76472 55156 76486 55244
rect 75808 54962 75868 55072
rect 76520 55156 76528 55244
rect 77132 57848 77144 57958
rect 77784 58020 77860 58116
rect 79002 58082 79078 58140
rect 79006 58034 79062 58082
rect 77178 57848 77188 57958
rect 77784 57938 77802 58020
rect 77132 57326 77188 57848
rect 77132 57154 77144 57326
rect 77178 57154 77188 57326
rect 77132 56632 77188 57154
rect 77132 56460 77144 56632
rect 77178 56460 77188 56632
rect 77132 55938 77188 56460
rect 77132 55766 77144 55938
rect 77178 55766 77188 55938
rect 77132 55244 77188 55766
rect 77132 55114 77144 55244
rect 76486 55056 76520 55072
rect 77136 55072 77144 55114
rect 77178 55202 77188 55244
rect 77786 57848 77802 57938
rect 77836 57938 77860 58020
rect 78722 57974 78938 58034
rect 77836 57848 77842 57938
rect 77786 57326 77842 57848
rect 77786 57154 77802 57326
rect 77836 57154 77842 57326
rect 77786 56632 77842 57154
rect 77786 56460 77802 56632
rect 77836 56460 77842 56632
rect 77786 55938 77842 56460
rect 77786 55766 77802 55938
rect 77836 55766 77842 55938
rect 77786 55244 77842 55766
rect 77178 55072 77196 55202
rect 77786 55118 77802 55244
rect 77136 54966 77196 55072
rect 77836 55118 77842 55244
rect 78722 55228 78752 57974
rect 78892 55228 78938 57974
rect 78722 55174 78938 55228
rect 79006 57862 79020 58034
rect 79054 57862 79062 58034
rect 79678 58034 79712 58050
rect 79006 57340 79062 57862
rect 79006 57168 79020 57340
rect 79054 57168 79062 57340
rect 79006 56646 79062 57168
rect 79006 56474 79020 56646
rect 79054 56474 79062 56646
rect 79006 55952 79062 56474
rect 79006 55780 79020 55952
rect 79054 55780 79062 55952
rect 79006 55362 79062 55780
rect 79668 57862 79678 58018
rect 80324 58034 80380 58140
rect 81634 58130 81820 58140
rect 79712 57862 79724 58018
rect 80324 58014 80336 58034
rect 79668 57340 79724 57862
rect 79668 57168 79678 57340
rect 79712 57168 79724 57340
rect 79668 56646 79724 57168
rect 79668 56474 79678 56646
rect 79712 56474 79724 56646
rect 79668 55952 79724 56474
rect 79668 55780 79678 55952
rect 79712 55780 79724 55952
rect 79006 55258 79086 55362
rect 79006 55186 79020 55258
rect 77802 55056 77836 55072
rect 79010 55086 79020 55186
rect 79054 55086 79086 55258
rect 79668 55258 79724 55780
rect 79668 55218 79678 55258
rect 77136 54962 77294 54966
rect 75808 54900 77294 54962
rect 75808 54894 75868 54900
rect 77136 54892 77196 54900
rect 77796 54404 77974 54414
rect 79010 54410 79086 55086
rect 79658 55086 79678 55218
rect 79712 55174 79724 55258
rect 80322 57862 80336 58014
rect 80370 57982 80380 58034
rect 80994 58034 81028 58050
rect 80370 57862 80378 57982
rect 80322 57340 80378 57862
rect 80322 57168 80336 57340
rect 80370 57168 80378 57340
rect 80322 56646 80378 57168
rect 80322 56474 80336 56646
rect 80370 56474 80378 56646
rect 80322 55952 80378 56474
rect 80322 55780 80336 55952
rect 80370 55780 80378 55952
rect 80322 55258 80378 55780
rect 79712 55086 79718 55174
rect 80322 55170 80336 55258
rect 79658 54976 79718 55086
rect 80370 55170 80378 55258
rect 80982 57862 80994 57972
rect 81634 58034 81710 58130
rect 81028 57862 81038 57972
rect 81634 57952 81652 58034
rect 80982 57340 81038 57862
rect 80982 57168 80994 57340
rect 81028 57168 81038 57340
rect 80982 56646 81038 57168
rect 80982 56474 80994 56646
rect 81028 56474 81038 56646
rect 80982 55952 81038 56474
rect 80982 55780 80994 55952
rect 81028 55780 81038 55952
rect 80982 55258 81038 55780
rect 80982 55128 80994 55258
rect 80336 55070 80370 55086
rect 80986 55086 80994 55128
rect 81028 55216 81038 55258
rect 81636 57862 81652 57952
rect 81686 57952 81710 58034
rect 81686 57862 81692 57952
rect 81636 57340 81692 57862
rect 81636 57168 81652 57340
rect 81686 57168 81692 57340
rect 81636 56646 81692 57168
rect 81636 56474 81652 56646
rect 81686 56474 81692 56646
rect 81636 55952 81692 56474
rect 81636 55780 81652 55952
rect 81686 55780 81692 55952
rect 81636 55258 81692 55780
rect 81028 55086 81046 55216
rect 81636 55132 81652 55258
rect 80986 54980 81046 55086
rect 81686 55132 81692 55258
rect 81652 55070 81686 55086
rect 80986 54976 81144 54980
rect 79658 54914 81144 54976
rect 81894 54946 81928 54954
rect 81894 54936 82128 54946
rect 81894 54918 81910 54936
rect 79658 54908 79718 54914
rect 80986 54906 81046 54914
rect 81646 54418 81824 54428
rect 81638 54410 81824 54418
rect 77788 54396 77974 54404
rect 71296 54300 71372 54374
rect 71296 54268 71352 54300
rect 71012 54208 71228 54268
rect 71012 51462 71042 54208
rect 71182 51462 71228 54208
rect 71012 51408 71228 51462
rect 71296 54096 71310 54268
rect 71344 54096 71352 54268
rect 71968 54268 72002 54284
rect 71296 53574 71352 54096
rect 71296 53402 71310 53574
rect 71344 53402 71352 53574
rect 71296 52880 71352 53402
rect 71296 52708 71310 52880
rect 71344 52708 71352 52880
rect 71296 52186 71352 52708
rect 71296 52014 71310 52186
rect 71344 52014 71352 52186
rect 71296 51492 71352 52014
rect 71296 51420 71310 51492
rect 71344 51420 71352 51492
rect 71958 54096 71968 54252
rect 72614 54268 72670 54374
rect 73924 54364 74110 54374
rect 72002 54096 72014 54252
rect 72614 54248 72626 54268
rect 71958 53574 72014 54096
rect 71958 53402 71968 53574
rect 72002 53402 72014 53574
rect 71958 52880 72014 53402
rect 71958 52708 71968 52880
rect 72002 52708 72014 52880
rect 71958 52186 72014 52708
rect 71958 52014 71968 52186
rect 72002 52014 72014 52186
rect 71958 51492 72014 52014
rect 71958 51452 71968 51492
rect 71310 51304 71344 51320
rect 71948 51320 71968 51452
rect 72002 51408 72014 51492
rect 72612 54096 72626 54248
rect 72660 54216 72670 54268
rect 73284 54268 73318 54284
rect 72660 54096 72668 54216
rect 72612 53574 72668 54096
rect 72612 53402 72626 53574
rect 72660 53402 72668 53574
rect 72612 52880 72668 53402
rect 72612 52708 72626 52880
rect 72660 52708 72668 52880
rect 72612 52186 72668 52708
rect 72612 52014 72626 52186
rect 72660 52014 72668 52186
rect 72612 51492 72668 52014
rect 72002 51320 72008 51408
rect 72612 51404 72626 51492
rect 71948 51210 72008 51320
rect 72660 51404 72668 51492
rect 73272 54096 73284 54206
rect 73924 54268 74000 54364
rect 75156 54354 77974 54396
rect 79006 54368 81824 54410
rect 73318 54096 73328 54206
rect 73924 54186 73942 54268
rect 73272 53574 73328 54096
rect 73272 53402 73284 53574
rect 73318 53402 73328 53574
rect 73272 52880 73328 53402
rect 73272 52708 73284 52880
rect 73318 52708 73328 52880
rect 73272 52186 73328 52708
rect 73272 52014 73284 52186
rect 73318 52014 73328 52186
rect 73272 51492 73328 52014
rect 73272 51362 73284 51492
rect 72626 51304 72660 51320
rect 73276 51320 73284 51362
rect 73318 51450 73328 51492
rect 73926 54096 73942 54186
rect 73976 54186 74000 54268
rect 75160 54280 75236 54354
rect 75160 54248 75216 54280
rect 74876 54188 75092 54248
rect 73976 54096 73982 54186
rect 73926 53574 73982 54096
rect 73926 53402 73942 53574
rect 73976 53402 73982 53574
rect 73926 52880 73982 53402
rect 73926 52708 73942 52880
rect 73976 52708 73982 52880
rect 73926 52186 73982 52708
rect 73926 52014 73942 52186
rect 73976 52014 73982 52186
rect 73926 51492 73982 52014
rect 73318 51320 73336 51450
rect 73926 51366 73942 51492
rect 73276 51214 73336 51320
rect 73976 51366 73982 51492
rect 74876 51442 74906 54188
rect 75046 51442 75092 54188
rect 74876 51388 75092 51442
rect 75160 54076 75174 54248
rect 75208 54076 75216 54248
rect 75832 54248 75866 54264
rect 75160 53554 75216 54076
rect 75160 53382 75174 53554
rect 75208 53382 75216 53554
rect 75160 52860 75216 53382
rect 75160 52688 75174 52860
rect 75208 52688 75216 52860
rect 75160 52166 75216 52688
rect 75160 51994 75174 52166
rect 75208 51994 75216 52166
rect 75160 51472 75216 51994
rect 75160 51400 75174 51472
rect 73942 51304 73976 51320
rect 75208 51400 75216 51472
rect 75822 54076 75832 54232
rect 76478 54248 76534 54354
rect 77788 54344 77974 54354
rect 75866 54076 75878 54232
rect 76478 54228 76490 54248
rect 75822 53554 75878 54076
rect 75822 53382 75832 53554
rect 75866 53382 75878 53554
rect 75822 52860 75878 53382
rect 75822 52688 75832 52860
rect 75866 52688 75878 52860
rect 75822 52166 75878 52688
rect 75822 51994 75832 52166
rect 75866 51994 75878 52166
rect 75822 51472 75878 51994
rect 75822 51432 75832 51472
rect 75174 51284 75208 51300
rect 75812 51300 75832 51432
rect 75866 51388 75878 51472
rect 76476 54076 76490 54228
rect 76524 54196 76534 54248
rect 77148 54248 77182 54264
rect 76524 54076 76532 54196
rect 76476 53554 76532 54076
rect 76476 53382 76490 53554
rect 76524 53382 76532 53554
rect 76476 52860 76532 53382
rect 76476 52688 76490 52860
rect 76524 52688 76532 52860
rect 76476 52166 76532 52688
rect 76476 51994 76490 52166
rect 76524 51994 76532 52166
rect 76476 51472 76532 51994
rect 75866 51300 75872 51388
rect 76476 51384 76490 51472
rect 73276 51210 73434 51214
rect 71948 51148 73434 51210
rect 75812 51190 75872 51300
rect 76524 51384 76532 51472
rect 77136 54076 77148 54186
rect 77788 54248 77864 54344
rect 79010 54294 79086 54368
rect 79010 54262 79066 54294
rect 77182 54076 77192 54186
rect 77788 54166 77806 54248
rect 77136 53554 77192 54076
rect 77136 53382 77148 53554
rect 77182 53382 77192 53554
rect 77136 52860 77192 53382
rect 77136 52688 77148 52860
rect 77182 52688 77192 52860
rect 77136 52166 77192 52688
rect 77136 51994 77148 52166
rect 77182 51994 77192 52166
rect 77136 51472 77192 51994
rect 77136 51342 77148 51472
rect 76490 51284 76524 51300
rect 77140 51300 77148 51342
rect 77182 51430 77192 51472
rect 77790 54076 77806 54166
rect 77840 54166 77864 54248
rect 78726 54202 78942 54262
rect 77840 54076 77846 54166
rect 77790 53554 77846 54076
rect 77790 53382 77806 53554
rect 77840 53382 77846 53554
rect 77790 52860 77846 53382
rect 77790 52688 77806 52860
rect 77840 52688 77846 52860
rect 77790 52166 77846 52688
rect 77790 51994 77806 52166
rect 77840 51994 77846 52166
rect 77790 51472 77846 51994
rect 77182 51300 77200 51430
rect 77790 51346 77806 51472
rect 77140 51194 77200 51300
rect 77840 51346 77846 51472
rect 78726 51456 78756 54202
rect 78896 51456 78942 54202
rect 78726 51402 78942 51456
rect 79010 54090 79024 54262
rect 79058 54090 79066 54262
rect 79682 54262 79716 54278
rect 79010 53568 79066 54090
rect 79010 53396 79024 53568
rect 79058 53396 79066 53568
rect 79010 52874 79066 53396
rect 79010 52702 79024 52874
rect 79058 52702 79066 52874
rect 79010 52180 79066 52702
rect 79010 52008 79024 52180
rect 79058 52008 79066 52180
rect 79010 51486 79066 52008
rect 79010 51414 79024 51486
rect 77806 51284 77840 51300
rect 79058 51414 79066 51486
rect 79672 54090 79682 54246
rect 80328 54262 80384 54368
rect 81638 54358 81824 54368
rect 79716 54090 79728 54246
rect 80328 54242 80340 54262
rect 79672 53568 79728 54090
rect 79672 53396 79682 53568
rect 79716 53396 79728 53568
rect 79672 52874 79728 53396
rect 79672 52702 79682 52874
rect 79716 52702 79728 52874
rect 79672 52180 79728 52702
rect 79672 52008 79682 52180
rect 79716 52008 79728 52180
rect 79672 51486 79728 52008
rect 79672 51446 79682 51486
rect 79024 51298 79058 51314
rect 79662 51314 79682 51446
rect 79716 51402 79728 51486
rect 80326 54090 80340 54242
rect 80374 54210 80384 54262
rect 80998 54262 81032 54278
rect 80374 54090 80382 54210
rect 80326 53568 80382 54090
rect 80326 53396 80340 53568
rect 80374 53396 80382 53568
rect 80326 52874 80382 53396
rect 80326 52702 80340 52874
rect 80374 52702 80382 52874
rect 80326 52180 80382 52702
rect 80326 52008 80340 52180
rect 80374 52008 80382 52180
rect 80326 51486 80382 52008
rect 79716 51314 79722 51402
rect 80326 51398 80340 51486
rect 79662 51204 79722 51314
rect 80374 51398 80382 51486
rect 80986 54090 80998 54200
rect 81638 54262 81714 54358
rect 81032 54090 81042 54200
rect 81638 54180 81656 54262
rect 80986 53568 81042 54090
rect 80986 53396 80998 53568
rect 81032 53396 81042 53568
rect 80986 52874 81042 53396
rect 80986 52702 80998 52874
rect 81032 52702 81042 52874
rect 80986 52180 81042 52702
rect 80986 52008 80998 52180
rect 81032 52008 81042 52180
rect 80986 51486 81042 52008
rect 80986 51356 80998 51486
rect 80340 51298 80374 51314
rect 80990 51314 80998 51356
rect 81032 51444 81042 51486
rect 81640 54090 81656 54180
rect 81690 54180 81714 54262
rect 81896 54182 81910 54918
rect 82086 54182 82128 54936
rect 81690 54090 81696 54180
rect 81896 54108 82128 54182
rect 81640 53568 81696 54090
rect 83272 54065 83303 54099
rect 83337 54065 83399 54099
rect 83433 54065 83495 54099
rect 83529 54065 83591 54099
rect 83625 54065 83687 54099
rect 83721 54065 83783 54099
rect 83817 54065 83879 54099
rect 83913 54065 83975 54099
rect 84009 54065 84071 54099
rect 84105 54065 84167 54099
rect 84201 54065 84263 54099
rect 84297 54065 84359 54099
rect 84393 54065 84455 54099
rect 84489 54065 84551 54099
rect 84585 54065 84647 54099
rect 84681 54065 84743 54099
rect 84777 54065 84839 54099
rect 84873 54065 84935 54099
rect 84969 54065 85031 54099
rect 85065 54065 85127 54099
rect 85161 54065 85223 54099
rect 85257 54065 85319 54099
rect 85353 54065 85415 54099
rect 85449 54065 85511 54099
rect 85545 54065 85607 54099
rect 85641 54065 85703 54099
rect 85737 54065 85799 54099
rect 85833 54065 85895 54099
rect 85929 54065 85991 54099
rect 86025 54065 86087 54099
rect 86121 54065 86183 54099
rect 86217 54065 86279 54099
rect 86313 54065 86344 54099
rect 83398 54003 83516 54009
rect 83398 53969 83404 54003
rect 83438 53969 83476 54003
rect 83510 53969 83516 54003
rect 81640 53396 81656 53568
rect 81690 53396 81696 53568
rect 81640 52874 81696 53396
rect 83294 53943 83360 53959
rect 83294 53909 83310 53943
rect 83344 53909 83360 53943
rect 83294 53851 83360 53909
rect 83294 53817 83310 53851
rect 83344 53817 83360 53851
rect 83294 53773 83360 53817
rect 83398 53947 83516 53969
rect 83398 53913 83466 53947
rect 83500 53913 83516 53947
rect 83398 53847 83516 53913
rect 83398 53813 83466 53847
rect 83500 53813 83516 53847
rect 83552 53995 83840 54029
rect 83552 53773 83586 53995
rect 83294 53757 83586 53773
rect 83294 53739 83536 53757
rect 83294 53434 83348 53739
rect 83520 53723 83536 53739
rect 83570 53723 83586 53757
rect 83448 53640 83450 53698
rect 83384 53621 83450 53640
rect 83520 53689 83586 53723
rect 83520 53655 83536 53689
rect 83570 53655 83586 53689
rect 83520 53639 83586 53655
rect 83622 53943 83672 53959
rect 83656 53909 83672 53943
rect 83622 53851 83672 53909
rect 83656 53817 83672 53851
rect 83622 53698 83672 53817
rect 83720 53942 83770 53959
rect 83720 53908 83736 53942
rect 83720 53836 83770 53908
rect 83806 53906 83840 53995
rect 83876 54003 83942 54009
rect 83876 53969 83882 54003
rect 83916 53976 83942 54003
rect 83876 53942 83892 53969
rect 83926 53942 83942 53976
rect 83978 53995 84326 54029
rect 83978 53906 84012 53995
rect 83806 53872 84012 53906
rect 84048 53942 84082 53959
rect 84188 53950 84254 53959
rect 84188 53916 84204 53950
rect 84238 53916 84254 53950
rect 84188 53908 84254 53916
rect 84048 53836 84082 53908
rect 83720 53802 84082 53836
rect 84118 53852 84162 53868
rect 84118 53818 84123 53852
rect 84157 53818 84162 53852
rect 84118 53802 84162 53818
rect 84048 53766 84082 53802
rect 83811 53710 83919 53766
rect 84048 53732 84092 53766
rect 83622 53692 83727 53698
rect 83622 53658 83687 53692
rect 83721 53658 83727 53692
rect 83622 53652 83727 53658
rect 83811 53676 83827 53710
rect 83861 53676 83919 53710
rect 83384 53587 83400 53621
rect 83434 53587 83450 53621
rect 83384 53553 83450 53587
rect 83384 53519 83400 53553
rect 83434 53519 83450 53553
rect 83384 53503 83450 53519
rect 83622 53467 83676 53652
rect 83811 53642 83919 53676
rect 83811 53608 83827 53642
rect 83861 53608 83919 53642
rect 83811 53592 83919 53608
rect 83294 53400 83314 53434
rect 83294 53367 83348 53400
rect 83384 53434 83574 53467
rect 83384 53400 83470 53434
rect 83504 53400 83574 53434
rect 83384 53381 83574 53400
rect 83384 53347 83390 53381
rect 83424 53347 83462 53381
rect 83496 53347 83534 53381
rect 83568 53347 83574 53381
rect 83610 53434 83676 53467
rect 83610 53400 83626 53434
rect 83660 53400 83676 53434
rect 83610 53367 83676 53400
rect 83712 53500 83830 53517
rect 83712 53466 83764 53500
rect 83798 53466 83830 53500
rect 83885 53498 83919 53592
rect 83955 53673 84021 53689
rect 83955 53639 83971 53673
rect 84005 53639 84021 53673
rect 83955 53606 84021 53639
rect 83955 53550 83970 53606
rect 84020 53550 84021 53606
rect 83712 53381 83830 53466
rect 83384 53341 83574 53347
rect 83712 53347 83718 53381
rect 83752 53347 83790 53381
rect 83824 53347 83830 53381
rect 83885 53394 83919 53460
rect 83955 53430 84021 53550
rect 84058 53533 84092 53732
rect 84128 53698 84162 53802
rect 84198 53768 84232 53908
rect 84292 53877 84326 53995
rect 84362 54003 84552 54009
rect 84362 53969 84368 54003
rect 84402 53969 84440 54003
rect 84474 53969 84512 54003
rect 84546 53969 84552 54003
rect 84362 53961 84552 53969
rect 84362 53927 84502 53961
rect 84536 53927 84552 53961
rect 84362 53913 84552 53927
rect 84588 53995 84794 54029
rect 84588 53877 84622 53995
rect 84292 53868 84622 53877
rect 84268 53852 84622 53868
rect 84268 53818 84284 53852
rect 84318 53843 84622 53852
rect 84658 53950 84724 53959
rect 84658 53916 84674 53950
rect 84708 53916 84724 53950
rect 84318 53818 84334 53843
rect 84268 53804 84334 53818
rect 84658 53807 84724 53916
rect 84760 53923 84794 53995
rect 84830 54003 85020 54019
rect 84830 53969 84836 54003
rect 84870 53998 84908 54003
rect 84880 53969 84908 53998
rect 84942 53969 84980 54003
rect 85014 53969 85020 54003
rect 84830 53964 84846 53969
rect 84880 53964 85020 53969
rect 84830 53959 85020 53964
rect 85158 54003 85208 54019
rect 85192 53969 85208 54003
rect 85158 53928 85208 53969
rect 84760 53889 85122 53923
rect 84370 53773 84724 53807
rect 84986 53819 85002 53853
rect 85036 53819 85052 53853
rect 84370 53768 84404 53773
rect 84198 53734 84404 53768
rect 84986 53737 85052 53819
rect 84128 53692 84333 53698
rect 84128 53658 84167 53692
rect 84201 53667 84333 53692
rect 84201 53658 84283 53667
rect 84128 53652 84283 53658
rect 84267 53633 84283 53652
rect 84317 53633 84333 53667
rect 84267 53599 84333 53633
rect 84267 53565 84283 53599
rect 84317 53565 84333 53599
rect 84267 53553 84333 53565
rect 84370 53597 84404 53734
rect 84440 53736 85052 53737
rect 84440 53702 84456 53736
rect 84490 53703 85052 53736
rect 84490 53702 84506 53703
rect 84440 53668 84506 53702
rect 84440 53634 84456 53668
rect 84490 53634 84506 53668
rect 84440 53633 84506 53634
rect 84593 53633 84609 53667
rect 84643 53633 84964 53667
rect 84370 53563 84844 53597
rect 84878 53563 84894 53597
rect 84058 53500 84112 53533
rect 84370 53517 84404 53563
rect 84930 53527 84964 53633
rect 84058 53466 84062 53500
rect 84096 53466 84112 53500
rect 84058 53433 84112 53466
rect 84202 53500 84404 53517
rect 84202 53466 84218 53500
rect 84252 53483 84404 53500
rect 84440 53493 84964 53527
rect 84252 53466 84268 53483
rect 84202 53433 84268 53466
rect 84440 53394 84474 53493
rect 83885 53360 84474 53394
rect 84704 53437 84894 53457
rect 84704 53403 84844 53437
rect 84878 53403 84894 53437
rect 84704 53381 84894 53403
rect 83712 53341 83830 53347
rect 84704 53347 84710 53381
rect 84744 53347 84782 53381
rect 84816 53347 84854 53381
rect 84888 53347 84894 53381
rect 84704 53341 84894 53347
rect 84930 53355 84964 53493
rect 85000 53533 85052 53703
rect 85088 53763 85122 53889
rect 85192 53894 85208 53928
rect 85158 53853 85208 53894
rect 85192 53837 85208 53853
rect 85369 54003 85559 54009
rect 85369 53969 85375 54003
rect 85409 53969 85447 54003
rect 85481 53969 85519 54003
rect 85553 53969 85559 54003
rect 85369 53870 85559 53969
rect 85726 54003 85905 54009
rect 85760 53969 85798 54003
rect 85832 53969 85870 54003
rect 85904 53969 85905 54003
rect 85192 53819 85333 53837
rect 85158 53803 85333 53819
rect 85369 53836 85479 53870
rect 85513 53836 85559 53870
rect 85369 53803 85559 53836
rect 85640 53870 85690 53903
rect 85640 53836 85656 53870
rect 85726 53883 85905 53969
rect 85726 53849 85812 53883
rect 85846 53849 85905 53883
rect 86027 54003 86216 54015
rect 86027 53969 86032 54003
rect 86066 53969 86104 54003
rect 86138 53999 86176 54003
rect 86150 53969 86176 53999
rect 86210 53969 86216 54003
rect 86027 53965 86116 53969
rect 86150 53965 86216 53969
rect 86027 53919 86216 53965
rect 86027 53885 86116 53919
rect 86150 53885 86216 53919
rect 85726 53845 85905 53849
rect 85941 53853 85991 53869
rect 85640 53809 85690 53836
rect 85975 53819 85991 53853
rect 85088 53695 85122 53729
rect 85088 53619 85122 53661
rect 85197 53739 85263 53755
rect 85197 53705 85213 53739
rect 85247 53705 85263 53739
rect 85299 53739 85333 53803
rect 85640 53775 85841 53809
rect 85299 53705 85721 53739
rect 85755 53705 85771 53739
rect 85197 53692 85263 53705
rect 85197 53658 85223 53692
rect 85257 53658 85263 53692
rect 85197 53655 85263 53658
rect 85088 53603 85322 53619
rect 85088 53585 85281 53603
rect 85265 53569 85281 53585
rect 85315 53569 85322 53603
rect 85265 53535 85322 53569
rect 85000 53517 85066 53533
rect 85000 53483 85016 53517
rect 85050 53483 85066 53517
rect 85000 53425 85066 53483
rect 85000 53391 85016 53425
rect 85050 53391 85066 53425
rect 85158 53517 85224 53533
rect 85158 53483 85174 53517
rect 85208 53483 85224 53517
rect 85265 53501 85281 53535
rect 85315 53501 85322 53535
rect 85265 53485 85322 53501
rect 85158 53425 85224 53483
rect 85358 53425 85392 53705
rect 85807 53669 85841 53775
rect 85433 53664 85841 53669
rect 85433 53630 85449 53664
rect 85483 53635 85841 53664
rect 85483 53630 85499 53635
rect 85433 53596 85499 53630
rect 85433 53562 85449 53596
rect 85483 53562 85499 53596
rect 85433 53557 85499 53562
rect 85563 53565 85579 53599
rect 85613 53565 85629 53599
rect 85563 53531 85629 53565
rect 85563 53521 85579 53531
rect 85158 53391 85174 53425
rect 85208 53391 85392 53425
rect 85428 53497 85579 53521
rect 85613 53497 85629 53531
rect 85428 53487 85629 53497
rect 85428 53355 85462 53487
rect 85796 53467 85841 53635
rect 85941 53753 85991 53819
rect 85975 53719 85991 53753
rect 85941 53669 85991 53719
rect 86027 53837 86216 53885
rect 86027 53803 86116 53837
rect 86150 53803 86216 53837
rect 86027 53757 86216 53803
rect 86027 53723 86116 53757
rect 86150 53723 86216 53757
rect 86027 53707 86216 53723
rect 86252 53999 86319 54015
rect 86252 53965 86272 53999
rect 86306 53965 86319 53999
rect 86252 53919 86319 53965
rect 86252 53885 86272 53919
rect 86306 53885 86319 53919
rect 86252 53837 86319 53885
rect 86252 53803 86272 53837
rect 86306 53803 86319 53837
rect 86252 53757 86319 53803
rect 86252 53723 86272 53757
rect 86306 53723 86319 53757
rect 85941 53653 86216 53669
rect 85941 53619 86166 53653
rect 86200 53619 86216 53653
rect 85941 53603 86216 53619
rect 86252 53630 86319 53723
rect 85941 53567 85983 53603
rect 86252 53586 86270 53630
rect 86316 53586 86319 53630
rect 85917 53534 85983 53567
rect 85917 53500 85933 53534
rect 85967 53500 85983 53534
rect 85917 53467 85983 53500
rect 86019 53551 86209 53567
rect 86019 53517 86112 53551
rect 86146 53517 86209 53551
rect 84930 53321 85462 53355
rect 85498 53434 85688 53451
rect 85498 53400 85514 53434
rect 85548 53400 85688 53434
rect 85498 53381 85688 53400
rect 85498 53347 85504 53381
rect 85538 53347 85576 53381
rect 85610 53347 85648 53381
rect 85682 53347 85688 53381
rect 85796 53434 85862 53467
rect 85796 53400 85812 53434
rect 85846 53400 85862 53434
rect 85796 53367 85862 53400
rect 86019 53451 86209 53517
rect 86019 53417 86112 53451
rect 86146 53417 86209 53451
rect 86019 53381 86209 53417
rect 86252 53551 86319 53586
rect 86252 53517 86268 53551
rect 86302 53517 86319 53551
rect 86252 53451 86319 53517
rect 86252 53417 86268 53451
rect 86302 53417 86319 53451
rect 86252 53401 86319 53417
rect 85498 53341 85688 53347
rect 86019 53347 86025 53381
rect 86059 53347 86097 53381
rect 86131 53347 86169 53381
rect 86203 53347 86209 53381
rect 86019 53341 86209 53347
rect 83272 53251 83303 53285
rect 83337 53251 83399 53285
rect 83433 53251 83495 53285
rect 83529 53251 83591 53285
rect 83625 53251 83687 53285
rect 83721 53251 83783 53285
rect 83817 53251 83879 53285
rect 83913 53251 83975 53285
rect 84009 53251 84071 53285
rect 84105 53251 84167 53285
rect 84201 53251 84263 53285
rect 84297 53251 84359 53285
rect 84393 53251 84455 53285
rect 84489 53251 84551 53285
rect 84585 53251 84647 53285
rect 84681 53251 84743 53285
rect 84777 53251 84839 53285
rect 84873 53251 84935 53285
rect 84969 53251 85031 53285
rect 85065 53251 85127 53285
rect 85161 53251 85223 53285
rect 85257 53251 85319 53285
rect 85353 53251 85415 53285
rect 85449 53251 85511 53285
rect 85545 53251 85607 53285
rect 85641 53251 85703 53285
rect 85737 53251 85799 53285
rect 85833 53251 85895 53285
rect 85929 53251 85991 53285
rect 86025 53251 86087 53285
rect 86121 53251 86183 53285
rect 86217 53251 86279 53285
rect 86313 53251 86344 53285
rect 81640 52702 81656 52874
rect 81690 52702 81696 52874
rect 81640 52180 81696 52702
rect 81640 52008 81656 52180
rect 81690 52008 81696 52180
rect 81640 51486 81696 52008
rect 81032 51314 81050 51444
rect 81640 51360 81656 51486
rect 80990 51208 81050 51314
rect 81690 51360 81696 51486
rect 81656 51298 81690 51314
rect 80990 51204 81148 51208
rect 77140 51190 77298 51194
rect 71948 51142 72008 51148
rect 73276 51140 73336 51148
rect 75812 51128 77298 51190
rect 79662 51142 81148 51204
rect 79662 51136 79722 51142
rect 80990 51134 81050 51142
rect 75812 51122 75872 51128
rect 75934 48690 76256 51128
rect 77140 51120 77200 51128
rect 77322 51022 77690 51054
rect 77322 50826 77348 51022
rect 77656 50826 77690 51022
rect 77322 50798 77690 50826
rect 58938 46342 66184 46504
rect 38714 45148 42794 45178
rect 24024 44998 25442 45070
rect 24024 44696 24240 44998
rect 25328 44696 25442 44998
rect 24024 44582 25442 44696
rect 38714 44424 38946 45148
rect 42360 44424 42794 45148
rect 38714 44308 42794 44424
rect 49454 43936 50070 44004
rect 11016 43736 11290 43774
rect 1910 43330 2046 43626
rect 11016 43606 11050 43736
rect 11240 43606 11290 43736
rect 11016 43566 11290 43606
rect 7240 43362 7376 43390
rect 4048 43330 4116 43346
rect 6172 43338 8648 43362
rect 10562 43338 10630 43354
rect 11078 43338 11192 43566
rect 12686 43352 12754 43370
rect 14964 43352 15032 43356
rect 12624 43346 15426 43352
rect 17068 43346 17136 43362
rect 19192 43346 19260 43378
rect 12624 43340 19260 43346
rect 20254 43340 20338 43350
rect 12624 43338 20338 43340
rect 6172 43330 20338 43338
rect 1910 43320 20338 43330
rect 1806 43256 20338 43320
rect 1806 43246 19116 43256
rect 1806 43240 15426 43246
rect 1806 43230 6096 43240
rect 6164 43238 15426 43240
rect 1910 43052 2046 43230
rect 1910 42760 1958 43052
rect 1992 42760 2046 43052
rect 3016 43052 3050 43068
rect 1910 41958 2046 42760
rect 1910 41666 1958 41958
rect 1992 41666 2046 41958
rect 1304 41518 1454 41644
rect 1304 40322 1326 41518
rect 1420 40322 1454 41518
rect 1304 39998 1454 40322
rect 1910 40864 2046 41666
rect 1910 40572 1958 40864
rect 1992 40572 2046 40864
rect 1910 39770 2046 40572
rect 1910 39478 1958 39770
rect 1992 39478 2046 39770
rect 1910 38676 2046 39478
rect 1910 38384 1958 38676
rect 1992 38384 2046 38676
rect 3012 42760 3016 42958
rect 4048 43052 4116 43230
rect 6164 43116 8648 43238
rect 4048 42964 4074 43052
rect 3050 42760 3058 42958
rect 3012 41958 3058 42760
rect 3012 41666 3016 41958
rect 3050 41666 3058 41958
rect 3012 40864 3058 41666
rect 3012 40572 3016 40864
rect 3050 40572 3058 40864
rect 3012 39770 3058 40572
rect 3012 39478 3016 39770
rect 3050 39478 3058 39770
rect 3012 38676 3058 39478
rect 3012 38596 3016 38676
rect 1910 37514 2046 38384
rect 2996 38384 3016 38484
rect 3050 38596 3058 38676
rect 4064 42760 4074 42964
rect 4108 43016 4116 43052
rect 5132 43052 5166 43068
rect 4108 42964 4122 43016
rect 4108 42760 4110 42964
rect 4064 41958 4110 42760
rect 4064 41666 4074 41958
rect 4108 41666 4110 41958
rect 4064 40864 4110 41666
rect 4064 40572 4074 40864
rect 4108 40572 4110 40864
rect 4064 39770 4110 40572
rect 4064 39478 4074 39770
rect 4108 39478 4110 39770
rect 4064 38676 4110 39478
rect 4064 38618 4074 38676
rect 3050 38384 3078 38484
rect 2996 38274 3078 38384
rect 4108 38618 4110 38676
rect 6164 43052 6248 43116
rect 5166 42760 5178 42964
rect 6164 42960 6190 43052
rect 5132 41958 5178 42760
rect 5166 41666 5178 41958
rect 5132 40864 5178 41666
rect 5166 40572 5178 40864
rect 5132 39770 5178 40572
rect 5166 39478 5178 39770
rect 5132 38676 5178 39478
rect 4074 38368 4108 38384
rect 5122 38384 5132 38456
rect 5166 38602 5178 38676
rect 6184 42760 6190 42960
rect 6224 42960 6248 43052
rect 7240 43052 7376 43116
rect 6224 42760 6230 42960
rect 6184 41958 6230 42760
rect 6184 41666 6190 41958
rect 6224 41666 6230 41958
rect 6184 40864 6230 41666
rect 6184 40572 6190 40864
rect 6224 40572 6230 40864
rect 6184 39770 6230 40572
rect 6184 39478 6190 39770
rect 6224 39478 6230 39770
rect 6184 38676 6230 39478
rect 6184 38646 6190 38676
rect 5166 38384 5204 38456
rect 5122 38274 5204 38384
rect 6224 38646 6230 38676
rect 7240 42760 7248 43052
rect 7282 42760 7376 43052
rect 7240 41958 7376 42760
rect 7240 41666 7248 41958
rect 7282 41666 7376 41958
rect 7240 40864 7376 41666
rect 8436 43060 8572 43116
rect 8436 42768 8472 43060
rect 8506 42768 8572 43060
rect 9530 43060 9564 43076
rect 8436 41966 8572 42768
rect 8436 41674 8472 41966
rect 8506 41674 8572 41966
rect 7240 40572 7248 40864
rect 7282 40572 7376 40864
rect 7240 39770 7376 40572
rect 7818 41526 7968 41652
rect 7818 40330 7840 41526
rect 7934 40330 7968 41526
rect 7818 40006 7968 40330
rect 8436 40872 8572 41674
rect 8436 40580 8472 40872
rect 8506 40580 8572 40872
rect 7240 39478 7248 39770
rect 7282 39478 7376 39770
rect 7240 38676 7376 39478
rect 7240 38478 7248 38676
rect 6190 38368 6224 38384
rect 7224 38384 7248 38478
rect 7282 38384 7376 38676
rect 7224 38274 7376 38384
rect 8436 39778 8572 40580
rect 8436 39486 8472 39778
rect 8506 39486 8572 39778
rect 8436 38684 8572 39486
rect 8436 38392 8472 38684
rect 8506 38392 8572 38684
rect 9526 42768 9530 42966
rect 10562 43060 10630 43238
rect 12578 43224 15426 43238
rect 10562 42972 10588 43060
rect 9564 42768 9572 42966
rect 9526 41966 9572 42768
rect 9526 41674 9530 41966
rect 9564 41674 9572 41966
rect 9526 40872 9572 41674
rect 9526 40580 9530 40872
rect 9564 40580 9572 40872
rect 9526 39778 9572 40580
rect 9526 39486 9530 39778
rect 9564 39486 9572 39778
rect 9526 38684 9572 39486
rect 9526 38604 9530 38684
rect 2996 38184 7446 38274
rect 3008 38178 7446 38184
rect 5122 38156 5204 38178
rect 4048 37514 4116 37530
rect 6172 37514 6240 37546
rect 1910 37504 6240 37514
rect 1806 37460 6240 37504
rect 1806 37424 6248 37460
rect 1806 37414 6096 37424
rect 1910 37236 2046 37414
rect 1910 36944 1958 37236
rect 1992 36944 2046 37236
rect 3016 37236 3050 37252
rect 1910 36142 2046 36944
rect 1910 35850 1958 36142
rect 1992 35850 2046 36142
rect 1304 35702 1454 35828
rect 1304 34506 1326 35702
rect 1420 34506 1454 35702
rect 1304 34182 1454 34506
rect 1910 35048 2046 35850
rect 1910 34756 1958 35048
rect 1992 34756 2046 35048
rect 1910 33954 2046 34756
rect 1910 33662 1958 33954
rect 1992 33662 2046 33954
rect 1910 32860 2046 33662
rect 1910 32568 1958 32860
rect 1992 32568 2046 32860
rect 3012 36944 3016 37142
rect 4048 37236 4116 37414
rect 4048 37148 4074 37236
rect 3050 36944 3058 37142
rect 3012 36142 3058 36944
rect 3012 35850 3016 36142
rect 3050 35850 3058 36142
rect 3012 35048 3058 35850
rect 3012 34756 3016 35048
rect 3050 34756 3058 35048
rect 3012 33954 3058 34756
rect 3012 33662 3016 33954
rect 3050 33662 3058 33954
rect 3012 32860 3058 33662
rect 3012 32780 3016 32860
rect 1910 31680 2046 32568
rect 2996 32568 3016 32668
rect 3050 32780 3058 32860
rect 4064 36944 4074 37148
rect 4108 37200 4116 37236
rect 5132 37236 5166 37252
rect 4108 37148 4122 37200
rect 4108 36944 4110 37148
rect 4064 36142 4110 36944
rect 4064 35850 4074 36142
rect 4108 35850 4110 36142
rect 4064 35048 4110 35850
rect 4064 34756 4074 35048
rect 4108 34756 4110 35048
rect 4064 33954 4110 34756
rect 4064 33662 4074 33954
rect 4108 33662 4110 33954
rect 4064 32860 4110 33662
rect 4064 32802 4074 32860
rect 3050 32568 3078 32668
rect 2996 32458 3078 32568
rect 4108 32802 4110 32860
rect 6164 37236 6248 37424
rect 5166 36944 5178 37148
rect 6164 37144 6190 37236
rect 5132 36142 5178 36944
rect 5166 35850 5178 36142
rect 5132 35048 5178 35850
rect 5166 34756 5178 35048
rect 5132 33954 5178 34756
rect 5166 33662 5178 33954
rect 5132 32860 5178 33662
rect 4074 32552 4108 32568
rect 5122 32568 5132 32640
rect 5166 32786 5178 32860
rect 6184 36944 6190 37144
rect 6224 37144 6248 37236
rect 7240 37236 7376 38178
rect 8436 37522 8572 38392
rect 9510 38392 9530 38492
rect 9564 38604 9572 38684
rect 10578 42768 10588 42972
rect 10622 43024 10630 43060
rect 11646 43060 11680 43076
rect 10622 42972 10636 43024
rect 10622 42768 10624 42972
rect 10578 41966 10624 42768
rect 10578 41674 10588 41966
rect 10622 41674 10624 41966
rect 10578 40872 10624 41674
rect 10578 40580 10588 40872
rect 10622 40580 10624 40872
rect 10578 39778 10624 40580
rect 10578 39486 10588 39778
rect 10622 39486 10624 39778
rect 10578 38684 10624 39486
rect 10578 38626 10588 38684
rect 9564 38392 9592 38492
rect 9510 38282 9592 38392
rect 10622 38626 10624 38684
rect 12678 43060 12762 43224
rect 11680 42768 11692 42972
rect 12678 42968 12704 43060
rect 11646 41966 11692 42768
rect 11680 41674 11692 41966
rect 11646 40872 11692 41674
rect 11680 40580 11692 40872
rect 11646 39778 11692 40580
rect 11680 39486 11692 39778
rect 11646 38684 11692 39486
rect 10588 38376 10622 38392
rect 11636 38392 11646 38464
rect 11680 38610 11692 38684
rect 12698 42768 12704 42968
rect 12738 42968 12762 43060
rect 13746 43060 13888 43224
rect 13746 43022 13762 43060
rect 13742 42972 13762 43022
rect 12738 42768 12744 42968
rect 12698 41966 12744 42768
rect 12698 41674 12704 41966
rect 12738 41674 12744 41966
rect 12698 40872 12744 41674
rect 12698 40580 12704 40872
rect 12738 40580 12744 40872
rect 12698 39778 12744 40580
rect 12698 39486 12704 39778
rect 12738 39486 12744 39778
rect 12698 38684 12744 39486
rect 12698 38654 12704 38684
rect 11680 38392 11718 38464
rect 11636 38282 11718 38392
rect 12738 38654 12744 38684
rect 13754 42768 13762 42972
rect 13796 43006 13888 43060
rect 14940 43068 15032 43224
rect 13796 42768 13874 43006
rect 13754 41966 13874 42768
rect 13754 41674 13762 41966
rect 13796 41674 13874 41966
rect 13754 40872 13874 41674
rect 14940 42776 14978 43068
rect 15012 42966 15032 43068
rect 16036 43068 16070 43084
rect 15012 42776 15028 42966
rect 14940 41974 15028 42776
rect 14940 41682 14978 41974
rect 15012 41682 15028 41974
rect 13754 40580 13762 40872
rect 13796 40580 13874 40872
rect 13754 39778 13874 40580
rect 14324 41534 14474 41660
rect 14324 40338 14346 41534
rect 14440 40338 14474 41534
rect 14324 40014 14474 40338
rect 14940 40880 15028 41682
rect 14940 40588 14978 40880
rect 15012 40588 15028 40880
rect 13754 39486 13762 39778
rect 13796 39486 13874 39778
rect 13754 38684 13874 39486
rect 13754 38626 13762 38684
rect 12704 38376 12738 38392
rect 13738 38392 13762 38486
rect 13796 38392 13874 38684
rect 13738 38282 13874 38392
rect 14940 39786 15028 40588
rect 14940 39494 14978 39786
rect 15012 39494 15028 39786
rect 14940 38692 15028 39494
rect 14940 38400 14978 38692
rect 15012 38400 15028 38692
rect 16032 42776 16036 42974
rect 17068 43068 17136 43246
rect 19182 43206 20338 43256
rect 17068 42980 17094 43068
rect 16070 42776 16078 42974
rect 16032 41974 16078 42776
rect 16032 41682 16036 41974
rect 16070 41682 16078 41974
rect 16032 40880 16078 41682
rect 16032 40588 16036 40880
rect 16070 40588 16078 40880
rect 16032 39786 16078 40588
rect 16032 39494 16036 39786
rect 16070 39494 16078 39786
rect 16032 38692 16078 39494
rect 16032 38612 16036 38692
rect 9510 38192 13960 38282
rect 9522 38186 13960 38192
rect 11636 38164 11718 38186
rect 10562 37522 10630 37538
rect 12686 37522 12754 37554
rect 8436 37512 12754 37522
rect 8320 37468 12754 37512
rect 8320 37432 12762 37468
rect 8320 37422 12610 37432
rect 6224 36944 6230 37144
rect 6184 36142 6230 36944
rect 6184 35850 6190 36142
rect 6224 35850 6230 36142
rect 6184 35048 6230 35850
rect 6184 34756 6190 35048
rect 6224 34756 6230 35048
rect 6184 33954 6230 34756
rect 6184 33662 6190 33954
rect 6224 33662 6230 33954
rect 6184 32860 6230 33662
rect 6184 32830 6190 32860
rect 5166 32568 5204 32640
rect 5122 32458 5204 32568
rect 6224 32830 6230 32860
rect 7240 36944 7248 37236
rect 7282 36944 7376 37236
rect 7240 36142 7376 36944
rect 7240 35850 7248 36142
rect 7282 35850 7376 36142
rect 7240 35048 7376 35850
rect 8436 37244 8572 37422
rect 8436 36952 8472 37244
rect 8506 36952 8572 37244
rect 9530 37244 9564 37260
rect 8436 36150 8572 36952
rect 8436 35858 8472 36150
rect 8506 35858 8572 36150
rect 7240 34756 7248 35048
rect 7282 34756 7376 35048
rect 7240 33954 7376 34756
rect 7818 35710 7968 35836
rect 7818 34514 7840 35710
rect 7934 34514 7968 35710
rect 7818 34190 7968 34514
rect 8436 35056 8572 35858
rect 8436 34764 8472 35056
rect 8506 34764 8572 35056
rect 7240 33662 7248 33954
rect 7282 33662 7376 33954
rect 7240 32860 7376 33662
rect 7240 32662 7248 32860
rect 6190 32552 6224 32568
rect 7224 32568 7248 32662
rect 7282 32568 7376 32860
rect 7224 32458 7376 32568
rect 8436 33962 8572 34764
rect 8436 33670 8472 33962
rect 8506 33670 8572 33962
rect 8436 32868 8572 33670
rect 8436 32576 8472 32868
rect 8506 32576 8572 32868
rect 9526 36952 9530 37150
rect 10562 37244 10630 37422
rect 10562 37156 10588 37244
rect 9564 36952 9572 37150
rect 9526 36150 9572 36952
rect 9526 35858 9530 36150
rect 9564 35858 9572 36150
rect 9526 35056 9572 35858
rect 9526 34764 9530 35056
rect 9564 34764 9572 35056
rect 9526 33962 9572 34764
rect 9526 33670 9530 33962
rect 9564 33670 9572 33962
rect 9526 32868 9572 33670
rect 9526 32788 9530 32868
rect 2996 32368 7446 32458
rect 3008 32362 7446 32368
rect 5122 32340 5204 32362
rect 4048 31680 4116 31696
rect 6172 31680 6240 31712
rect 1910 31670 6240 31680
rect 1806 31626 6240 31670
rect 1806 31590 6248 31626
rect 1806 31580 6096 31590
rect 1910 31402 2046 31580
rect 1910 31110 1958 31402
rect 1992 31110 2046 31402
rect 3016 31402 3050 31418
rect 1910 30308 2046 31110
rect 1910 30016 1958 30308
rect 1992 30016 2046 30308
rect 1304 29868 1454 29994
rect 1304 28672 1326 29868
rect 1420 28672 1454 29868
rect 1304 28348 1454 28672
rect 1910 29214 2046 30016
rect 1910 28922 1958 29214
rect 1992 28922 2046 29214
rect 1910 28120 2046 28922
rect 1910 27828 1958 28120
rect 1992 27828 2046 28120
rect 1910 27026 2046 27828
rect 1910 26734 1958 27026
rect 1992 26734 2046 27026
rect 3012 31110 3016 31308
rect 4048 31402 4116 31580
rect 4048 31314 4074 31402
rect 3050 31110 3058 31308
rect 3012 30308 3058 31110
rect 3012 30016 3016 30308
rect 3050 30016 3058 30308
rect 3012 29214 3058 30016
rect 3012 28922 3016 29214
rect 3050 28922 3058 29214
rect 3012 28120 3058 28922
rect 3012 27828 3016 28120
rect 3050 27828 3058 28120
rect 3012 27026 3058 27828
rect 3012 26946 3016 27026
rect 1910 25844 2046 26734
rect 2996 26734 3016 26834
rect 3050 26946 3058 27026
rect 4064 31110 4074 31314
rect 4108 31366 4116 31402
rect 5132 31402 5166 31418
rect 4108 31314 4122 31366
rect 4108 31110 4110 31314
rect 4064 30308 4110 31110
rect 4064 30016 4074 30308
rect 4108 30016 4110 30308
rect 4064 29214 4110 30016
rect 4064 28922 4074 29214
rect 4108 28922 4110 29214
rect 4064 28120 4110 28922
rect 4064 27828 4074 28120
rect 4108 27828 4110 28120
rect 4064 27026 4110 27828
rect 4064 26968 4074 27026
rect 3050 26734 3078 26834
rect 2996 26624 3078 26734
rect 4108 26968 4110 27026
rect 6164 31402 6248 31590
rect 5166 31110 5178 31314
rect 6164 31310 6190 31402
rect 5132 30308 5178 31110
rect 5166 30016 5178 30308
rect 5132 29214 5178 30016
rect 5166 28922 5178 29214
rect 5132 28120 5178 28922
rect 5166 27828 5178 28120
rect 5132 27026 5178 27828
rect 4074 26718 4108 26734
rect 5122 26734 5132 26806
rect 5166 26952 5178 27026
rect 6184 31110 6190 31310
rect 6224 31310 6248 31402
rect 7240 31402 7376 32362
rect 8436 31688 8572 32576
rect 9510 32576 9530 32676
rect 9564 32788 9572 32868
rect 10578 36952 10588 37156
rect 10622 37208 10630 37244
rect 11646 37244 11680 37260
rect 10622 37156 10636 37208
rect 10622 36952 10624 37156
rect 10578 36150 10624 36952
rect 10578 35858 10588 36150
rect 10622 35858 10624 36150
rect 10578 35056 10624 35858
rect 10578 34764 10588 35056
rect 10622 34764 10624 35056
rect 10578 33962 10624 34764
rect 10578 33670 10588 33962
rect 10622 33670 10624 33962
rect 10578 32868 10624 33670
rect 10578 32810 10588 32868
rect 9564 32576 9592 32676
rect 9510 32466 9592 32576
rect 10622 32810 10624 32868
rect 12678 37244 12762 37432
rect 13768 37260 13874 38186
rect 14940 37540 15028 38400
rect 16016 38400 16036 38500
rect 16070 38612 16078 38692
rect 17084 42776 17094 42980
rect 17128 43032 17136 43068
rect 18152 43068 18186 43084
rect 17128 42980 17142 43032
rect 17128 42776 17130 42980
rect 17084 41974 17130 42776
rect 17084 41682 17094 41974
rect 17128 41682 17130 41974
rect 17084 40880 17130 41682
rect 17084 40588 17094 40880
rect 17128 40588 17130 40880
rect 17084 39786 17130 40588
rect 17084 39494 17094 39786
rect 17128 39494 17130 39786
rect 17084 38692 17130 39494
rect 17084 38634 17094 38692
rect 16070 38400 16098 38500
rect 16016 38290 16098 38400
rect 17128 38634 17130 38692
rect 19184 43068 19268 43206
rect 18186 42776 18198 42980
rect 19184 42976 19210 43068
rect 18152 41974 18198 42776
rect 18186 41682 18198 41974
rect 18152 40880 18198 41682
rect 18186 40588 18198 40880
rect 18152 39786 18198 40588
rect 18186 39494 18198 39786
rect 18152 38692 18198 39494
rect 17094 38384 17128 38400
rect 18142 38400 18152 38472
rect 18186 38618 18198 38692
rect 19204 42776 19210 42976
rect 19244 42976 19268 43068
rect 20242 43068 20338 43206
rect 20942 43320 21394 43634
rect 21454 43330 21522 43340
rect 23558 43330 23626 43346
rect 25682 43332 25750 43362
rect 27976 43346 28044 43356
rect 30080 43346 30148 43362
rect 32204 43354 32272 43378
rect 34486 43354 34554 43362
rect 34612 43354 34872 43372
rect 32170 43352 35080 43354
rect 36590 43352 36658 43368
rect 38714 43352 38782 43384
rect 32170 43346 38782 43352
rect 27976 43344 38782 43346
rect 27976 43336 38792 43344
rect 27838 43332 38792 43336
rect 25660 43330 38792 43332
rect 21454 43320 38792 43330
rect 20942 43256 38792 43320
rect 20942 43246 32128 43256
rect 32170 43252 38792 43256
rect 20942 43240 28240 43246
rect 20942 43230 25606 43240
rect 20942 43074 21394 43230
rect 19244 42776 19250 42976
rect 19204 41974 19250 42776
rect 19204 41682 19210 41974
rect 19244 41682 19250 41974
rect 19204 40880 19250 41682
rect 19204 40588 19210 40880
rect 19244 40588 19250 40880
rect 19204 39786 19250 40588
rect 19204 39494 19210 39786
rect 19244 39494 19250 39786
rect 19204 38692 19250 39494
rect 19204 38662 19210 38692
rect 18186 38400 18224 38472
rect 18142 38290 18224 38400
rect 19244 38662 19250 38692
rect 20242 42776 20268 43068
rect 20302 42986 20338 43068
rect 21454 43052 21522 43230
rect 20302 42776 20336 42986
rect 20242 41974 20336 42776
rect 20242 41682 20268 41974
rect 20302 41682 20336 41974
rect 20242 40880 20336 41682
rect 21454 42760 21468 43052
rect 21502 42950 21522 43052
rect 22526 43052 22560 43068
rect 21454 42744 21502 42760
rect 22522 42760 22526 42958
rect 23558 43052 23626 43230
rect 25660 43194 28240 43240
rect 23558 42964 23584 43052
rect 22560 42760 22568 42958
rect 21454 41974 21500 42744
rect 21454 41958 21502 41974
rect 21454 41666 21468 41958
rect 21454 41650 21502 41666
rect 22522 41958 22568 42760
rect 22522 41666 22526 41958
rect 22560 41666 22568 41958
rect 20242 40588 20268 40880
rect 20302 40588 20336 40880
rect 20242 39786 20336 40588
rect 20814 41518 20964 41644
rect 20814 40322 20836 41518
rect 20930 40322 20964 41518
rect 20814 39998 20964 40322
rect 21454 40880 21500 41650
rect 21454 40864 21502 40880
rect 21454 40572 21468 40864
rect 21454 40556 21502 40572
rect 22522 40864 22568 41666
rect 22522 40572 22526 40864
rect 22560 40572 22568 40864
rect 20242 39494 20268 39786
rect 20302 39494 20336 39786
rect 20242 38692 20336 39494
rect 21454 39786 21500 40556
rect 21454 39770 21502 39786
rect 21454 39478 21468 39770
rect 21454 39462 21502 39478
rect 22522 39770 22568 40572
rect 22522 39478 22526 39770
rect 22560 39478 22568 39770
rect 21454 38716 21500 39462
rect 19210 38384 19244 38400
rect 20242 38400 20268 38692
rect 20302 38400 20336 38692
rect 20242 38290 20336 38400
rect 21426 38676 21558 38716
rect 21426 38384 21468 38676
rect 21502 38384 21558 38676
rect 22522 38676 22568 39478
rect 22522 38596 22526 38676
rect 16016 38200 20466 38290
rect 16028 38194 20466 38200
rect 18142 38172 18224 38194
rect 14940 37530 15032 37540
rect 17068 37530 17136 37546
rect 19192 37530 19260 37562
rect 14940 37520 19260 37530
rect 14826 37476 19260 37520
rect 14826 37440 19268 37476
rect 14826 37430 19116 37440
rect 11680 36952 11692 37156
rect 12678 37152 12704 37244
rect 11646 36150 11692 36952
rect 11680 35858 11692 36150
rect 11646 35056 11692 35858
rect 11680 34764 11692 35056
rect 11646 33962 11692 34764
rect 11680 33670 11692 33962
rect 11646 32868 11692 33670
rect 10588 32560 10622 32576
rect 11636 32576 11646 32648
rect 11680 32794 11692 32868
rect 12698 36952 12704 37152
rect 12738 37152 12762 37244
rect 13762 37244 13874 37260
rect 12738 36952 12744 37152
rect 12698 36150 12744 36952
rect 12698 35858 12704 36150
rect 12738 35858 12744 36150
rect 12698 35056 12744 35858
rect 12698 34764 12704 35056
rect 12738 34764 12744 35056
rect 12698 33962 12744 34764
rect 12698 33670 12704 33962
rect 12738 33670 12744 33962
rect 12698 32868 12744 33670
rect 12698 32838 12704 32868
rect 11680 32576 11718 32648
rect 11636 32466 11718 32576
rect 12738 32838 12744 32868
rect 13754 36952 13762 37172
rect 13796 36952 13874 37244
rect 13754 36150 13874 36952
rect 13754 35858 13762 36150
rect 13796 35858 13874 36150
rect 13754 35056 13874 35858
rect 14940 37252 15032 37430
rect 14940 36960 14978 37252
rect 15012 37150 15032 37252
rect 16036 37252 16070 37268
rect 15012 36960 15028 37150
rect 14940 36158 15028 36960
rect 14940 35866 14978 36158
rect 15012 35866 15028 36158
rect 13754 34764 13762 35056
rect 13796 34764 13874 35056
rect 13754 33962 13874 34764
rect 14324 35718 14474 35844
rect 14324 34522 14346 35718
rect 14440 34522 14474 35718
rect 14324 34198 14474 34522
rect 14940 35064 15028 35866
rect 14940 34772 14978 35064
rect 15012 34772 15028 35064
rect 13754 33670 13762 33962
rect 13796 33670 13874 33962
rect 13754 32868 13874 33670
rect 13754 32810 13762 32868
rect 12704 32560 12738 32576
rect 13738 32576 13762 32670
rect 13796 32576 13874 32868
rect 13738 32466 13874 32576
rect 14940 33970 15028 34772
rect 14940 33678 14978 33970
rect 15012 33678 15028 33970
rect 14940 32876 15028 33678
rect 14940 32584 14978 32876
rect 15012 32584 15028 32876
rect 16032 36960 16036 37158
rect 17068 37252 17136 37430
rect 17068 37164 17094 37252
rect 16070 36960 16078 37158
rect 16032 36158 16078 36960
rect 16032 35866 16036 36158
rect 16070 35866 16078 36158
rect 16032 35064 16078 35866
rect 16032 34772 16036 35064
rect 16070 34772 16078 35064
rect 16032 33970 16078 34772
rect 16032 33678 16036 33970
rect 16070 33678 16078 33970
rect 16032 32876 16078 33678
rect 16032 32796 16036 32876
rect 9510 32376 13960 32466
rect 9522 32370 13960 32376
rect 11636 32348 11718 32370
rect 10562 31688 10630 31704
rect 12686 31688 12754 31720
rect 8436 31678 12754 31688
rect 8320 31634 12754 31678
rect 8320 31598 12762 31634
rect 8320 31588 12610 31598
rect 6224 31110 6230 31310
rect 6184 30308 6230 31110
rect 6184 30016 6190 30308
rect 6224 30016 6230 30308
rect 6184 29214 6230 30016
rect 6184 28922 6190 29214
rect 6224 28922 6230 29214
rect 6184 28120 6230 28922
rect 6184 27828 6190 28120
rect 6224 27828 6230 28120
rect 6184 27026 6230 27828
rect 6184 26996 6190 27026
rect 5166 26734 5204 26806
rect 5122 26624 5204 26734
rect 6224 26996 6230 27026
rect 7240 31110 7248 31402
rect 7282 31110 7376 31402
rect 7240 30308 7376 31110
rect 7240 30016 7248 30308
rect 7282 30016 7376 30308
rect 7240 29214 7376 30016
rect 8436 31410 8572 31588
rect 8436 31118 8472 31410
rect 8506 31118 8572 31410
rect 9530 31410 9564 31426
rect 8436 30316 8572 31118
rect 8436 30024 8472 30316
rect 8506 30024 8572 30316
rect 7240 28922 7248 29214
rect 7282 28922 7376 29214
rect 7240 28120 7376 28922
rect 7818 29876 7968 30002
rect 7818 28680 7840 29876
rect 7934 28680 7968 29876
rect 7818 28356 7968 28680
rect 8436 29222 8572 30024
rect 8436 28930 8472 29222
rect 8506 28930 8572 29222
rect 7240 27828 7248 28120
rect 7282 27828 7376 28120
rect 7240 27026 7376 27828
rect 7240 26828 7248 27026
rect 6190 26718 6224 26734
rect 7224 26734 7248 26828
rect 7282 26734 7376 27026
rect 7224 26624 7376 26734
rect 8436 28128 8572 28930
rect 8436 27836 8472 28128
rect 8506 27836 8572 28128
rect 8436 27034 8572 27836
rect 8436 26742 8472 27034
rect 8506 26742 8572 27034
rect 9526 31118 9530 31316
rect 10562 31410 10630 31588
rect 10562 31322 10588 31410
rect 9564 31118 9572 31316
rect 9526 30316 9572 31118
rect 9526 30024 9530 30316
rect 9564 30024 9572 30316
rect 9526 29222 9572 30024
rect 9526 28930 9530 29222
rect 9564 28930 9572 29222
rect 9526 28128 9572 28930
rect 9526 27836 9530 28128
rect 9564 27836 9572 28128
rect 9526 27034 9572 27836
rect 9526 26954 9530 27034
rect 2996 26534 7446 26624
rect 3008 26528 7446 26534
rect 5122 26506 5204 26528
rect 4048 25844 4116 25860
rect 6172 25844 6240 25876
rect 1910 25834 6240 25844
rect 1806 25790 6240 25834
rect 1806 25754 6248 25790
rect 1806 25744 6096 25754
rect 1910 25566 2046 25744
rect 1910 25274 1958 25566
rect 1992 25274 2046 25566
rect 3016 25566 3050 25582
rect 1910 24472 2046 25274
rect 1910 24180 1958 24472
rect 1992 24180 2046 24472
rect 1304 24032 1454 24158
rect 1304 22836 1326 24032
rect 1420 22836 1454 24032
rect 1304 22512 1454 22836
rect 1910 23378 2046 24180
rect 1910 23086 1958 23378
rect 1992 23086 2046 23378
rect 1910 22284 2046 23086
rect 1910 21992 1958 22284
rect 1992 21992 2046 22284
rect 1910 21190 2046 21992
rect 1910 20898 1958 21190
rect 1992 20898 2046 21190
rect 3012 25274 3016 25472
rect 4048 25566 4116 25744
rect 4048 25478 4074 25566
rect 3050 25274 3058 25472
rect 3012 24472 3058 25274
rect 3012 24180 3016 24472
rect 3050 24180 3058 24472
rect 3012 23378 3058 24180
rect 3012 23086 3016 23378
rect 3050 23086 3058 23378
rect 3012 22284 3058 23086
rect 3012 21992 3016 22284
rect 3050 21992 3058 22284
rect 3012 21190 3058 21992
rect 3012 21110 3016 21190
rect 1910 19980 2046 20898
rect 2996 20898 3016 20998
rect 3050 21110 3058 21190
rect 4064 25274 4074 25478
rect 4108 25530 4116 25566
rect 5132 25566 5166 25582
rect 4108 25478 4122 25530
rect 4108 25274 4110 25478
rect 4064 24472 4110 25274
rect 4064 24180 4074 24472
rect 4108 24180 4110 24472
rect 4064 23378 4110 24180
rect 4064 23086 4074 23378
rect 4108 23086 4110 23378
rect 4064 22284 4110 23086
rect 4064 21992 4074 22284
rect 4108 21992 4110 22284
rect 4064 21190 4110 21992
rect 4064 21132 4074 21190
rect 3050 20898 3078 20998
rect 2996 20788 3078 20898
rect 4108 21132 4110 21190
rect 6164 25566 6248 25754
rect 5166 25274 5178 25478
rect 6164 25474 6190 25566
rect 5132 24472 5178 25274
rect 5166 24180 5178 24472
rect 5132 23378 5178 24180
rect 5166 23086 5178 23378
rect 5132 22284 5178 23086
rect 5166 21992 5178 22284
rect 5132 21190 5178 21992
rect 4074 20882 4108 20898
rect 5122 20898 5132 20970
rect 5166 21116 5178 21190
rect 6184 25274 6190 25474
rect 6224 25474 6248 25566
rect 7240 25566 7376 26528
rect 8436 25852 8572 26742
rect 9510 26742 9530 26842
rect 9564 26954 9572 27034
rect 10578 31118 10588 31322
rect 10622 31374 10630 31410
rect 11646 31410 11680 31426
rect 10622 31322 10636 31374
rect 10622 31118 10624 31322
rect 10578 30316 10624 31118
rect 10578 30024 10588 30316
rect 10622 30024 10624 30316
rect 10578 29222 10624 30024
rect 10578 28930 10588 29222
rect 10622 28930 10624 29222
rect 10578 28128 10624 28930
rect 10578 27836 10588 28128
rect 10622 27836 10624 28128
rect 10578 27034 10624 27836
rect 10578 26976 10588 27034
rect 9564 26742 9592 26842
rect 9510 26632 9592 26742
rect 10622 26976 10624 27034
rect 12678 31410 12762 31598
rect 13768 31426 13874 32370
rect 14940 31706 15028 32584
rect 16016 32584 16036 32684
rect 16070 32796 16078 32876
rect 17084 36960 17094 37164
rect 17128 37216 17136 37252
rect 18152 37252 18186 37268
rect 17128 37164 17142 37216
rect 17128 36960 17130 37164
rect 17084 36158 17130 36960
rect 17084 35866 17094 36158
rect 17128 35866 17130 36158
rect 17084 35064 17130 35866
rect 17084 34772 17094 35064
rect 17128 34772 17130 35064
rect 17084 33970 17130 34772
rect 17084 33678 17094 33970
rect 17128 33678 17130 33970
rect 17084 32876 17130 33678
rect 17084 32818 17094 32876
rect 16070 32584 16098 32684
rect 16016 32474 16098 32584
rect 17128 32818 17130 32876
rect 19184 37252 19268 37440
rect 18186 36960 18198 37164
rect 19184 37160 19210 37252
rect 18152 36158 18198 36960
rect 18186 35866 18198 36158
rect 18152 35064 18198 35866
rect 18186 34772 18198 35064
rect 18152 33970 18198 34772
rect 18186 33678 18198 33970
rect 18152 32876 18198 33678
rect 17094 32568 17128 32584
rect 18142 32584 18152 32656
rect 18186 32802 18198 32876
rect 19204 36960 19210 37160
rect 19244 37160 19268 37252
rect 20242 37252 20336 38194
rect 21426 37514 21558 38384
rect 22506 38384 22526 38484
rect 22560 38596 22568 38676
rect 23574 42760 23584 42964
rect 23618 43016 23626 43052
rect 24642 43052 24676 43068
rect 23618 42964 23632 43016
rect 23618 42760 23620 42964
rect 23574 41958 23620 42760
rect 23574 41666 23584 41958
rect 23618 41666 23620 41958
rect 23574 40864 23620 41666
rect 23574 40572 23584 40864
rect 23618 40572 23620 40864
rect 23574 39770 23620 40572
rect 23574 39478 23584 39770
rect 23618 39478 23620 39770
rect 23574 38676 23620 39478
rect 23574 38618 23584 38676
rect 22560 38384 22588 38484
rect 22506 38274 22588 38384
rect 23618 38618 23620 38676
rect 25674 43052 25758 43194
rect 27976 43068 28044 43194
rect 24676 42760 24688 42964
rect 25674 42960 25700 43052
rect 24642 41958 24688 42760
rect 24676 41666 24688 41958
rect 24642 40864 24688 41666
rect 24676 40572 24688 40864
rect 24642 39770 24688 40572
rect 24676 39478 24688 39770
rect 24642 38676 24688 39478
rect 23584 38368 23618 38384
rect 24632 38384 24642 38456
rect 24676 38602 24688 38676
rect 25694 42760 25700 42960
rect 25734 42960 25758 43052
rect 26758 43052 26792 43068
rect 25734 42760 25740 42960
rect 25694 41958 25740 42760
rect 25694 41666 25700 41958
rect 25734 41666 25740 41958
rect 25694 40864 25740 41666
rect 25694 40572 25700 40864
rect 25734 40572 25740 40864
rect 25694 39770 25740 40572
rect 25694 39478 25700 39770
rect 25734 39478 25740 39770
rect 25694 38676 25740 39478
rect 25694 38646 25700 38676
rect 24676 38384 24714 38456
rect 24632 38274 24714 38384
rect 25734 38646 25740 38676
rect 26750 42760 26758 42980
rect 26792 42760 26796 42980
rect 26750 41958 26796 42760
rect 26750 41666 26758 41958
rect 26792 41666 26796 41958
rect 26750 40864 26796 41666
rect 27976 42776 27990 43068
rect 28024 42966 28044 43068
rect 29048 43068 29082 43084
rect 27976 42760 28024 42776
rect 29044 42776 29048 42974
rect 30080 43068 30148 43246
rect 32170 43162 35080 43252
rect 30080 42980 30106 43068
rect 29082 42776 29090 42974
rect 27976 41990 28022 42760
rect 27976 41974 28024 41990
rect 27976 41682 27990 41974
rect 27976 41666 28024 41682
rect 29044 41974 29090 42776
rect 29044 41682 29048 41974
rect 29082 41682 29090 41974
rect 26750 40572 26758 40864
rect 26792 40572 26796 40864
rect 26750 39770 26796 40572
rect 27336 41534 27486 41660
rect 27336 40338 27358 41534
rect 27452 40338 27486 41534
rect 27336 40014 27486 40338
rect 27976 40896 28022 41666
rect 27976 40880 28024 40896
rect 27976 40588 27990 40880
rect 27976 40572 28024 40588
rect 29044 40880 29090 41682
rect 29044 40588 29048 40880
rect 29082 40588 29090 40880
rect 26750 39478 26758 39770
rect 26792 39478 26796 39770
rect 26750 38676 26796 39478
rect 27976 39802 28022 40572
rect 27976 39786 28024 39802
rect 27976 39494 27990 39786
rect 27976 39478 28024 39494
rect 29044 39786 29090 40588
rect 29044 39494 29048 39786
rect 29082 39494 29090 39786
rect 27976 38798 28022 39478
rect 26750 38618 26758 38676
rect 25700 38368 25734 38384
rect 26704 38384 26758 38530
rect 26792 38618 26796 38676
rect 27970 38692 28102 38798
rect 26792 38384 26836 38530
rect 26704 38274 26836 38384
rect 27970 38400 27990 38692
rect 28024 38400 28102 38692
rect 29044 38692 29090 39494
rect 29044 38612 29048 38692
rect 22506 38184 26956 38274
rect 22518 38178 26956 38184
rect 24632 38156 24714 38178
rect 23558 37514 23626 37530
rect 25682 37514 25750 37546
rect 21426 37504 25750 37514
rect 21316 37460 25750 37504
rect 21316 37424 25758 37460
rect 21316 37414 25606 37424
rect 21426 37308 21558 37414
rect 19244 36960 19250 37160
rect 19204 36158 19250 36960
rect 19204 35866 19210 36158
rect 19244 35866 19250 36158
rect 19204 35064 19250 35866
rect 19204 34772 19210 35064
rect 19244 34772 19250 35064
rect 19204 33970 19250 34772
rect 19204 33678 19210 33970
rect 19244 33678 19250 33970
rect 19204 32876 19250 33678
rect 19204 32846 19210 32876
rect 18186 32584 18224 32656
rect 18142 32474 18224 32584
rect 19244 32846 19250 32876
rect 20242 36960 20268 37252
rect 20302 36960 20336 37252
rect 20242 36158 20336 36960
rect 20242 35866 20268 36158
rect 20302 35866 20336 36158
rect 20242 35064 20336 35866
rect 21454 37236 21522 37308
rect 21454 36944 21468 37236
rect 21502 37134 21522 37236
rect 22526 37236 22560 37252
rect 21454 36928 21502 36944
rect 22522 36944 22526 37142
rect 23558 37236 23626 37414
rect 23558 37148 23584 37236
rect 22560 36944 22568 37142
rect 21454 36158 21500 36928
rect 21454 36142 21502 36158
rect 21454 35850 21468 36142
rect 21454 35834 21502 35850
rect 22522 36142 22568 36944
rect 22522 35850 22526 36142
rect 22560 35850 22568 36142
rect 20242 34772 20268 35064
rect 20302 34772 20336 35064
rect 20242 33970 20336 34772
rect 20814 35702 20964 35828
rect 20814 34506 20836 35702
rect 20930 34506 20964 35702
rect 20814 34182 20964 34506
rect 21454 35064 21500 35834
rect 21454 35048 21502 35064
rect 21454 34756 21468 35048
rect 21454 34740 21502 34756
rect 22522 35048 22568 35850
rect 22522 34756 22526 35048
rect 22560 34756 22568 35048
rect 20242 33678 20268 33970
rect 20302 33678 20336 33970
rect 20242 32876 20336 33678
rect 21454 33970 21500 34740
rect 21454 33954 21502 33970
rect 21454 33662 21468 33954
rect 21454 33646 21502 33662
rect 22522 33954 22568 34756
rect 22522 33662 22526 33954
rect 22560 33662 22568 33954
rect 21454 32916 21500 33646
rect 19210 32568 19244 32584
rect 20242 32584 20268 32876
rect 20302 32730 20336 32876
rect 21440 32860 21572 32916
rect 20302 32584 20380 32730
rect 20242 32474 20380 32584
rect 21440 32568 21468 32860
rect 21502 32568 21572 32860
rect 22522 32860 22568 33662
rect 22522 32780 22526 32860
rect 16016 32384 20466 32474
rect 16028 32378 20466 32384
rect 18142 32356 18224 32378
rect 14940 31696 15032 31706
rect 17068 31696 17136 31712
rect 19192 31696 19260 31728
rect 14940 31686 19260 31696
rect 14826 31642 19260 31686
rect 14826 31606 19268 31642
rect 14826 31596 19116 31606
rect 11680 31118 11692 31322
rect 12678 31318 12704 31410
rect 11646 30316 11692 31118
rect 11680 30024 11692 30316
rect 11646 29222 11692 30024
rect 11680 28930 11692 29222
rect 11646 28128 11692 28930
rect 11680 27836 11692 28128
rect 11646 27034 11692 27836
rect 10588 26726 10622 26742
rect 11636 26742 11646 26814
rect 11680 26960 11692 27034
rect 12698 31118 12704 31318
rect 12738 31318 12762 31410
rect 13762 31410 13874 31426
rect 12738 31118 12744 31318
rect 12698 30316 12744 31118
rect 12698 30024 12704 30316
rect 12738 30024 12744 30316
rect 12698 29222 12744 30024
rect 12698 28930 12704 29222
rect 12738 28930 12744 29222
rect 12698 28128 12744 28930
rect 12698 27836 12704 28128
rect 12738 27836 12744 28128
rect 12698 27034 12744 27836
rect 12698 27004 12704 27034
rect 11680 26742 11718 26814
rect 11636 26632 11718 26742
rect 12738 27004 12744 27034
rect 13754 31118 13762 31338
rect 13796 31118 13874 31410
rect 13754 30316 13874 31118
rect 13754 30024 13762 30316
rect 13796 30024 13874 30316
rect 13754 29222 13874 30024
rect 14940 31418 15032 31596
rect 14940 31126 14978 31418
rect 15012 31316 15032 31418
rect 16036 31418 16070 31434
rect 15012 31126 15028 31316
rect 14940 30324 15028 31126
rect 14940 30032 14978 30324
rect 15012 30032 15028 30324
rect 13754 28930 13762 29222
rect 13796 28930 13874 29222
rect 13754 28128 13874 28930
rect 14324 29884 14474 30010
rect 14324 28688 14346 29884
rect 14440 28688 14474 29884
rect 14324 28364 14474 28688
rect 14940 29230 15028 30032
rect 14940 28938 14978 29230
rect 15012 28938 15028 29230
rect 13754 27836 13762 28128
rect 13796 27836 13874 28128
rect 13754 27034 13874 27836
rect 13754 26976 13762 27034
rect 12704 26726 12738 26742
rect 13738 26742 13762 26836
rect 13796 26742 13874 27034
rect 13738 26632 13874 26742
rect 14940 28136 15028 28938
rect 14940 27844 14978 28136
rect 15012 27844 15028 28136
rect 14940 27042 15028 27844
rect 14940 26750 14978 27042
rect 15012 26750 15028 27042
rect 16032 31126 16036 31324
rect 17068 31418 17136 31596
rect 17068 31330 17094 31418
rect 16070 31126 16078 31324
rect 16032 30324 16078 31126
rect 16032 30032 16036 30324
rect 16070 30032 16078 30324
rect 16032 29230 16078 30032
rect 16032 28938 16036 29230
rect 16070 28938 16078 29230
rect 16032 28136 16078 28938
rect 16032 27844 16036 28136
rect 16070 27844 16078 28136
rect 16032 27042 16078 27844
rect 16032 26962 16036 27042
rect 9510 26542 13960 26632
rect 9522 26536 13960 26542
rect 11636 26514 11718 26536
rect 10562 25852 10630 25868
rect 12686 25852 12754 25884
rect 8436 25842 12754 25852
rect 8320 25798 12754 25842
rect 8320 25762 12762 25798
rect 8320 25752 12610 25762
rect 6224 25274 6230 25474
rect 6184 24472 6230 25274
rect 6184 24180 6190 24472
rect 6224 24180 6230 24472
rect 6184 23378 6230 24180
rect 6184 23086 6190 23378
rect 6224 23086 6230 23378
rect 6184 22284 6230 23086
rect 6184 21992 6190 22284
rect 6224 21992 6230 22284
rect 6184 21190 6230 21992
rect 6184 21160 6190 21190
rect 5166 20898 5204 20970
rect 5122 20788 5204 20898
rect 6224 21160 6230 21190
rect 7240 25274 7248 25566
rect 7282 25274 7376 25566
rect 7240 24472 7376 25274
rect 7240 24180 7248 24472
rect 7282 24180 7376 24472
rect 7240 23378 7376 24180
rect 8436 25574 8572 25752
rect 8436 25282 8472 25574
rect 8506 25282 8572 25574
rect 9530 25574 9564 25590
rect 8436 24480 8572 25282
rect 8436 24188 8472 24480
rect 8506 24188 8572 24480
rect 7240 23086 7248 23378
rect 7282 23086 7376 23378
rect 7240 22284 7376 23086
rect 7818 24040 7968 24166
rect 7818 22844 7840 24040
rect 7934 22844 7968 24040
rect 7818 22520 7968 22844
rect 8436 23386 8572 24188
rect 8436 23094 8472 23386
rect 8506 23094 8572 23386
rect 7240 21992 7248 22284
rect 7282 21992 7376 22284
rect 7240 21190 7376 21992
rect 7240 20992 7248 21190
rect 6190 20882 6224 20898
rect 7224 20898 7248 20992
rect 7282 20898 7376 21190
rect 7224 20788 7376 20898
rect 8436 22292 8572 23094
rect 8436 22000 8472 22292
rect 8506 22000 8572 22292
rect 8436 21198 8572 22000
rect 8436 20906 8472 21198
rect 8506 20906 8572 21198
rect 9526 25282 9530 25480
rect 10562 25574 10630 25752
rect 10562 25486 10588 25574
rect 9564 25282 9572 25480
rect 9526 24480 9572 25282
rect 9526 24188 9530 24480
rect 9564 24188 9572 24480
rect 9526 23386 9572 24188
rect 9526 23094 9530 23386
rect 9564 23094 9572 23386
rect 9526 22292 9572 23094
rect 9526 22000 9530 22292
rect 9564 22000 9572 22292
rect 9526 21198 9572 22000
rect 9526 21118 9530 21198
rect 2996 20698 7446 20788
rect 3008 20692 7446 20698
rect 5122 20670 5204 20692
rect 4048 19980 4116 19996
rect 6172 19980 6240 20012
rect 1910 19970 6240 19980
rect 1806 19926 6240 19970
rect 1806 19890 6248 19926
rect 1806 19880 6096 19890
rect 1910 19702 2046 19880
rect 1910 19410 1958 19702
rect 1992 19410 2046 19702
rect 3016 19702 3050 19718
rect 1910 18608 2046 19410
rect 1910 18316 1958 18608
rect 1992 18316 2046 18608
rect 1304 18168 1454 18294
rect 1304 16972 1326 18168
rect 1420 16972 1454 18168
rect 1304 16648 1454 16972
rect 1910 17514 2046 18316
rect 1910 17222 1958 17514
rect 1992 17222 2046 17514
rect 1910 16420 2046 17222
rect 1910 16128 1958 16420
rect 1992 16128 2046 16420
rect 1910 15326 2046 16128
rect 1910 15034 1958 15326
rect 1992 15034 2046 15326
rect 3012 19410 3016 19608
rect 4048 19702 4116 19880
rect 4048 19614 4074 19702
rect 3050 19410 3058 19608
rect 3012 18608 3058 19410
rect 3012 18316 3016 18608
rect 3050 18316 3058 18608
rect 3012 17514 3058 18316
rect 3012 17222 3016 17514
rect 3050 17222 3058 17514
rect 3012 16420 3058 17222
rect 3012 16128 3016 16420
rect 3050 16128 3058 16420
rect 3012 15326 3058 16128
rect 3012 15246 3016 15326
rect 1910 14124 2046 15034
rect 2996 15034 3016 15134
rect 3050 15246 3058 15326
rect 4064 19410 4074 19614
rect 4108 19666 4116 19702
rect 5132 19702 5166 19718
rect 4108 19614 4122 19666
rect 4108 19410 4110 19614
rect 4064 18608 4110 19410
rect 4064 18316 4074 18608
rect 4108 18316 4110 18608
rect 4064 17514 4110 18316
rect 4064 17222 4074 17514
rect 4108 17222 4110 17514
rect 4064 16420 4110 17222
rect 4064 16128 4074 16420
rect 4108 16128 4110 16420
rect 4064 15326 4110 16128
rect 4064 15268 4074 15326
rect 3050 15034 3078 15134
rect 2996 14924 3078 15034
rect 4108 15268 4110 15326
rect 6164 19702 6248 19890
rect 5166 19410 5178 19614
rect 6164 19610 6190 19702
rect 5132 18608 5178 19410
rect 5166 18316 5178 18608
rect 5132 17514 5178 18316
rect 5166 17222 5178 17514
rect 5132 16420 5178 17222
rect 5166 16128 5178 16420
rect 5132 15326 5178 16128
rect 4074 15018 4108 15034
rect 5122 15034 5132 15106
rect 5166 15252 5178 15326
rect 6184 19410 6190 19610
rect 6224 19610 6248 19702
rect 7240 19702 7376 20692
rect 8436 19988 8572 20906
rect 9510 20906 9530 21006
rect 9564 21118 9572 21198
rect 10578 25282 10588 25486
rect 10622 25538 10630 25574
rect 11646 25574 11680 25590
rect 10622 25486 10636 25538
rect 10622 25282 10624 25486
rect 10578 24480 10624 25282
rect 10578 24188 10588 24480
rect 10622 24188 10624 24480
rect 10578 23386 10624 24188
rect 10578 23094 10588 23386
rect 10622 23094 10624 23386
rect 10578 22292 10624 23094
rect 10578 22000 10588 22292
rect 10622 22000 10624 22292
rect 10578 21198 10624 22000
rect 10578 21140 10588 21198
rect 9564 20906 9592 21006
rect 9510 20796 9592 20906
rect 10622 21140 10624 21198
rect 12678 25574 12762 25762
rect 13768 25590 13874 26536
rect 14940 25870 15028 26750
rect 16016 26750 16036 26850
rect 16070 26962 16078 27042
rect 17084 31126 17094 31330
rect 17128 31382 17136 31418
rect 18152 31418 18186 31434
rect 17128 31330 17142 31382
rect 17128 31126 17130 31330
rect 17084 30324 17130 31126
rect 17084 30032 17094 30324
rect 17128 30032 17130 30324
rect 17084 29230 17130 30032
rect 17084 28938 17094 29230
rect 17128 28938 17130 29230
rect 17084 28136 17130 28938
rect 17084 27844 17094 28136
rect 17128 27844 17130 28136
rect 17084 27042 17130 27844
rect 17084 26984 17094 27042
rect 16070 26750 16098 26850
rect 16016 26640 16098 26750
rect 17128 26984 17130 27042
rect 19184 31418 19268 31606
rect 18186 31126 18198 31330
rect 19184 31326 19210 31418
rect 18152 30324 18198 31126
rect 18186 30032 18198 30324
rect 18152 29230 18198 30032
rect 18186 28938 18198 29230
rect 18152 28136 18198 28938
rect 18186 27844 18198 28136
rect 18152 27042 18198 27844
rect 17094 26734 17128 26750
rect 18142 26750 18152 26822
rect 18186 26968 18198 27042
rect 19204 31126 19210 31326
rect 19244 31326 19268 31418
rect 20242 31418 20380 32378
rect 21440 31680 21572 32568
rect 22506 32568 22526 32668
rect 22560 32780 22568 32860
rect 23574 36944 23584 37148
rect 23618 37200 23626 37236
rect 24642 37236 24676 37252
rect 23618 37148 23632 37200
rect 23618 36944 23620 37148
rect 23574 36142 23620 36944
rect 23574 35850 23584 36142
rect 23618 35850 23620 36142
rect 23574 35048 23620 35850
rect 23574 34756 23584 35048
rect 23618 34756 23620 35048
rect 23574 33954 23620 34756
rect 23574 33662 23584 33954
rect 23618 33662 23620 33954
rect 23574 32860 23620 33662
rect 23574 32802 23584 32860
rect 22560 32568 22588 32668
rect 22506 32458 22588 32568
rect 23618 32802 23620 32860
rect 25674 37236 25758 37424
rect 24676 36944 24688 37148
rect 25674 37144 25700 37236
rect 24642 36142 24688 36944
rect 24676 35850 24688 36142
rect 24642 35048 24688 35850
rect 24676 34756 24688 35048
rect 24642 33954 24688 34756
rect 24676 33662 24688 33954
rect 24642 32860 24688 33662
rect 23584 32552 23618 32568
rect 24632 32568 24642 32640
rect 24676 32786 24688 32860
rect 25694 36944 25700 37144
rect 25734 37144 25758 37236
rect 26704 37236 26836 38178
rect 27970 37530 28102 38400
rect 29028 38400 29048 38500
rect 29082 38612 29090 38692
rect 30096 42776 30106 42980
rect 30140 43032 30148 43068
rect 31164 43068 31198 43084
rect 30140 42980 30154 43032
rect 30140 42776 30142 42980
rect 30096 41974 30142 42776
rect 30096 41682 30106 41974
rect 30140 41682 30142 41974
rect 30096 40880 30142 41682
rect 30096 40588 30106 40880
rect 30140 40588 30142 40880
rect 30096 39786 30142 40588
rect 30096 39494 30106 39786
rect 30140 39494 30142 39786
rect 30096 38692 30142 39494
rect 30096 38634 30106 38692
rect 29082 38400 29110 38500
rect 29028 38290 29110 38400
rect 30140 38634 30142 38692
rect 32196 43068 32280 43162
rect 31198 42776 31210 42980
rect 32196 42976 32222 43068
rect 31164 41974 31210 42776
rect 31198 41682 31210 41974
rect 31164 40880 31210 41682
rect 31198 40588 31210 40880
rect 31164 39786 31210 40588
rect 31198 39494 31210 39786
rect 31164 38692 31210 39494
rect 30106 38384 30140 38400
rect 31154 38400 31164 38472
rect 31198 38618 31210 38692
rect 32216 42776 32222 42976
rect 32256 42976 32280 43068
rect 33280 43068 33314 43084
rect 32256 42776 32262 42976
rect 32216 41974 32262 42776
rect 32216 41682 32222 41974
rect 32256 41682 32262 41974
rect 32216 40880 32262 41682
rect 32216 40588 32222 40880
rect 32256 40588 32262 40880
rect 32216 39786 32262 40588
rect 32216 39494 32222 39786
rect 32256 39494 32262 39786
rect 32216 38692 32262 39494
rect 32216 38662 32222 38692
rect 31198 38400 31236 38472
rect 31154 38290 31236 38400
rect 32256 38662 32262 38692
rect 33272 42776 33280 42996
rect 34486 43074 34554 43162
rect 33314 42776 33318 42996
rect 33272 41974 33318 42776
rect 33272 41682 33280 41974
rect 33314 41682 33318 41974
rect 33272 40880 33318 41682
rect 34486 42782 34500 43074
rect 34534 42972 34554 43074
rect 35558 43074 35592 43090
rect 34486 42766 34534 42782
rect 35554 42782 35558 42980
rect 36590 43074 36658 43252
rect 38462 43162 38792 43252
rect 36590 42986 36616 43074
rect 35592 42782 35600 42980
rect 34486 41996 34532 42766
rect 34486 41980 34534 41996
rect 34486 41688 34500 41980
rect 34486 41672 34534 41688
rect 35554 41980 35600 42782
rect 35554 41688 35558 41980
rect 35592 41688 35600 41980
rect 33272 40588 33280 40880
rect 33314 40588 33318 40880
rect 33272 39786 33318 40588
rect 33846 41540 33996 41666
rect 33846 40344 33868 41540
rect 33962 40344 33996 41540
rect 33846 40020 33996 40344
rect 34486 40902 34532 41672
rect 34486 40886 34534 40902
rect 34486 40594 34500 40886
rect 34486 40578 34534 40594
rect 35554 40886 35600 41688
rect 35554 40594 35558 40886
rect 35592 40594 35600 40886
rect 33272 39494 33280 39786
rect 33314 39494 33318 39786
rect 33272 38692 33318 39494
rect 34486 39808 34532 40578
rect 34486 39792 34534 39808
rect 34486 39500 34500 39792
rect 34486 39484 34534 39500
rect 35554 39792 35600 40594
rect 35554 39500 35558 39792
rect 35592 39500 35600 39792
rect 34486 38718 34532 39484
rect 33272 38634 33280 38692
rect 32222 38384 32256 38400
rect 33250 38400 33280 38494
rect 33314 38634 33318 38692
rect 34444 38698 34566 38718
rect 33314 38400 33382 38494
rect 34444 38462 34500 38698
rect 33250 38290 33382 38400
rect 34450 38406 34500 38462
rect 34534 38510 34566 38698
rect 35554 38698 35600 39500
rect 35554 38618 35558 38698
rect 34534 38406 34576 38510
rect 29028 38200 33478 38290
rect 29040 38194 33478 38200
rect 31154 38172 31236 38194
rect 30080 37530 30148 37546
rect 32204 37530 32272 37562
rect 27970 37520 32272 37530
rect 27838 37476 32272 37520
rect 27838 37440 32280 37476
rect 27838 37430 32128 37440
rect 27970 37390 28102 37430
rect 25734 36944 25740 37144
rect 26704 37122 26758 37236
rect 25694 36142 25740 36944
rect 25694 35850 25700 36142
rect 25734 35850 25740 36142
rect 25694 35048 25740 35850
rect 25694 34756 25700 35048
rect 25734 34756 25740 35048
rect 25694 33954 25740 34756
rect 25694 33662 25700 33954
rect 25734 33662 25740 33954
rect 25694 32860 25740 33662
rect 25694 32830 25700 32860
rect 24676 32568 24714 32640
rect 24632 32458 24714 32568
rect 25734 32830 25740 32860
rect 26750 36944 26758 37122
rect 26792 37122 26836 37236
rect 27976 37252 28044 37390
rect 26792 36944 26796 37122
rect 26750 36142 26796 36944
rect 26750 35850 26758 36142
rect 26792 35850 26796 36142
rect 26750 35048 26796 35850
rect 27976 36960 27990 37252
rect 28024 37150 28044 37252
rect 29048 37252 29082 37268
rect 27976 36944 28024 36960
rect 29044 36960 29048 37158
rect 30080 37252 30148 37430
rect 30080 37164 30106 37252
rect 29082 36960 29090 37158
rect 27976 36174 28022 36944
rect 27976 36158 28024 36174
rect 27976 35866 27990 36158
rect 27976 35850 28024 35866
rect 29044 36158 29090 36960
rect 29044 35866 29048 36158
rect 29082 35866 29090 36158
rect 26750 34756 26758 35048
rect 26792 34756 26796 35048
rect 26750 33954 26796 34756
rect 27336 35718 27486 35844
rect 27336 34522 27358 35718
rect 27452 34522 27486 35718
rect 27336 34198 27486 34522
rect 27976 35080 28022 35850
rect 27976 35064 28024 35080
rect 27976 34772 27990 35064
rect 27976 34756 28024 34772
rect 29044 35064 29090 35866
rect 29044 34772 29048 35064
rect 29082 34772 29090 35064
rect 26750 33662 26758 33954
rect 26792 33662 26796 33954
rect 26750 32860 26796 33662
rect 27976 33986 28022 34756
rect 27976 33970 28024 33986
rect 27976 33678 27990 33970
rect 27976 33662 28024 33678
rect 29044 33970 29090 34772
rect 29044 33678 29048 33970
rect 29082 33678 29090 33970
rect 27976 32954 28022 33662
rect 26750 32802 26758 32860
rect 25700 32552 25734 32568
rect 26734 32568 26758 32662
rect 26792 32802 26796 32860
rect 27948 32876 28080 32954
rect 26792 32648 26816 32662
rect 26792 32568 26880 32648
rect 26734 32458 26880 32568
rect 27948 32584 27990 32876
rect 28024 32584 28080 32876
rect 29044 32876 29090 33678
rect 29044 32796 29048 32876
rect 22506 32368 26956 32458
rect 22518 32362 26956 32368
rect 24632 32340 24714 32362
rect 23558 31680 23626 31696
rect 25682 31680 25750 31712
rect 21440 31670 25750 31680
rect 21316 31626 25750 31670
rect 21316 31590 25758 31626
rect 21316 31580 25606 31590
rect 21440 31508 21572 31580
rect 19244 31126 19250 31326
rect 19204 30324 19250 31126
rect 19204 30032 19210 30324
rect 19244 30032 19250 30324
rect 19204 29230 19250 30032
rect 19204 28938 19210 29230
rect 19244 28938 19250 29230
rect 19204 28136 19250 28938
rect 19204 27844 19210 28136
rect 19244 27844 19250 28136
rect 19204 27042 19250 27844
rect 19204 27012 19210 27042
rect 18186 26750 18224 26822
rect 18142 26640 18224 26750
rect 19244 27012 19250 27042
rect 20242 31126 20268 31418
rect 20302 31322 20380 31418
rect 21454 31402 21522 31508
rect 20302 31126 20336 31322
rect 20242 30324 20336 31126
rect 20242 30032 20268 30324
rect 20302 30032 20336 30324
rect 20242 29230 20336 30032
rect 21454 31110 21468 31402
rect 21502 31300 21522 31402
rect 22526 31402 22560 31418
rect 21454 31094 21502 31110
rect 22522 31110 22526 31308
rect 23558 31402 23626 31580
rect 23558 31314 23584 31402
rect 22560 31110 22568 31308
rect 21454 30324 21500 31094
rect 21454 30308 21502 30324
rect 21454 30016 21468 30308
rect 21454 30000 21502 30016
rect 22522 30308 22568 31110
rect 22522 30016 22526 30308
rect 22560 30016 22568 30308
rect 20242 28938 20268 29230
rect 20302 28938 20336 29230
rect 20242 28136 20336 28938
rect 20814 29868 20964 29994
rect 20814 28672 20836 29868
rect 20930 28672 20964 29868
rect 20814 28348 20964 28672
rect 21454 29230 21500 30000
rect 21454 29214 21502 29230
rect 21454 28922 21468 29214
rect 21454 28906 21502 28922
rect 22522 29214 22568 30016
rect 22522 28922 22526 29214
rect 22560 28922 22568 29214
rect 20242 27844 20268 28136
rect 20302 27844 20336 28136
rect 20242 27042 20336 27844
rect 21454 28136 21500 28906
rect 21454 28120 21502 28136
rect 21454 27828 21468 28120
rect 21454 27812 21502 27828
rect 22522 28120 22568 28922
rect 22522 27828 22526 28120
rect 22560 27828 22568 28120
rect 21454 27072 21500 27812
rect 20242 26864 20268 27042
rect 19210 26734 19244 26750
rect 20240 26750 20268 26864
rect 20302 26864 20336 27042
rect 21410 27026 21542 27072
rect 20302 26750 20372 26864
rect 20240 26640 20372 26750
rect 21410 26734 21468 27026
rect 21502 26734 21542 27026
rect 22522 27026 22568 27828
rect 22522 26946 22526 27026
rect 16016 26550 20466 26640
rect 16028 26544 20466 26550
rect 18142 26522 18224 26544
rect 14940 25860 15032 25870
rect 17068 25860 17136 25876
rect 19192 25860 19260 25892
rect 14940 25850 19260 25860
rect 14826 25806 19260 25850
rect 14826 25770 19268 25806
rect 14826 25760 19116 25770
rect 11680 25282 11692 25486
rect 12678 25482 12704 25574
rect 11646 24480 11692 25282
rect 11680 24188 11692 24480
rect 11646 23386 11692 24188
rect 11680 23094 11692 23386
rect 11646 22292 11692 23094
rect 11680 22000 11692 22292
rect 11646 21198 11692 22000
rect 10588 20890 10622 20906
rect 11636 20906 11646 20978
rect 11680 21124 11692 21198
rect 12698 25282 12704 25482
rect 12738 25482 12762 25574
rect 13762 25574 13874 25590
rect 12738 25282 12744 25482
rect 12698 24480 12744 25282
rect 12698 24188 12704 24480
rect 12738 24188 12744 24480
rect 12698 23386 12744 24188
rect 12698 23094 12704 23386
rect 12738 23094 12744 23386
rect 12698 22292 12744 23094
rect 12698 22000 12704 22292
rect 12738 22000 12744 22292
rect 12698 21198 12744 22000
rect 12698 21168 12704 21198
rect 11680 20906 11718 20978
rect 11636 20796 11718 20906
rect 12738 21168 12744 21198
rect 13754 25282 13762 25502
rect 13796 25282 13874 25574
rect 13754 24480 13874 25282
rect 13754 24188 13762 24480
rect 13796 24188 13874 24480
rect 13754 23386 13874 24188
rect 14940 25582 15032 25760
rect 14940 25290 14978 25582
rect 15012 25480 15032 25582
rect 16036 25582 16070 25598
rect 15012 25290 15028 25480
rect 14940 24488 15028 25290
rect 14940 24196 14978 24488
rect 15012 24196 15028 24488
rect 13754 23094 13762 23386
rect 13796 23094 13874 23386
rect 13754 22292 13874 23094
rect 14324 24048 14474 24174
rect 14324 22852 14346 24048
rect 14440 22852 14474 24048
rect 14324 22528 14474 22852
rect 14940 23394 15028 24196
rect 14940 23102 14978 23394
rect 15012 23102 15028 23394
rect 13754 22000 13762 22292
rect 13796 22000 13874 22292
rect 13754 21198 13874 22000
rect 13754 21140 13762 21198
rect 12704 20890 12738 20906
rect 13738 20906 13762 21000
rect 13796 20906 13874 21198
rect 13738 20796 13874 20906
rect 14940 22300 15028 23102
rect 14940 22008 14978 22300
rect 15012 22008 15028 22300
rect 14940 21206 15028 22008
rect 14940 20914 14978 21206
rect 15012 20914 15028 21206
rect 16032 25290 16036 25488
rect 17068 25582 17136 25760
rect 17068 25494 17094 25582
rect 16070 25290 16078 25488
rect 16032 24488 16078 25290
rect 16032 24196 16036 24488
rect 16070 24196 16078 24488
rect 16032 23394 16078 24196
rect 16032 23102 16036 23394
rect 16070 23102 16078 23394
rect 16032 22300 16078 23102
rect 16032 22008 16036 22300
rect 16070 22008 16078 22300
rect 16032 21206 16078 22008
rect 16032 21126 16036 21206
rect 9510 20706 13960 20796
rect 9522 20700 13960 20706
rect 11636 20678 11718 20700
rect 10562 19988 10630 20004
rect 12686 19988 12754 20020
rect 8436 19978 12754 19988
rect 8320 19934 12754 19978
rect 8320 19898 12762 19934
rect 8320 19888 12610 19898
rect 6224 19410 6230 19610
rect 6184 18608 6230 19410
rect 6184 18316 6190 18608
rect 6224 18316 6230 18608
rect 6184 17514 6230 18316
rect 6184 17222 6190 17514
rect 6224 17222 6230 17514
rect 6184 16420 6230 17222
rect 6184 16128 6190 16420
rect 6224 16128 6230 16420
rect 6184 15326 6230 16128
rect 6184 15296 6190 15326
rect 5166 15034 5204 15106
rect 5122 14924 5204 15034
rect 6224 15296 6230 15326
rect 7240 19410 7248 19702
rect 7282 19410 7376 19702
rect 7240 18608 7376 19410
rect 7240 18316 7248 18608
rect 7282 18316 7376 18608
rect 7240 17514 7376 18316
rect 8436 19710 8572 19888
rect 8436 19418 8472 19710
rect 8506 19418 8572 19710
rect 9530 19710 9564 19726
rect 8436 18616 8572 19418
rect 8436 18324 8472 18616
rect 8506 18324 8572 18616
rect 7240 17222 7248 17514
rect 7282 17222 7376 17514
rect 7240 16420 7376 17222
rect 7818 18176 7968 18302
rect 7818 16980 7840 18176
rect 7934 16980 7968 18176
rect 7818 16656 7968 16980
rect 8436 17522 8572 18324
rect 8436 17230 8472 17522
rect 8506 17230 8572 17522
rect 7240 16128 7248 16420
rect 7282 16128 7376 16420
rect 7240 15326 7376 16128
rect 7240 15128 7248 15326
rect 6190 15018 6224 15034
rect 7224 15034 7248 15128
rect 7282 15034 7376 15326
rect 7224 14924 7376 15034
rect 8436 16428 8572 17230
rect 8436 16136 8472 16428
rect 8506 16136 8572 16428
rect 8436 15334 8572 16136
rect 8436 15042 8472 15334
rect 8506 15042 8572 15334
rect 9526 19418 9530 19616
rect 10562 19710 10630 19888
rect 10562 19622 10588 19710
rect 9564 19418 9572 19616
rect 9526 18616 9572 19418
rect 9526 18324 9530 18616
rect 9564 18324 9572 18616
rect 9526 17522 9572 18324
rect 9526 17230 9530 17522
rect 9564 17230 9572 17522
rect 9526 16428 9572 17230
rect 9526 16136 9530 16428
rect 9564 16136 9572 16428
rect 9526 15334 9572 16136
rect 9526 15254 9530 15334
rect 2996 14834 7446 14924
rect 3008 14828 7446 14834
rect 5122 14806 5204 14828
rect 4058 14124 4126 14140
rect 6182 14124 6250 14156
rect 1910 14114 6250 14124
rect 1816 14070 6250 14114
rect 1816 14034 6258 14070
rect 1816 14024 6106 14034
rect 1910 13846 2046 14024
rect 1910 13554 1968 13846
rect 2002 13554 2046 13846
rect 3026 13846 3060 13862
rect 1910 12752 2046 13554
rect 1910 12460 1968 12752
rect 2002 12460 2046 12752
rect 1314 12312 1464 12438
rect 1314 11116 1336 12312
rect 1430 11116 1464 12312
rect 1314 10792 1464 11116
rect 1910 11658 2046 12460
rect 1910 11366 1968 11658
rect 2002 11366 2046 11658
rect 1910 10564 2046 11366
rect 1910 10272 1968 10564
rect 2002 10272 2046 10564
rect 1910 9470 2046 10272
rect 1910 9178 1968 9470
rect 2002 9178 2046 9470
rect 3022 13554 3026 13752
rect 4058 13846 4126 14024
rect 4058 13758 4084 13846
rect 3060 13554 3068 13752
rect 3022 12752 3068 13554
rect 3022 12460 3026 12752
rect 3060 12460 3068 12752
rect 3022 11658 3068 12460
rect 3022 11366 3026 11658
rect 3060 11366 3068 11658
rect 3022 10564 3068 11366
rect 3022 10272 3026 10564
rect 3060 10272 3068 10564
rect 3022 9470 3068 10272
rect 3022 9390 3026 9470
rect 1910 8216 2046 9178
rect 3006 9178 3026 9278
rect 3060 9390 3068 9470
rect 4074 13554 4084 13758
rect 4118 13810 4126 13846
rect 5142 13846 5176 13862
rect 4118 13758 4132 13810
rect 4118 13554 4120 13758
rect 4074 12752 4120 13554
rect 4074 12460 4084 12752
rect 4118 12460 4120 12752
rect 4074 11658 4120 12460
rect 4074 11366 4084 11658
rect 4118 11366 4120 11658
rect 4074 10564 4120 11366
rect 4074 10272 4084 10564
rect 4118 10272 4120 10564
rect 4074 9470 4120 10272
rect 4074 9412 4084 9470
rect 3060 9178 3088 9278
rect 3006 9068 3088 9178
rect 4118 9412 4120 9470
rect 6174 13846 6258 14034
rect 5176 13554 5188 13758
rect 6174 13754 6200 13846
rect 5142 12752 5188 13554
rect 5176 12460 5188 12752
rect 5142 11658 5188 12460
rect 5176 11366 5188 11658
rect 5142 10564 5188 11366
rect 5176 10272 5188 10564
rect 5142 9470 5188 10272
rect 4084 9162 4118 9178
rect 5132 9178 5142 9250
rect 5176 9396 5188 9470
rect 6194 13554 6200 13754
rect 6234 13754 6258 13846
rect 7240 13846 7376 14828
rect 8436 14132 8572 15042
rect 9510 15042 9530 15142
rect 9564 15254 9572 15334
rect 10578 19418 10588 19622
rect 10622 19674 10630 19710
rect 11646 19710 11680 19726
rect 10622 19622 10636 19674
rect 10622 19418 10624 19622
rect 10578 18616 10624 19418
rect 10578 18324 10588 18616
rect 10622 18324 10624 18616
rect 10578 17522 10624 18324
rect 10578 17230 10588 17522
rect 10622 17230 10624 17522
rect 10578 16428 10624 17230
rect 10578 16136 10588 16428
rect 10622 16136 10624 16428
rect 10578 15334 10624 16136
rect 10578 15276 10588 15334
rect 9564 15042 9592 15142
rect 9510 14932 9592 15042
rect 10622 15276 10624 15334
rect 12678 19710 12762 19898
rect 13768 19726 13874 20700
rect 14940 20006 15028 20914
rect 16016 20914 16036 21014
rect 16070 21126 16078 21206
rect 17084 25290 17094 25494
rect 17128 25546 17136 25582
rect 18152 25582 18186 25598
rect 17128 25494 17142 25546
rect 17128 25290 17130 25494
rect 17084 24488 17130 25290
rect 17084 24196 17094 24488
rect 17128 24196 17130 24488
rect 17084 23394 17130 24196
rect 17084 23102 17094 23394
rect 17128 23102 17130 23394
rect 17084 22300 17130 23102
rect 17084 22008 17094 22300
rect 17128 22008 17130 22300
rect 17084 21206 17130 22008
rect 17084 21148 17094 21206
rect 16070 20914 16098 21014
rect 16016 20804 16098 20914
rect 17128 21148 17130 21206
rect 19184 25582 19268 25770
rect 18186 25290 18198 25494
rect 19184 25490 19210 25582
rect 18152 24488 18198 25290
rect 18186 24196 18198 24488
rect 18152 23394 18198 24196
rect 18186 23102 18198 23394
rect 18152 22300 18198 23102
rect 18186 22008 18198 22300
rect 18152 21206 18198 22008
rect 17094 20898 17128 20914
rect 18142 20914 18152 20986
rect 18186 21132 18198 21206
rect 19204 25290 19210 25490
rect 19244 25490 19268 25582
rect 20240 25582 20372 26544
rect 21410 25844 21542 26734
rect 22506 26734 22526 26834
rect 22560 26946 22568 27026
rect 23574 31110 23584 31314
rect 23618 31366 23626 31402
rect 24642 31402 24676 31418
rect 23618 31314 23632 31366
rect 23618 31110 23620 31314
rect 23574 30308 23620 31110
rect 23574 30016 23584 30308
rect 23618 30016 23620 30308
rect 23574 29214 23620 30016
rect 23574 28922 23584 29214
rect 23618 28922 23620 29214
rect 23574 28120 23620 28922
rect 23574 27828 23584 28120
rect 23618 27828 23620 28120
rect 23574 27026 23620 27828
rect 23574 26968 23584 27026
rect 22560 26734 22588 26834
rect 22506 26624 22588 26734
rect 23618 26968 23620 27026
rect 25674 31402 25758 31590
rect 24676 31110 24688 31314
rect 25674 31310 25700 31402
rect 24642 30308 24688 31110
rect 24676 30016 24688 30308
rect 24642 29214 24688 30016
rect 24676 28922 24688 29214
rect 24642 28120 24688 28922
rect 24676 27828 24688 28120
rect 24642 27026 24688 27828
rect 23584 26718 23618 26734
rect 24632 26734 24642 26806
rect 24676 26952 24688 27026
rect 25694 31110 25700 31310
rect 25734 31310 25758 31402
rect 26748 31402 26880 32362
rect 27948 31696 28080 32584
rect 29028 32584 29048 32684
rect 29082 32796 29090 32876
rect 30096 36960 30106 37164
rect 30140 37216 30148 37252
rect 31164 37252 31198 37268
rect 30140 37164 30154 37216
rect 30140 36960 30142 37164
rect 30096 36158 30142 36960
rect 30096 35866 30106 36158
rect 30140 35866 30142 36158
rect 30096 35064 30142 35866
rect 30096 34772 30106 35064
rect 30140 34772 30142 35064
rect 30096 33970 30142 34772
rect 30096 33678 30106 33970
rect 30140 33678 30142 33970
rect 30096 32876 30142 33678
rect 30096 32818 30106 32876
rect 29082 32584 29110 32684
rect 29028 32474 29110 32584
rect 30140 32818 30142 32876
rect 32196 37252 32280 37440
rect 31198 36960 31210 37164
rect 32196 37160 32222 37252
rect 31164 36158 31210 36960
rect 31198 35866 31210 36158
rect 31164 35064 31210 35866
rect 31198 34772 31210 35064
rect 31164 33970 31210 34772
rect 31198 33678 31210 33970
rect 31164 32876 31210 33678
rect 30106 32568 30140 32584
rect 31154 32584 31164 32656
rect 31198 32802 31210 32876
rect 32216 36960 32222 37160
rect 32256 37160 32280 37252
rect 33250 37252 33382 38194
rect 34450 37536 34576 38406
rect 35538 38406 35558 38506
rect 35592 38618 35600 38698
rect 36606 42782 36616 42986
rect 36650 43038 36658 43074
rect 37674 43074 37708 43090
rect 36650 42986 36664 43038
rect 36650 42782 36652 42986
rect 36606 41980 36652 42782
rect 36606 41688 36616 41980
rect 36650 41688 36652 41980
rect 36606 40886 36652 41688
rect 36606 40594 36616 40886
rect 36650 40594 36652 40886
rect 36606 39792 36652 40594
rect 36606 39500 36616 39792
rect 36650 39500 36652 39792
rect 36606 38698 36652 39500
rect 36606 38640 36616 38698
rect 35592 38406 35620 38506
rect 35538 38296 35620 38406
rect 36650 38640 36652 38698
rect 38706 43074 38790 43162
rect 39704 43110 40048 43878
rect 49454 43672 49550 43936
rect 49974 43672 50070 43936
rect 49454 43614 50070 43672
rect 63792 43632 64238 43652
rect 40976 43352 41044 43362
rect 43080 43352 43148 43368
rect 45204 43352 45272 43384
rect 47564 43374 47632 43384
rect 49642 43374 49838 43614
rect 63792 43466 63810 43632
rect 64200 43466 64238 43632
rect 51792 43374 51860 43406
rect 54078 43388 54146 43398
rect 56182 43388 56250 43404
rect 58306 43388 58374 43420
rect 54078 43380 58374 43388
rect 59348 43380 59446 43456
rect 63792 43444 64238 43466
rect 66242 43532 66422 46248
rect 68276 43950 69060 43984
rect 68276 43808 68330 43950
rect 68980 43808 69060 43950
rect 68276 43782 69060 43808
rect 67732 43614 68038 43628
rect 71570 43614 71878 43638
rect 67732 43584 68228 43614
rect 54078 43378 59446 43380
rect 47564 43364 51860 43374
rect 40976 43344 45272 43352
rect 40868 43342 45272 43344
rect 40838 43338 45272 43342
rect 47426 43360 51860 43364
rect 53940 43360 59446 43378
rect 47426 43338 59446 43360
rect 40838 43298 59446 43338
rect 40838 43288 58230 43298
rect 40838 43284 54496 43288
rect 40838 43274 51716 43284
rect 40838 43262 47900 43274
rect 40838 43252 45128 43262
rect 40868 43162 41130 43252
rect 37708 42782 37720 42986
rect 38706 42982 38732 43074
rect 37674 41980 37720 42782
rect 37708 41688 37720 41980
rect 37674 40886 37720 41688
rect 37708 40594 37720 40886
rect 37674 39792 37720 40594
rect 37708 39500 37720 39792
rect 37674 38698 37720 39500
rect 36616 38390 36650 38406
rect 37664 38406 37674 38478
rect 37708 38624 37720 38698
rect 38726 42782 38732 42982
rect 38766 42982 38790 43074
rect 39758 43074 39922 43110
rect 38766 42782 38772 42982
rect 38726 41980 38772 42782
rect 39758 42782 39790 43074
rect 39824 42782 39922 43074
rect 39758 42730 39922 42782
rect 40976 43074 41044 43162
rect 40976 42782 40990 43074
rect 41024 42972 41044 43074
rect 42048 43074 42082 43090
rect 40976 42766 41024 42782
rect 42044 42782 42048 42980
rect 43080 43074 43148 43252
rect 45182 43240 47900 43262
rect 43080 42986 43106 43074
rect 42082 42782 42090 42980
rect 38726 41688 38732 41980
rect 38766 41688 38772 41980
rect 38726 40886 38772 41688
rect 38726 40594 38732 40886
rect 38766 40594 38772 40886
rect 38726 39792 38772 40594
rect 38726 39500 38732 39792
rect 38766 39500 38772 39792
rect 38726 38698 38772 39500
rect 38726 38668 38732 38698
rect 37708 38406 37746 38478
rect 37664 38296 37746 38406
rect 38766 38668 38772 38698
rect 39782 41980 39828 42730
rect 39782 41688 39790 41980
rect 39824 41688 39828 41980
rect 39782 40886 39828 41688
rect 40976 41996 41022 42766
rect 40976 41980 41024 41996
rect 40976 41688 40990 41980
rect 40976 41672 41024 41688
rect 42044 41980 42090 42782
rect 42044 41688 42048 41980
rect 42082 41688 42090 41980
rect 39782 40594 39790 40886
rect 39824 40594 39828 40886
rect 39782 39792 39828 40594
rect 40336 41540 40486 41666
rect 40336 40344 40358 41540
rect 40452 40344 40486 41540
rect 40336 40020 40486 40344
rect 40976 40902 41022 41672
rect 40976 40886 41024 40902
rect 40976 40594 40990 40886
rect 40976 40578 41024 40594
rect 42044 40886 42090 41688
rect 42044 40594 42048 40886
rect 42082 40594 42090 40886
rect 39782 39500 39790 39792
rect 39824 39500 39828 39792
rect 39782 38698 39828 39500
rect 39782 38640 39790 38698
rect 38732 38390 38766 38406
rect 39766 38406 39790 38500
rect 39824 38640 39828 38698
rect 40976 39808 41022 40578
rect 40976 39792 41024 39808
rect 40976 39500 40990 39792
rect 40976 39484 41024 39500
rect 42044 39792 42090 40594
rect 42044 39500 42048 39792
rect 42082 39500 42090 39792
rect 40976 38714 41022 39484
rect 40976 38698 41024 38714
rect 40976 38640 40990 38698
rect 39824 38496 39848 38500
rect 39824 38406 39894 38496
rect 39766 38296 39894 38406
rect 40962 38406 40990 38596
rect 42044 38698 42090 39500
rect 42044 38618 42048 38698
rect 41024 38406 41088 38596
rect 35538 38206 39988 38296
rect 35550 38200 39988 38206
rect 37664 38178 37746 38200
rect 36590 37536 36658 37552
rect 38714 37536 38782 37568
rect 34450 37526 38782 37536
rect 34348 37482 38782 37526
rect 34348 37446 38790 37482
rect 34348 37436 38638 37446
rect 32256 36960 32262 37160
rect 33250 37086 33280 37252
rect 32216 36158 32262 36960
rect 32216 35866 32222 36158
rect 32256 35866 32262 36158
rect 32216 35064 32262 35866
rect 32216 34772 32222 35064
rect 32256 34772 32262 35064
rect 32216 33970 32262 34772
rect 32216 33678 32222 33970
rect 32256 33678 32262 33970
rect 32216 32876 32262 33678
rect 32216 32846 32222 32876
rect 31198 32584 31236 32656
rect 31154 32474 31236 32584
rect 32256 32846 32262 32876
rect 33272 36960 33280 37086
rect 33314 37086 33382 37252
rect 34450 37258 34576 37436
rect 34450 37126 34500 37258
rect 33314 36960 33318 37086
rect 33272 36158 33318 36960
rect 33272 35866 33280 36158
rect 33314 35866 33318 36158
rect 33272 35064 33318 35866
rect 34486 36966 34500 37126
rect 34534 37126 34576 37258
rect 35558 37258 35592 37274
rect 34486 36950 34534 36966
rect 35554 36966 35558 37164
rect 36590 37258 36658 37436
rect 36590 37170 36616 37258
rect 35592 36966 35600 37164
rect 34486 36180 34532 36950
rect 34486 36164 34534 36180
rect 34486 35872 34500 36164
rect 34486 35856 34534 35872
rect 35554 36164 35600 36966
rect 35554 35872 35558 36164
rect 35592 35872 35600 36164
rect 33272 34772 33280 35064
rect 33314 34772 33318 35064
rect 33272 33970 33318 34772
rect 33846 35724 33996 35850
rect 33846 34528 33868 35724
rect 33962 34528 33996 35724
rect 33846 34204 33996 34528
rect 34486 35086 34532 35856
rect 34486 35070 34534 35086
rect 34486 34778 34500 35070
rect 34486 34762 34534 34778
rect 35554 35070 35600 35872
rect 35554 34778 35558 35070
rect 35592 34778 35600 35070
rect 33272 33678 33280 33970
rect 33314 33678 33318 33970
rect 33272 32876 33318 33678
rect 33272 32818 33280 32876
rect 33256 32640 33280 32678
rect 32222 32568 32256 32584
rect 33228 32584 33280 32640
rect 33314 32818 33318 32876
rect 34486 33992 34532 34762
rect 34486 33976 34534 33992
rect 34486 33684 34500 33976
rect 34486 33668 34534 33684
rect 35554 33976 35600 34778
rect 35554 33684 35558 33976
rect 35592 33684 35600 33976
rect 34486 32898 34532 33668
rect 34486 32882 34534 32898
rect 34486 32824 34500 32882
rect 33314 32640 33338 32678
rect 33314 32584 33360 32640
rect 33228 32474 33360 32584
rect 34450 32590 34500 32772
rect 35554 32882 35600 33684
rect 35554 32802 35558 32882
rect 34534 32590 34576 32772
rect 29028 32384 33478 32474
rect 29040 32378 33478 32384
rect 31154 32356 31236 32378
rect 30080 31696 30148 31712
rect 32204 31696 32272 31728
rect 27948 31686 32272 31696
rect 27838 31642 32272 31686
rect 27838 31606 32280 31642
rect 27838 31596 32128 31606
rect 27948 31546 28080 31596
rect 25734 31110 25740 31310
rect 26748 31240 26758 31402
rect 25694 30308 25740 31110
rect 25694 30016 25700 30308
rect 25734 30016 25740 30308
rect 25694 29214 25740 30016
rect 25694 28922 25700 29214
rect 25734 28922 25740 29214
rect 25694 28120 25740 28922
rect 25694 27828 25700 28120
rect 25734 27828 25740 28120
rect 25694 27026 25740 27828
rect 25694 26996 25700 27026
rect 24676 26734 24714 26806
rect 24632 26624 24714 26734
rect 25734 26996 25740 27026
rect 26750 31110 26758 31240
rect 26792 31240 26880 31402
rect 27976 31418 28044 31546
rect 26792 31110 26796 31240
rect 26750 30308 26796 31110
rect 26750 30016 26758 30308
rect 26792 30016 26796 30308
rect 26750 29214 26796 30016
rect 27976 31126 27990 31418
rect 28024 31316 28044 31418
rect 29048 31418 29082 31434
rect 27976 31110 28024 31126
rect 29044 31126 29048 31324
rect 30080 31418 30148 31596
rect 30080 31330 30106 31418
rect 29082 31126 29090 31324
rect 27976 30340 28022 31110
rect 27976 30324 28024 30340
rect 27976 30032 27990 30324
rect 27976 30016 28024 30032
rect 29044 30324 29090 31126
rect 29044 30032 29048 30324
rect 29082 30032 29090 30324
rect 26750 28922 26758 29214
rect 26792 28922 26796 29214
rect 26750 28120 26796 28922
rect 27336 29884 27486 30010
rect 27336 28688 27358 29884
rect 27452 28688 27486 29884
rect 27336 28364 27486 28688
rect 27976 29246 28022 30016
rect 27976 29230 28024 29246
rect 27976 28938 27990 29230
rect 27976 28922 28024 28938
rect 29044 29230 29090 30032
rect 29044 28938 29048 29230
rect 29082 28938 29090 29230
rect 26750 27828 26758 28120
rect 26792 27828 26796 28120
rect 26750 27026 26796 27828
rect 27976 28152 28022 28922
rect 27976 28136 28024 28152
rect 27976 27844 27990 28136
rect 27976 27828 28024 27844
rect 29044 28136 29090 28938
rect 29044 27844 29048 28136
rect 29082 27844 29090 28136
rect 27976 27080 28022 27828
rect 26750 26968 26758 27026
rect 26740 26828 26758 26878
rect 25700 26718 25734 26734
rect 26734 26734 26758 26828
rect 26792 26968 26796 27026
rect 27964 27042 28096 27080
rect 26792 26734 26872 26878
rect 26734 26624 26872 26734
rect 27964 26750 27990 27042
rect 28024 26750 28096 27042
rect 29044 27042 29090 27844
rect 29044 26962 29048 27042
rect 22506 26534 26956 26624
rect 22518 26528 26956 26534
rect 24632 26506 24714 26528
rect 23558 25844 23626 25860
rect 25682 25844 25750 25876
rect 21410 25834 25750 25844
rect 21316 25790 25750 25834
rect 21316 25754 25758 25790
rect 21316 25744 25606 25754
rect 21410 25664 21542 25744
rect 19244 25290 19250 25490
rect 20240 25456 20268 25582
rect 19204 24488 19250 25290
rect 19204 24196 19210 24488
rect 19244 24196 19250 24488
rect 19204 23394 19250 24196
rect 19204 23102 19210 23394
rect 19244 23102 19250 23394
rect 19204 22300 19250 23102
rect 19204 22008 19210 22300
rect 19244 22008 19250 22300
rect 19204 21206 19250 22008
rect 19204 21176 19210 21206
rect 18186 20914 18224 20986
rect 18142 20804 18224 20914
rect 19244 21176 19250 21206
rect 20242 25290 20268 25456
rect 20302 25456 20372 25582
rect 21454 25566 21522 25664
rect 20302 25290 20336 25456
rect 20242 24488 20336 25290
rect 20242 24196 20268 24488
rect 20302 24196 20336 24488
rect 20242 23394 20336 24196
rect 21454 25274 21468 25566
rect 21502 25464 21522 25566
rect 22526 25566 22560 25582
rect 21454 25258 21502 25274
rect 22522 25274 22526 25472
rect 23558 25566 23626 25744
rect 23558 25478 23584 25566
rect 22560 25274 22568 25472
rect 21454 24488 21500 25258
rect 21454 24472 21502 24488
rect 21454 24180 21468 24472
rect 21454 24164 21502 24180
rect 22522 24472 22568 25274
rect 22522 24180 22526 24472
rect 22560 24180 22568 24472
rect 20242 23102 20268 23394
rect 20302 23102 20336 23394
rect 20242 22300 20336 23102
rect 20814 24032 20964 24158
rect 20814 22836 20836 24032
rect 20930 22836 20964 24032
rect 20814 22512 20964 22836
rect 21454 23394 21500 24164
rect 21454 23378 21502 23394
rect 21454 23086 21468 23378
rect 21454 23070 21502 23086
rect 22522 23378 22568 24180
rect 22522 23086 22526 23378
rect 22560 23086 22568 23378
rect 20242 22008 20268 22300
rect 20302 22008 20336 22300
rect 20242 21206 20336 22008
rect 19210 20898 19244 20914
rect 20242 20914 20268 21206
rect 20302 20914 20336 21206
rect 21454 22300 21500 23070
rect 21454 22284 21502 22300
rect 21454 21992 21468 22284
rect 21454 21976 21502 21992
rect 22522 22284 22568 23086
rect 22522 21992 22526 22284
rect 22560 21992 22568 22284
rect 21454 21206 21500 21976
rect 21454 21190 21502 21206
rect 21454 21134 21468 21190
rect 20242 20804 20336 20914
rect 21410 20898 21468 21134
rect 22522 21190 22568 21992
rect 21502 20898 21542 21134
rect 22522 21110 22526 21190
rect 16016 20714 20466 20804
rect 16028 20708 20466 20714
rect 18142 20686 18224 20708
rect 14940 19996 15032 20006
rect 17068 19996 17136 20012
rect 19192 19996 19260 20028
rect 14940 19986 19260 19996
rect 14826 19942 19260 19986
rect 14826 19906 19268 19942
rect 14826 19896 19116 19906
rect 11680 19418 11692 19622
rect 12678 19618 12704 19710
rect 11646 18616 11692 19418
rect 11680 18324 11692 18616
rect 11646 17522 11692 18324
rect 11680 17230 11692 17522
rect 11646 16428 11692 17230
rect 11680 16136 11692 16428
rect 11646 15334 11692 16136
rect 10588 15026 10622 15042
rect 11636 15042 11646 15114
rect 11680 15260 11692 15334
rect 12698 19418 12704 19618
rect 12738 19618 12762 19710
rect 13762 19710 13874 19726
rect 12738 19418 12744 19618
rect 12698 18616 12744 19418
rect 12698 18324 12704 18616
rect 12738 18324 12744 18616
rect 12698 17522 12744 18324
rect 12698 17230 12704 17522
rect 12738 17230 12744 17522
rect 12698 16428 12744 17230
rect 12698 16136 12704 16428
rect 12738 16136 12744 16428
rect 12698 15334 12744 16136
rect 12698 15304 12704 15334
rect 11680 15042 11718 15114
rect 11636 14932 11718 15042
rect 12738 15304 12744 15334
rect 13754 19418 13762 19638
rect 13796 19418 13874 19710
rect 13754 18616 13874 19418
rect 13754 18324 13762 18616
rect 13796 18324 13874 18616
rect 13754 17522 13874 18324
rect 14940 19718 15032 19896
rect 14940 19426 14978 19718
rect 15012 19616 15032 19718
rect 16036 19718 16070 19734
rect 15012 19426 15028 19616
rect 14940 18624 15028 19426
rect 14940 18332 14978 18624
rect 15012 18332 15028 18624
rect 13754 17230 13762 17522
rect 13796 17230 13874 17522
rect 13754 16428 13874 17230
rect 14324 18184 14474 18310
rect 14324 16988 14346 18184
rect 14440 16988 14474 18184
rect 14324 16664 14474 16988
rect 14940 17530 15028 18332
rect 14940 17238 14978 17530
rect 15012 17238 15028 17530
rect 13754 16136 13762 16428
rect 13796 16136 13874 16428
rect 13754 15334 13874 16136
rect 13754 15276 13762 15334
rect 12704 15026 12738 15042
rect 13738 15042 13762 15136
rect 13796 15042 13874 15334
rect 13738 14932 13874 15042
rect 14940 16436 15028 17238
rect 14940 16144 14978 16436
rect 15012 16144 15028 16436
rect 14940 15342 15028 16144
rect 14940 15050 14978 15342
rect 15012 15050 15028 15342
rect 16032 19426 16036 19624
rect 17068 19718 17136 19896
rect 17068 19630 17094 19718
rect 16070 19426 16078 19624
rect 16032 18624 16078 19426
rect 16032 18332 16036 18624
rect 16070 18332 16078 18624
rect 16032 17530 16078 18332
rect 16032 17238 16036 17530
rect 16070 17238 16078 17530
rect 16032 16436 16078 17238
rect 16032 16144 16036 16436
rect 16070 16144 16078 16436
rect 16032 15342 16078 16144
rect 16032 15262 16036 15342
rect 9510 14842 13960 14932
rect 9522 14836 13960 14842
rect 11636 14814 11718 14836
rect 10572 14132 10640 14148
rect 12696 14132 12764 14164
rect 8436 14122 12764 14132
rect 8330 14078 12764 14122
rect 8330 14042 12772 14078
rect 8330 14032 12620 14042
rect 6234 13554 6240 13754
rect 6194 12752 6240 13554
rect 6194 12460 6200 12752
rect 6234 12460 6240 12752
rect 6194 11658 6240 12460
rect 6194 11366 6200 11658
rect 6234 11366 6240 11658
rect 6194 10564 6240 11366
rect 6194 10272 6200 10564
rect 6234 10272 6240 10564
rect 6194 9470 6240 10272
rect 6194 9440 6200 9470
rect 5176 9178 5214 9250
rect 5132 9068 5214 9178
rect 6234 9440 6240 9470
rect 7240 13554 7258 13846
rect 7292 13554 7376 13846
rect 7240 12752 7376 13554
rect 7240 12460 7258 12752
rect 7292 12460 7376 12752
rect 7240 11658 7376 12460
rect 8436 13854 8572 14032
rect 8436 13562 8482 13854
rect 8516 13562 8572 13854
rect 9540 13854 9574 13870
rect 8436 12760 8572 13562
rect 8436 12468 8482 12760
rect 8516 12468 8572 12760
rect 7240 11366 7258 11658
rect 7292 11366 7376 11658
rect 7240 10564 7376 11366
rect 7828 12320 7978 12446
rect 7828 11124 7850 12320
rect 7944 11124 7978 12320
rect 7828 10800 7978 11124
rect 8436 11666 8572 12468
rect 8436 11374 8482 11666
rect 8516 11374 8572 11666
rect 7240 10272 7258 10564
rect 7292 10272 7376 10564
rect 7240 9470 7376 10272
rect 7240 9272 7258 9470
rect 6200 9162 6234 9178
rect 7234 9178 7258 9272
rect 7292 9178 7376 9470
rect 7234 9068 7376 9178
rect 8436 10572 8572 11374
rect 8436 10280 8482 10572
rect 8516 10280 8572 10572
rect 8436 9478 8572 10280
rect 8436 9186 8482 9478
rect 8516 9186 8572 9478
rect 9536 13562 9540 13760
rect 10572 13854 10640 14032
rect 10572 13766 10598 13854
rect 9574 13562 9582 13760
rect 9536 12760 9582 13562
rect 9536 12468 9540 12760
rect 9574 12468 9582 12760
rect 9536 11666 9582 12468
rect 9536 11374 9540 11666
rect 9574 11374 9582 11666
rect 9536 10572 9582 11374
rect 9536 10280 9540 10572
rect 9574 10280 9582 10572
rect 9536 9478 9582 10280
rect 9536 9398 9540 9478
rect 3006 8978 7456 9068
rect 3018 8972 7456 8978
rect 5132 8950 5214 8972
rect 4076 8216 4144 8232
rect 6200 8216 6268 8248
rect 1910 8206 6268 8216
rect 1834 8162 6268 8206
rect 1834 8126 6276 8162
rect 1834 8116 6124 8126
rect 1910 8008 2046 8116
rect 1972 7938 2040 8008
rect 1972 7646 1986 7938
rect 2020 7836 2040 7938
rect 3044 7938 3078 7954
rect 1972 7630 2020 7646
rect 3040 7646 3044 7844
rect 4076 7938 4144 8116
rect 4076 7850 4102 7938
rect 3078 7646 3086 7844
rect 1972 6860 2018 7630
rect 1972 6844 2020 6860
rect 1972 6552 1986 6844
rect 1972 6536 2020 6552
rect 3040 6844 3086 7646
rect 3040 6552 3044 6844
rect 3078 6552 3086 6844
rect 1332 6404 1482 6530
rect 1332 5208 1354 6404
rect 1448 5208 1482 6404
rect 1332 4884 1482 5208
rect 1972 5766 2018 6536
rect 1972 5750 2020 5766
rect 1972 5458 1986 5750
rect 1972 5442 2020 5458
rect 3040 5750 3086 6552
rect 3040 5458 3044 5750
rect 3078 5458 3086 5750
rect 1972 4672 2018 5442
rect 1972 4656 2020 4672
rect 1972 4364 1986 4656
rect 1972 4348 2020 4364
rect 3040 4656 3086 5458
rect 3040 4364 3044 4656
rect 3078 4364 3086 4656
rect 1972 3578 2018 4348
rect 1972 3562 2020 3578
rect 1972 3504 1986 3562
rect 3040 3562 3086 4364
rect 3040 3482 3044 3562
rect 1986 3254 2020 3270
rect 3024 3270 3044 3370
rect 3078 3482 3086 3562
rect 4092 7646 4102 7850
rect 4136 7902 4144 7938
rect 5160 7938 5194 7954
rect 4136 7850 4150 7902
rect 4136 7646 4138 7850
rect 4092 6844 4138 7646
rect 4092 6552 4102 6844
rect 4136 6552 4138 6844
rect 4092 5750 4138 6552
rect 4092 5458 4102 5750
rect 4136 5458 4138 5750
rect 4092 4656 4138 5458
rect 4092 4364 4102 4656
rect 4136 4364 4138 4656
rect 4092 3562 4138 4364
rect 4092 3504 4102 3562
rect 3078 3270 3106 3370
rect 3024 3160 3106 3270
rect 4136 3504 4138 3562
rect 6192 7938 6276 8126
rect 5194 7646 5206 7850
rect 6192 7846 6218 7938
rect 5160 6844 5206 7646
rect 5194 6552 5206 6844
rect 5160 5750 5206 6552
rect 5194 5458 5206 5750
rect 5160 4656 5206 5458
rect 5194 4364 5206 4656
rect 5160 3562 5206 4364
rect 4102 3254 4136 3270
rect 5150 3270 5160 3342
rect 5194 3488 5206 3562
rect 6212 7646 6218 7846
rect 6252 7846 6276 7938
rect 7240 7938 7376 8972
rect 8436 8224 8572 9186
rect 9520 9186 9540 9286
rect 9574 9398 9582 9478
rect 10588 13562 10598 13766
rect 10632 13818 10640 13854
rect 11656 13854 11690 13870
rect 10632 13766 10646 13818
rect 10632 13562 10634 13766
rect 10588 12760 10634 13562
rect 10588 12468 10598 12760
rect 10632 12468 10634 12760
rect 10588 11666 10634 12468
rect 10588 11374 10598 11666
rect 10632 11374 10634 11666
rect 10588 10572 10634 11374
rect 10588 10280 10598 10572
rect 10632 10280 10634 10572
rect 10588 9478 10634 10280
rect 10588 9420 10598 9478
rect 9574 9186 9602 9286
rect 9520 9076 9602 9186
rect 10632 9420 10634 9478
rect 12688 13854 12772 14042
rect 11690 13562 11702 13766
rect 12688 13762 12714 13854
rect 11656 12760 11702 13562
rect 11690 12468 11702 12760
rect 11656 11666 11702 12468
rect 11690 11374 11702 11666
rect 11656 10572 11702 11374
rect 11690 10280 11702 10572
rect 11656 9478 11702 10280
rect 10598 9170 10632 9186
rect 11646 9186 11656 9258
rect 11690 9404 11702 9478
rect 12708 13562 12714 13762
rect 12748 13762 12772 13854
rect 13768 13854 13874 14836
rect 14940 14150 15028 15050
rect 16016 15050 16036 15150
rect 16070 15262 16078 15342
rect 17084 19426 17094 19630
rect 17128 19682 17136 19718
rect 18152 19718 18186 19734
rect 17128 19630 17142 19682
rect 17128 19426 17130 19630
rect 17084 18624 17130 19426
rect 17084 18332 17094 18624
rect 17128 18332 17130 18624
rect 17084 17530 17130 18332
rect 17084 17238 17094 17530
rect 17128 17238 17130 17530
rect 17084 16436 17130 17238
rect 17084 16144 17094 16436
rect 17128 16144 17130 16436
rect 17084 15342 17130 16144
rect 17084 15284 17094 15342
rect 16070 15050 16098 15150
rect 16016 14940 16098 15050
rect 17128 15284 17130 15342
rect 19184 19718 19268 19906
rect 18186 19426 18198 19630
rect 19184 19626 19210 19718
rect 18152 18624 18198 19426
rect 18186 18332 18198 18624
rect 18152 17530 18198 18332
rect 18186 17238 18198 17530
rect 18152 16436 18198 17238
rect 18186 16144 18198 16436
rect 18152 15342 18198 16144
rect 17094 15034 17128 15050
rect 18142 15050 18152 15122
rect 18186 15268 18198 15342
rect 19204 19426 19210 19626
rect 19244 19626 19268 19718
rect 20242 19718 20336 20708
rect 21410 19980 21542 20898
rect 22506 20898 22526 20998
rect 22560 21110 22568 21190
rect 23574 25274 23584 25478
rect 23618 25530 23626 25566
rect 24642 25566 24676 25582
rect 23618 25478 23632 25530
rect 23618 25274 23620 25478
rect 23574 24472 23620 25274
rect 23574 24180 23584 24472
rect 23618 24180 23620 24472
rect 23574 23378 23620 24180
rect 23574 23086 23584 23378
rect 23618 23086 23620 23378
rect 23574 22284 23620 23086
rect 23574 21992 23584 22284
rect 23618 21992 23620 22284
rect 23574 21190 23620 21992
rect 23574 21132 23584 21190
rect 22560 20898 22588 20998
rect 22506 20788 22588 20898
rect 23618 21132 23620 21190
rect 25674 25566 25758 25754
rect 24676 25274 24688 25478
rect 25674 25474 25700 25566
rect 24642 24472 24688 25274
rect 24676 24180 24688 24472
rect 24642 23378 24688 24180
rect 24676 23086 24688 23378
rect 24642 22284 24688 23086
rect 24676 21992 24688 22284
rect 24642 21190 24688 21992
rect 23584 20882 23618 20898
rect 24632 20898 24642 20970
rect 24676 21116 24688 21190
rect 25694 25274 25700 25474
rect 25734 25474 25758 25566
rect 26740 25566 26872 26528
rect 27964 25860 28096 26750
rect 29028 26750 29048 26850
rect 29082 26962 29090 27042
rect 30096 31126 30106 31330
rect 30140 31382 30148 31418
rect 31164 31418 31198 31434
rect 30140 31330 30154 31382
rect 30140 31126 30142 31330
rect 30096 30324 30142 31126
rect 30096 30032 30106 30324
rect 30140 30032 30142 30324
rect 30096 29230 30142 30032
rect 30096 28938 30106 29230
rect 30140 28938 30142 29230
rect 30096 28136 30142 28938
rect 30096 27844 30106 28136
rect 30140 27844 30142 28136
rect 30096 27042 30142 27844
rect 30096 26984 30106 27042
rect 29082 26750 29110 26850
rect 29028 26640 29110 26750
rect 30140 26984 30142 27042
rect 32196 31418 32280 31606
rect 31198 31126 31210 31330
rect 32196 31326 32222 31418
rect 31164 30324 31210 31126
rect 31198 30032 31210 30324
rect 31164 29230 31210 30032
rect 31198 28938 31210 29230
rect 31164 28136 31210 28938
rect 31198 27844 31210 28136
rect 31164 27042 31210 27844
rect 30106 26734 30140 26750
rect 31154 26750 31164 26822
rect 31198 26968 31210 27042
rect 32216 31126 32222 31326
rect 32256 31326 32280 31418
rect 33228 31418 33360 32378
rect 34450 31702 34576 32590
rect 35538 32590 35558 32690
rect 35592 32802 35600 32882
rect 36606 36966 36616 37170
rect 36650 37222 36658 37258
rect 37674 37258 37708 37274
rect 36650 37170 36664 37222
rect 36650 36966 36652 37170
rect 36606 36164 36652 36966
rect 36606 35872 36616 36164
rect 36650 35872 36652 36164
rect 36606 35070 36652 35872
rect 36606 34778 36616 35070
rect 36650 34778 36652 35070
rect 36606 33976 36652 34778
rect 36606 33684 36616 33976
rect 36650 33684 36652 33976
rect 36606 32882 36652 33684
rect 36606 32824 36616 32882
rect 35592 32590 35620 32690
rect 35538 32480 35620 32590
rect 36650 32824 36652 32882
rect 38706 37258 38790 37446
rect 37708 36966 37720 37170
rect 38706 37166 38732 37258
rect 37674 36164 37720 36966
rect 37708 35872 37720 36164
rect 37674 35070 37720 35872
rect 37708 34778 37720 35070
rect 37674 33976 37720 34778
rect 37708 33684 37720 33976
rect 37674 32882 37720 33684
rect 36616 32574 36650 32590
rect 37664 32590 37674 32662
rect 37708 32808 37720 32882
rect 38726 36966 38732 37166
rect 38766 37166 38790 37258
rect 39768 37258 39894 38200
rect 40962 37536 41088 38406
rect 42028 38406 42048 38506
rect 42082 38618 42090 38698
rect 43096 42782 43106 42986
rect 43140 43038 43148 43074
rect 44164 43074 44198 43090
rect 43140 42986 43154 43038
rect 43140 42782 43142 42986
rect 43096 41980 43142 42782
rect 43096 41688 43106 41980
rect 43140 41688 43142 41980
rect 43096 40886 43142 41688
rect 43096 40594 43106 40886
rect 43140 40594 43142 40886
rect 43096 39792 43142 40594
rect 43096 39500 43106 39792
rect 43140 39500 43142 39792
rect 43096 38698 43142 39500
rect 43096 38640 43106 38698
rect 42082 38406 42110 38506
rect 42028 38296 42110 38406
rect 43140 38640 43142 38698
rect 45196 43074 45280 43240
rect 44198 42782 44210 42986
rect 45196 42982 45222 43074
rect 44164 41980 44210 42782
rect 44198 41688 44210 41980
rect 44164 40886 44210 41688
rect 44198 40594 44210 40886
rect 44164 39792 44210 40594
rect 44198 39500 44210 39792
rect 44164 38698 44210 39500
rect 43106 38390 43140 38406
rect 44154 38406 44164 38478
rect 44198 38624 44210 38698
rect 45216 42782 45222 42982
rect 45256 42982 45280 43074
rect 46256 43074 46386 43240
rect 45256 42782 45262 42982
rect 45216 41980 45262 42782
rect 46256 42782 46280 43074
rect 46314 42782 46386 43074
rect 46256 42554 46386 42782
rect 47564 43096 47632 43240
rect 47564 42804 47578 43096
rect 47612 42994 47632 43096
rect 48636 43096 48670 43112
rect 47564 42788 47612 42804
rect 48632 42804 48636 43002
rect 49668 43096 49736 43274
rect 51778 43262 54496 43284
rect 49668 43008 49694 43096
rect 48670 42804 48678 43002
rect 45216 41688 45222 41980
rect 45256 41688 45262 41980
rect 45216 40886 45262 41688
rect 45216 40594 45222 40886
rect 45256 40594 45262 40886
rect 45216 39792 45262 40594
rect 45216 39500 45222 39792
rect 45256 39500 45262 39792
rect 45216 38698 45262 39500
rect 45216 38668 45222 38698
rect 44198 38406 44236 38478
rect 44154 38296 44236 38406
rect 45256 38668 45262 38698
rect 46272 41980 46318 42554
rect 46272 41688 46280 41980
rect 46314 41688 46318 41980
rect 47564 42018 47610 42788
rect 47564 42002 47612 42018
rect 47564 41710 47578 42002
rect 47564 41694 47612 41710
rect 48632 42002 48678 42804
rect 48632 41710 48636 42002
rect 48670 41710 48678 42002
rect 46272 40886 46318 41688
rect 46272 40594 46280 40886
rect 46314 40594 46318 40886
rect 46272 39792 46318 40594
rect 46924 41562 47074 41688
rect 46924 40366 46946 41562
rect 47040 40366 47074 41562
rect 46924 40042 47074 40366
rect 47564 40924 47610 41694
rect 47564 40908 47612 40924
rect 47564 40616 47578 40908
rect 47564 40600 47612 40616
rect 48632 40908 48678 41710
rect 48632 40616 48636 40908
rect 48670 40616 48678 40908
rect 46272 39500 46280 39792
rect 46314 39500 46318 39792
rect 46272 38698 46318 39500
rect 46272 38640 46280 38698
rect 45222 38390 45256 38406
rect 46242 38406 46280 38512
rect 46314 38640 46318 38698
rect 47564 39830 47610 40600
rect 47564 39814 47612 39830
rect 47564 39522 47578 39814
rect 47564 39506 47612 39522
rect 48632 39814 48678 40616
rect 48632 39522 48636 39814
rect 48670 39522 48678 39814
rect 47564 38736 47610 39506
rect 47564 38720 47612 38736
rect 47564 38662 47578 38720
rect 46314 38406 46368 38512
rect 46242 38296 46368 38406
rect 47548 38428 47578 38604
rect 48632 38720 48678 39522
rect 48632 38640 48636 38720
rect 47612 38428 47680 38604
rect 42028 38206 46478 38296
rect 42040 38200 46478 38206
rect 44154 38178 44236 38200
rect 43080 37536 43148 37552
rect 45204 37536 45272 37568
rect 40962 37526 45272 37536
rect 40838 37482 45272 37526
rect 40838 37446 45280 37482
rect 40838 37436 45128 37446
rect 38766 36966 38772 37166
rect 39768 37112 39790 37258
rect 38726 36164 38772 36966
rect 38726 35872 38732 36164
rect 38766 35872 38772 36164
rect 38726 35070 38772 35872
rect 38726 34778 38732 35070
rect 38766 34778 38772 35070
rect 38726 33976 38772 34778
rect 38726 33684 38732 33976
rect 38766 33684 38772 33976
rect 38726 32882 38772 33684
rect 38726 32852 38732 32882
rect 37708 32590 37746 32662
rect 37664 32480 37746 32590
rect 38766 32852 38772 32882
rect 39782 36966 39790 37112
rect 39824 37112 39894 37258
rect 40962 37258 41088 37436
rect 40962 37212 40990 37258
rect 39824 36966 39828 37112
rect 39782 36164 39828 36966
rect 39782 35872 39790 36164
rect 39824 35872 39828 36164
rect 39782 35070 39828 35872
rect 40976 36966 40990 37212
rect 41024 37212 41088 37258
rect 42048 37258 42082 37274
rect 41024 37156 41044 37212
rect 40976 36950 41024 36966
rect 42044 36966 42048 37164
rect 43080 37258 43148 37436
rect 43080 37170 43106 37258
rect 42082 36966 42090 37164
rect 40976 36180 41022 36950
rect 40976 36164 41024 36180
rect 40976 35872 40990 36164
rect 40976 35856 41024 35872
rect 42044 36164 42090 36966
rect 42044 35872 42048 36164
rect 42082 35872 42090 36164
rect 39782 34778 39790 35070
rect 39824 34778 39828 35070
rect 39782 33976 39828 34778
rect 40336 35724 40486 35850
rect 40336 34528 40358 35724
rect 40452 34528 40486 35724
rect 40336 34204 40486 34528
rect 40976 35086 41022 35856
rect 40976 35070 41024 35086
rect 40976 34778 40990 35070
rect 40976 34762 41024 34778
rect 42044 35070 42090 35872
rect 42044 34778 42048 35070
rect 42082 34778 42090 35070
rect 39782 33684 39790 33976
rect 39824 33684 39828 33976
rect 39782 32882 39828 33684
rect 39782 32824 39790 32882
rect 38732 32574 38766 32590
rect 39754 32590 39790 32716
rect 39824 32824 39828 32882
rect 40976 33992 41022 34762
rect 40976 33976 41024 33992
rect 40976 33684 40990 33976
rect 40976 33668 41024 33684
rect 42044 33976 42090 34778
rect 42044 33684 42048 33976
rect 42082 33684 42090 33976
rect 40976 32898 41022 33668
rect 40976 32882 41024 32898
rect 40976 32824 40990 32882
rect 39824 32590 39880 32716
rect 39754 32480 39880 32590
rect 40962 32590 40990 32702
rect 42044 32882 42090 33684
rect 42044 32802 42048 32882
rect 41024 32590 41088 32702
rect 35538 32390 39988 32480
rect 35550 32384 39988 32390
rect 37664 32362 37746 32384
rect 36590 31702 36658 31718
rect 38714 31702 38782 31734
rect 34450 31692 38782 31702
rect 34348 31648 38782 31692
rect 34348 31612 38790 31648
rect 34348 31602 38638 31612
rect 32256 31126 32262 31326
rect 33228 31232 33280 31418
rect 32216 30324 32262 31126
rect 32216 30032 32222 30324
rect 32256 30032 32262 30324
rect 32216 29230 32262 30032
rect 32216 28938 32222 29230
rect 32256 28938 32262 29230
rect 32216 28136 32262 28938
rect 32216 27844 32222 28136
rect 32256 27844 32262 28136
rect 32216 27042 32262 27844
rect 32216 27012 32222 27042
rect 31198 26750 31236 26822
rect 31154 26640 31236 26750
rect 32256 27012 32262 27042
rect 33272 31126 33280 31232
rect 33314 31232 33360 31418
rect 34450 31424 34576 31602
rect 34450 31388 34500 31424
rect 33314 31126 33318 31232
rect 33272 30324 33318 31126
rect 33272 30032 33280 30324
rect 33314 30032 33318 30324
rect 33272 29230 33318 30032
rect 34486 31132 34500 31388
rect 34534 31388 34576 31424
rect 35558 31424 35592 31440
rect 34534 31322 34554 31388
rect 34486 31116 34534 31132
rect 35554 31132 35558 31330
rect 36590 31424 36658 31602
rect 36590 31336 36616 31424
rect 35592 31132 35600 31330
rect 34486 30346 34532 31116
rect 34486 30330 34534 30346
rect 34486 30038 34500 30330
rect 34486 30022 34534 30038
rect 35554 30330 35600 31132
rect 35554 30038 35558 30330
rect 35592 30038 35600 30330
rect 33272 28938 33280 29230
rect 33314 28938 33318 29230
rect 33272 28136 33318 28938
rect 33846 29890 33996 30016
rect 33846 28694 33868 29890
rect 33962 28694 33996 29890
rect 33846 28370 33996 28694
rect 34486 29252 34532 30022
rect 34486 29236 34534 29252
rect 34486 28944 34500 29236
rect 34486 28928 34534 28944
rect 35554 29236 35600 30038
rect 35554 28944 35558 29236
rect 35592 28944 35600 29236
rect 33272 27844 33280 28136
rect 33314 27844 33318 28136
rect 33272 27042 33318 27844
rect 33272 26984 33280 27042
rect 32222 26734 32256 26750
rect 33256 26750 33280 26844
rect 33314 26984 33318 27042
rect 34486 28158 34532 28928
rect 34486 28142 34534 28158
rect 34486 27850 34500 28142
rect 34486 27834 34534 27850
rect 35554 28142 35600 28944
rect 35554 27850 35558 28142
rect 35592 27850 35600 28142
rect 34486 27064 34532 27834
rect 34486 27048 34534 27064
rect 34486 26990 34500 27048
rect 33314 26824 33338 26844
rect 33314 26750 33384 26824
rect 33256 26640 33384 26750
rect 34450 26756 34500 26936
rect 35554 27048 35600 27850
rect 35554 26968 35558 27048
rect 34534 26756 34576 26936
rect 29028 26550 33478 26640
rect 29040 26544 33478 26550
rect 31154 26522 31236 26544
rect 30080 25860 30148 25876
rect 32204 25860 32272 25892
rect 27964 25850 32272 25860
rect 27838 25806 32272 25850
rect 27838 25770 32280 25806
rect 27838 25760 32128 25770
rect 27964 25672 28096 25760
rect 25734 25274 25740 25474
rect 26740 25470 26758 25566
rect 25694 24472 25740 25274
rect 25694 24180 25700 24472
rect 25734 24180 25740 24472
rect 25694 23378 25740 24180
rect 25694 23086 25700 23378
rect 25734 23086 25740 23378
rect 25694 22284 25740 23086
rect 25694 21992 25700 22284
rect 25734 21992 25740 22284
rect 25694 21190 25740 21992
rect 25694 21160 25700 21190
rect 24676 20898 24714 20970
rect 24632 20788 24714 20898
rect 25734 21160 25740 21190
rect 26750 25274 26758 25470
rect 26792 25470 26872 25566
rect 27976 25582 28044 25672
rect 26792 25274 26796 25470
rect 26750 24472 26796 25274
rect 26750 24180 26758 24472
rect 26792 24180 26796 24472
rect 26750 23378 26796 24180
rect 27976 25290 27990 25582
rect 28024 25480 28044 25582
rect 29048 25582 29082 25598
rect 27976 25274 28024 25290
rect 29044 25290 29048 25488
rect 30080 25582 30148 25760
rect 30080 25494 30106 25582
rect 29082 25290 29090 25488
rect 27976 24504 28022 25274
rect 27976 24488 28024 24504
rect 27976 24196 27990 24488
rect 27976 24180 28024 24196
rect 29044 24488 29090 25290
rect 29044 24196 29048 24488
rect 29082 24196 29090 24488
rect 26750 23086 26758 23378
rect 26792 23086 26796 23378
rect 26750 22284 26796 23086
rect 27336 24048 27486 24174
rect 27336 22852 27358 24048
rect 27452 22852 27486 24048
rect 27336 22528 27486 22852
rect 27976 23410 28022 24180
rect 27976 23394 28024 23410
rect 27976 23102 27990 23394
rect 27976 23086 28024 23102
rect 29044 23394 29090 24196
rect 29044 23102 29048 23394
rect 29082 23102 29090 23394
rect 26750 21992 26758 22284
rect 26792 21992 26796 22284
rect 26750 21190 26796 21992
rect 27976 22316 28022 23086
rect 27976 22300 28024 22316
rect 27976 22008 27990 22300
rect 27976 21992 28024 22008
rect 29044 22300 29090 23102
rect 29044 22008 29048 22300
rect 29082 22008 29090 22300
rect 27976 21258 28022 21992
rect 26750 21132 26758 21190
rect 25700 20882 25734 20898
rect 26688 20898 26758 21004
rect 26792 21132 26796 21190
rect 27926 21206 28058 21258
rect 26792 20898 26820 21004
rect 26688 20788 26820 20898
rect 27926 20914 27990 21206
rect 28024 20914 28058 21206
rect 29044 21206 29090 22008
rect 29044 21126 29048 21206
rect 22506 20698 26956 20788
rect 22518 20692 26956 20698
rect 24632 20670 24714 20692
rect 23558 19980 23626 19996
rect 25682 19980 25750 20012
rect 21410 19970 25750 19980
rect 21316 19926 25750 19970
rect 21316 19890 25758 19926
rect 21316 19880 25606 19890
rect 19244 19426 19250 19626
rect 19204 18624 19250 19426
rect 19204 18332 19210 18624
rect 19244 18332 19250 18624
rect 19204 17530 19250 18332
rect 19204 17238 19210 17530
rect 19244 17238 19250 17530
rect 19204 16436 19250 17238
rect 19204 16144 19210 16436
rect 19244 16144 19250 16436
rect 19204 15342 19250 16144
rect 19204 15312 19210 15342
rect 18186 15050 18224 15122
rect 18142 14940 18224 15050
rect 19244 15312 19250 15342
rect 20242 19426 20268 19718
rect 20302 19426 20336 19718
rect 21410 19702 21542 19880
rect 21410 19692 21468 19702
rect 20242 18624 20336 19426
rect 20242 18332 20268 18624
rect 20302 18332 20336 18624
rect 20242 17530 20336 18332
rect 21454 19410 21468 19692
rect 21502 19692 21542 19702
rect 22526 19702 22560 19718
rect 21502 19600 21522 19692
rect 21454 19394 21502 19410
rect 22522 19410 22526 19608
rect 23558 19702 23626 19880
rect 23558 19614 23584 19702
rect 22560 19410 22568 19608
rect 21454 18624 21500 19394
rect 21454 18608 21502 18624
rect 21454 18316 21468 18608
rect 21454 18300 21502 18316
rect 22522 18608 22568 19410
rect 22522 18316 22526 18608
rect 22560 18316 22568 18608
rect 20242 17238 20268 17530
rect 20302 17238 20336 17530
rect 20242 16436 20336 17238
rect 20814 18168 20964 18294
rect 20814 16972 20836 18168
rect 20930 16972 20964 18168
rect 20814 16648 20964 16972
rect 21454 17530 21500 18300
rect 21454 17514 21502 17530
rect 21454 17222 21468 17514
rect 21454 17206 21502 17222
rect 22522 17514 22568 18316
rect 22522 17222 22526 17514
rect 22560 17222 22568 17514
rect 20242 16144 20268 16436
rect 20302 16144 20336 16436
rect 20242 15342 20336 16144
rect 19210 15034 19244 15050
rect 20242 15050 20268 15342
rect 20302 15050 20336 15342
rect 21454 16436 21500 17206
rect 21454 16420 21502 16436
rect 21454 16128 21468 16420
rect 21454 16112 21502 16128
rect 22522 16420 22568 17222
rect 22522 16128 22526 16420
rect 22560 16128 22568 16420
rect 21454 15342 21500 16112
rect 21454 15330 21502 15342
rect 20242 14940 20336 15050
rect 21440 15326 21572 15330
rect 21440 15034 21468 15326
rect 21502 15034 21572 15326
rect 22522 15326 22568 16128
rect 22522 15246 22526 15326
rect 16016 14850 20466 14940
rect 16028 14844 20466 14850
rect 18142 14822 18224 14844
rect 14940 14140 15042 14150
rect 17078 14140 17146 14156
rect 19202 14140 19270 14172
rect 14940 14130 19270 14140
rect 14836 14086 19270 14130
rect 14836 14050 19278 14086
rect 14836 14040 19126 14050
rect 13768 13782 13772 13854
rect 12748 13562 12754 13762
rect 12708 12760 12754 13562
rect 12708 12468 12714 12760
rect 12748 12468 12754 12760
rect 12708 11666 12754 12468
rect 12708 11374 12714 11666
rect 12748 11374 12754 11666
rect 12708 10572 12754 11374
rect 12708 10280 12714 10572
rect 12748 10280 12754 10572
rect 12708 9478 12754 10280
rect 12708 9448 12714 9478
rect 11690 9186 11728 9258
rect 11646 9076 11728 9186
rect 12748 9448 12754 9478
rect 13764 13562 13772 13782
rect 13806 13562 13874 13854
rect 13764 12760 13874 13562
rect 13764 12468 13772 12760
rect 13806 12468 13874 12760
rect 13764 11666 13874 12468
rect 14940 13862 15042 14040
rect 14940 13570 14988 13862
rect 15022 13760 15042 13862
rect 16046 13862 16080 13878
rect 15022 13570 15028 13760
rect 14940 12768 15028 13570
rect 14940 12476 14988 12768
rect 15022 12476 15028 12768
rect 13764 11374 13772 11666
rect 13806 11374 13874 11666
rect 13764 10572 13874 11374
rect 14334 12328 14484 12454
rect 14334 11132 14356 12328
rect 14450 11132 14484 12328
rect 14334 10808 14484 11132
rect 14940 11674 15028 12476
rect 14940 11382 14988 11674
rect 15022 11382 15028 11674
rect 13764 10280 13772 10572
rect 13806 10280 13874 10572
rect 13764 9478 13874 10280
rect 13764 9420 13772 9478
rect 13768 9280 13772 9420
rect 12714 9170 12748 9186
rect 13748 9186 13772 9280
rect 13806 9186 13874 9478
rect 13748 9076 13874 9186
rect 14940 10580 15028 11382
rect 14940 10288 14988 10580
rect 15022 10288 15028 10580
rect 14940 9486 15028 10288
rect 14940 9194 14988 9486
rect 15022 9240 15028 9486
rect 16042 13570 16046 13768
rect 17078 13862 17146 14040
rect 17078 13774 17104 13862
rect 16080 13570 16088 13768
rect 16042 12768 16088 13570
rect 16042 12476 16046 12768
rect 16080 12476 16088 12768
rect 16042 11674 16088 12476
rect 16042 11382 16046 11674
rect 16080 11382 16088 11674
rect 16042 10580 16088 11382
rect 16042 10288 16046 10580
rect 16080 10288 16088 10580
rect 16042 9486 16088 10288
rect 16042 9406 16046 9486
rect 15022 9194 15072 9240
rect 9520 8986 13970 9076
rect 9532 8980 13970 8986
rect 11646 8958 11728 8980
rect 10590 8224 10658 8240
rect 12714 8224 12782 8256
rect 8436 8214 12782 8224
rect 8348 8170 12782 8214
rect 8348 8134 12790 8170
rect 8348 8124 12638 8134
rect 6252 7646 6258 7846
rect 7240 7772 7276 7938
rect 6212 6844 6258 7646
rect 6212 6552 6218 6844
rect 6252 6552 6258 6844
rect 6212 5750 6258 6552
rect 6212 5458 6218 5750
rect 6252 5458 6258 5750
rect 6212 4656 6258 5458
rect 6212 4364 6218 4656
rect 6252 4364 6258 4656
rect 6212 3562 6258 4364
rect 6212 3532 6218 3562
rect 5194 3270 5232 3342
rect 5150 3160 5232 3270
rect 6252 3532 6258 3562
rect 7268 7646 7276 7772
rect 7310 7772 7376 7938
rect 8436 7946 8572 8124
rect 7310 7646 7314 7772
rect 8436 7688 8500 7946
rect 7268 6844 7314 7646
rect 7268 6552 7276 6844
rect 7310 6552 7314 6844
rect 7268 5750 7314 6552
rect 8486 7654 8500 7688
rect 8534 7688 8572 7946
rect 9558 7946 9592 7962
rect 8486 7638 8534 7654
rect 9554 7654 9558 7852
rect 10590 7946 10658 8124
rect 10590 7858 10616 7946
rect 9592 7654 9600 7852
rect 8486 6868 8532 7638
rect 8486 6852 8534 6868
rect 8486 6560 8500 6852
rect 8486 6544 8534 6560
rect 9554 6852 9600 7654
rect 9554 6560 9558 6852
rect 9592 6560 9600 6852
rect 7268 5458 7276 5750
rect 7310 5458 7314 5750
rect 7268 4656 7314 5458
rect 7846 6412 7996 6538
rect 7846 5216 7868 6412
rect 7962 5216 7996 6412
rect 7846 4892 7996 5216
rect 8486 5774 8532 6544
rect 8486 5758 8534 5774
rect 8486 5466 8500 5758
rect 8486 5450 8534 5466
rect 9554 5758 9600 6560
rect 9554 5466 9558 5758
rect 9592 5466 9600 5758
rect 7268 4364 7276 4656
rect 7310 4364 7314 4656
rect 7268 3562 7314 4364
rect 7268 3504 7276 3562
rect 6218 3254 6252 3270
rect 7252 3270 7276 3364
rect 7310 3504 7314 3562
rect 8486 4680 8532 5450
rect 8486 4664 8534 4680
rect 8486 4372 8500 4664
rect 8486 4356 8534 4372
rect 9554 4664 9600 5466
rect 9554 4372 9558 4664
rect 9592 4372 9600 4664
rect 8486 3586 8532 4356
rect 8486 3570 8534 3586
rect 8486 3512 8500 3570
rect 7310 3270 7334 3364
rect 7252 3160 7334 3270
rect 9554 3570 9600 4372
rect 9554 3490 9558 3570
rect 8500 3262 8534 3278
rect 9538 3278 9558 3378
rect 9592 3490 9600 3570
rect 10606 7654 10616 7858
rect 10650 7910 10658 7946
rect 11674 7946 11708 7962
rect 10650 7858 10664 7910
rect 10650 7654 10652 7858
rect 10606 6852 10652 7654
rect 10606 6560 10616 6852
rect 10650 6560 10652 6852
rect 10606 5758 10652 6560
rect 10606 5466 10616 5758
rect 10650 5466 10652 5758
rect 10606 4664 10652 5466
rect 10606 4372 10616 4664
rect 10650 4372 10652 4664
rect 10606 3570 10652 4372
rect 10606 3512 10616 3570
rect 9592 3278 9620 3378
rect 9538 3168 9620 3278
rect 10650 3512 10652 3570
rect 12706 7946 12790 8134
rect 11708 7654 11720 7858
rect 12706 7854 12732 7946
rect 11674 6852 11720 7654
rect 11708 6560 11720 6852
rect 11674 5758 11720 6560
rect 11708 5466 11720 5758
rect 11674 4664 11720 5466
rect 11708 4372 11720 4664
rect 11674 3570 11720 4372
rect 10616 3262 10650 3278
rect 11664 3278 11674 3350
rect 11708 3496 11720 3570
rect 12726 7654 12732 7854
rect 12766 7854 12790 7946
rect 13768 7946 13874 8980
rect 14940 8232 15072 9194
rect 16026 9194 16046 9294
rect 16080 9406 16088 9486
rect 17094 13570 17104 13774
rect 17138 13826 17146 13862
rect 18162 13862 18196 13878
rect 17138 13774 17152 13826
rect 17138 13570 17140 13774
rect 17094 12768 17140 13570
rect 17094 12476 17104 12768
rect 17138 12476 17140 12768
rect 17094 11674 17140 12476
rect 17094 11382 17104 11674
rect 17138 11382 17140 11674
rect 17094 10580 17140 11382
rect 17094 10288 17104 10580
rect 17138 10288 17140 10580
rect 17094 9486 17140 10288
rect 17094 9428 17104 9486
rect 16080 9194 16108 9294
rect 16026 9084 16108 9194
rect 17138 9428 17140 9486
rect 19194 13862 19278 14050
rect 18196 13570 18208 13774
rect 19194 13770 19220 13862
rect 18162 12768 18208 13570
rect 18196 12476 18208 12768
rect 18162 11674 18208 12476
rect 18196 11382 18208 11674
rect 18162 10580 18208 11382
rect 18196 10288 18208 10580
rect 18162 9486 18208 10288
rect 17104 9178 17138 9194
rect 18152 9194 18162 9266
rect 18196 9412 18208 9486
rect 19214 13570 19220 13770
rect 19254 13770 19278 13862
rect 20242 13862 20336 14844
rect 21440 14124 21572 15034
rect 22506 15034 22526 15134
rect 22560 15246 22568 15326
rect 23574 19410 23584 19614
rect 23618 19666 23626 19702
rect 24642 19702 24676 19718
rect 23618 19614 23632 19666
rect 23618 19410 23620 19614
rect 23574 18608 23620 19410
rect 23574 18316 23584 18608
rect 23618 18316 23620 18608
rect 23574 17514 23620 18316
rect 23574 17222 23584 17514
rect 23618 17222 23620 17514
rect 23574 16420 23620 17222
rect 23574 16128 23584 16420
rect 23618 16128 23620 16420
rect 23574 15326 23620 16128
rect 23574 15268 23584 15326
rect 22560 15034 22588 15134
rect 22506 14924 22588 15034
rect 23618 15268 23620 15326
rect 25674 19702 25758 19890
rect 24676 19410 24688 19614
rect 25674 19610 25700 19702
rect 24642 18608 24688 19410
rect 24676 18316 24688 18608
rect 24642 17514 24688 18316
rect 24676 17222 24688 17514
rect 24642 16420 24688 17222
rect 24676 16128 24688 16420
rect 24642 15326 24688 16128
rect 23584 15018 23618 15034
rect 24632 15034 24642 15106
rect 24676 15252 24688 15326
rect 25694 19410 25700 19610
rect 25734 19610 25758 19702
rect 26688 19702 26820 20692
rect 27926 19996 28058 20914
rect 29028 20914 29048 21014
rect 29082 21126 29090 21206
rect 30096 25290 30106 25494
rect 30140 25546 30148 25582
rect 31164 25582 31198 25598
rect 30140 25494 30154 25546
rect 30140 25290 30142 25494
rect 30096 24488 30142 25290
rect 30096 24196 30106 24488
rect 30140 24196 30142 24488
rect 30096 23394 30142 24196
rect 30096 23102 30106 23394
rect 30140 23102 30142 23394
rect 30096 22300 30142 23102
rect 30096 22008 30106 22300
rect 30140 22008 30142 22300
rect 30096 21206 30142 22008
rect 30096 21148 30106 21206
rect 29082 20914 29110 21014
rect 29028 20804 29110 20914
rect 30140 21148 30142 21206
rect 32196 25582 32280 25770
rect 31198 25290 31210 25494
rect 32196 25490 32222 25582
rect 31164 24488 31210 25290
rect 31198 24196 31210 24488
rect 31164 23394 31210 24196
rect 31198 23102 31210 23394
rect 31164 22300 31210 23102
rect 31198 22008 31210 22300
rect 31164 21206 31210 22008
rect 30106 20898 30140 20914
rect 31154 20914 31164 20986
rect 31198 21132 31210 21206
rect 32216 25290 32222 25490
rect 32256 25490 32280 25582
rect 33258 25582 33384 26544
rect 34450 25866 34576 26756
rect 35538 26756 35558 26856
rect 35592 26968 35600 27048
rect 36606 31132 36616 31336
rect 36650 31388 36658 31424
rect 37674 31424 37708 31440
rect 36650 31336 36664 31388
rect 36650 31132 36652 31336
rect 36606 30330 36652 31132
rect 36606 30038 36616 30330
rect 36650 30038 36652 30330
rect 36606 29236 36652 30038
rect 36606 28944 36616 29236
rect 36650 28944 36652 29236
rect 36606 28142 36652 28944
rect 36606 27850 36616 28142
rect 36650 27850 36652 28142
rect 36606 27048 36652 27850
rect 36606 26990 36616 27048
rect 35592 26756 35620 26856
rect 35538 26646 35620 26756
rect 36650 26990 36652 27048
rect 38706 31424 38790 31612
rect 37708 31132 37720 31336
rect 38706 31332 38732 31424
rect 37674 30330 37720 31132
rect 37708 30038 37720 30330
rect 37674 29236 37720 30038
rect 37708 28944 37720 29236
rect 37674 28142 37720 28944
rect 37708 27850 37720 28142
rect 37674 27048 37720 27850
rect 36616 26740 36650 26756
rect 37664 26756 37674 26828
rect 37708 26974 37720 27048
rect 38726 31132 38732 31332
rect 38766 31332 38790 31424
rect 39754 31424 39880 32384
rect 40962 31702 41088 32590
rect 42028 32590 42048 32690
rect 42082 32802 42090 32882
rect 43096 36966 43106 37170
rect 43140 37222 43148 37258
rect 44164 37258 44198 37274
rect 43140 37170 43154 37222
rect 43140 36966 43142 37170
rect 43096 36164 43142 36966
rect 43096 35872 43106 36164
rect 43140 35872 43142 36164
rect 43096 35070 43142 35872
rect 43096 34778 43106 35070
rect 43140 34778 43142 35070
rect 43096 33976 43142 34778
rect 43096 33684 43106 33976
rect 43140 33684 43142 33976
rect 43096 32882 43142 33684
rect 43096 32824 43106 32882
rect 42082 32590 42110 32690
rect 42028 32480 42110 32590
rect 43140 32824 43142 32882
rect 45196 37258 45280 37446
rect 44198 36966 44210 37170
rect 45196 37166 45222 37258
rect 44164 36164 44210 36966
rect 44198 35872 44210 36164
rect 44164 35070 44210 35872
rect 44198 34778 44210 35070
rect 44164 33976 44210 34778
rect 44198 33684 44210 33976
rect 44164 32882 44210 33684
rect 43106 32574 43140 32590
rect 44154 32590 44164 32662
rect 44198 32808 44210 32882
rect 45216 36966 45222 37166
rect 45256 37166 45280 37258
rect 46242 37258 46368 38200
rect 47548 37558 47680 38428
rect 48616 38428 48636 38528
rect 48670 38640 48678 38720
rect 49684 42804 49694 43008
rect 49728 43060 49736 43096
rect 50752 43096 50786 43112
rect 49728 43008 49742 43060
rect 49728 42804 49730 43008
rect 49684 42002 49730 42804
rect 49684 41710 49694 42002
rect 49728 41710 49730 42002
rect 49684 40908 49730 41710
rect 49684 40616 49694 40908
rect 49728 40616 49730 40908
rect 49684 39814 49730 40616
rect 49684 39522 49694 39814
rect 49728 39522 49730 39814
rect 49684 38720 49730 39522
rect 49684 38662 49694 38720
rect 48670 38428 48698 38528
rect 48616 38318 48698 38428
rect 49728 38662 49730 38720
rect 51784 43096 51868 43262
rect 50786 42804 50798 43008
rect 51784 43004 51810 43096
rect 50752 42002 50798 42804
rect 50786 41710 50798 42002
rect 50752 40908 50798 41710
rect 50786 40616 50798 40908
rect 50752 39814 50798 40616
rect 50786 39522 50798 39814
rect 50752 38720 50798 39522
rect 49694 38412 49728 38428
rect 50742 38428 50752 38500
rect 50786 38646 50798 38720
rect 51804 42804 51810 43004
rect 51844 43004 51868 43096
rect 52830 43096 52960 43262
rect 51844 42804 51850 43004
rect 51804 42002 51850 42804
rect 52830 42804 52868 43096
rect 52902 42804 52960 43096
rect 52830 42574 52960 42804
rect 54078 43110 54146 43262
rect 54078 42818 54092 43110
rect 54126 43008 54146 43110
rect 55150 43110 55184 43126
rect 54078 42802 54126 42818
rect 55146 42818 55150 43016
rect 56182 43110 56250 43288
rect 58296 43198 59446 43298
rect 62498 43284 62560 43294
rect 56182 43022 56208 43110
rect 55184 42818 55192 43016
rect 51804 41710 51810 42002
rect 51844 41710 51850 42002
rect 51804 40908 51850 41710
rect 51804 40616 51810 40908
rect 51844 40616 51850 40908
rect 51804 39814 51850 40616
rect 51804 39522 51810 39814
rect 51844 39522 51850 39814
rect 51804 38720 51850 39522
rect 51804 38690 51810 38720
rect 50786 38428 50824 38500
rect 50742 38318 50824 38428
rect 51844 38690 51850 38720
rect 52860 42002 52906 42574
rect 52860 41710 52868 42002
rect 52902 41710 52906 42002
rect 52860 40908 52906 41710
rect 54078 42032 54124 42802
rect 54078 42016 54126 42032
rect 54078 41724 54092 42016
rect 54078 41708 54126 41724
rect 55146 42016 55192 42818
rect 55146 41724 55150 42016
rect 55184 41724 55192 42016
rect 52860 40616 52868 40908
rect 52902 40616 52906 40908
rect 52860 39814 52906 40616
rect 53438 41576 53588 41702
rect 53438 40380 53460 41576
rect 53554 40380 53588 41576
rect 53438 40056 53588 40380
rect 54078 40938 54124 41708
rect 54078 40922 54126 40938
rect 54078 40630 54092 40922
rect 54078 40614 54126 40630
rect 55146 40922 55192 41724
rect 55146 40630 55150 40922
rect 55184 40630 55192 40922
rect 52860 39522 52868 39814
rect 52902 39522 52906 39814
rect 52860 38720 52906 39522
rect 52860 38662 52868 38720
rect 52850 38522 52868 38536
rect 51810 38412 51844 38428
rect 52844 38428 52868 38522
rect 52902 38662 52906 38720
rect 54078 39844 54124 40614
rect 54078 39828 54126 39844
rect 54078 39536 54092 39828
rect 54078 39520 54126 39536
rect 55146 39828 55192 40630
rect 55146 39536 55150 39828
rect 55184 39536 55192 39828
rect 54078 38750 54124 39520
rect 54078 38734 54126 38750
rect 54078 38676 54092 38734
rect 52902 38428 52946 38536
rect 52844 38318 52946 38428
rect 54062 38442 54092 38602
rect 55146 38734 55192 39536
rect 55146 38654 55150 38734
rect 54126 38442 54158 38602
rect 48616 38228 53066 38318
rect 48628 38222 53066 38228
rect 50742 38200 50824 38222
rect 49668 37558 49736 37574
rect 51792 37558 51860 37590
rect 47548 37548 51860 37558
rect 47426 37504 51860 37548
rect 47426 37468 51868 37504
rect 47426 37458 51716 37468
rect 45256 36966 45262 37166
rect 46242 37128 46280 37258
rect 45216 36164 45262 36966
rect 45216 35872 45222 36164
rect 45256 35872 45262 36164
rect 45216 35070 45262 35872
rect 45216 34778 45222 35070
rect 45256 34778 45262 35070
rect 45216 33976 45262 34778
rect 45216 33684 45222 33976
rect 45256 33684 45262 33976
rect 45216 32882 45262 33684
rect 45216 32852 45222 32882
rect 44198 32590 44236 32662
rect 44154 32480 44236 32590
rect 45256 32852 45262 32882
rect 46272 36966 46280 37128
rect 46314 37128 46368 37258
rect 47548 37280 47680 37458
rect 47548 37196 47578 37280
rect 46314 36966 46318 37128
rect 46272 36164 46318 36966
rect 46272 35872 46280 36164
rect 46314 35872 46318 36164
rect 47564 36988 47578 37196
rect 47612 37196 47680 37280
rect 48636 37280 48670 37296
rect 47612 37178 47632 37196
rect 47564 36972 47612 36988
rect 48632 36988 48636 37186
rect 49668 37280 49736 37458
rect 49668 37192 49694 37280
rect 48670 36988 48678 37186
rect 47564 36202 47610 36972
rect 47564 36186 47612 36202
rect 47564 35894 47578 36186
rect 47564 35878 47612 35894
rect 48632 36186 48678 36988
rect 48632 35894 48636 36186
rect 48670 35894 48678 36186
rect 46272 35070 46318 35872
rect 46272 34778 46280 35070
rect 46314 34778 46318 35070
rect 46272 33976 46318 34778
rect 46924 35746 47074 35872
rect 46924 34550 46946 35746
rect 47040 34550 47074 35746
rect 46924 34226 47074 34550
rect 47564 35108 47610 35878
rect 47564 35092 47612 35108
rect 47564 34800 47578 35092
rect 47564 34784 47612 34800
rect 48632 35092 48678 35894
rect 48632 34800 48636 35092
rect 48670 34800 48678 35092
rect 46272 33684 46280 33976
rect 46314 33684 46318 33976
rect 46272 32882 46318 33684
rect 46272 32824 46280 32882
rect 46256 32632 46280 32684
rect 45222 32574 45256 32590
rect 46242 32590 46280 32632
rect 46314 32824 46318 32882
rect 47564 34014 47610 34784
rect 47564 33998 47612 34014
rect 47564 33706 47578 33998
rect 47564 33690 47612 33706
rect 48632 33998 48678 34800
rect 48632 33706 48636 33998
rect 48670 33706 48678 33998
rect 47564 32920 47610 33690
rect 47564 32904 47612 32920
rect 47564 32846 47578 32904
rect 46314 32632 46338 32684
rect 46314 32590 46368 32632
rect 46242 32480 46368 32590
rect 47524 32612 47578 32790
rect 48632 32904 48678 33706
rect 48632 32824 48636 32904
rect 47612 32612 47656 32790
rect 42028 32390 46478 32480
rect 42040 32384 46478 32390
rect 44154 32362 44236 32384
rect 43080 31702 43148 31718
rect 45204 31702 45272 31734
rect 40962 31692 45272 31702
rect 40838 31648 45272 31692
rect 40838 31612 45280 31648
rect 40838 31602 45128 31612
rect 39754 31332 39790 31424
rect 38766 31132 38772 31332
rect 38726 30330 38772 31132
rect 38726 30038 38732 30330
rect 38766 30038 38772 30330
rect 38726 29236 38772 30038
rect 38726 28944 38732 29236
rect 38766 28944 38772 29236
rect 38726 28142 38772 28944
rect 38726 27850 38732 28142
rect 38766 27850 38772 28142
rect 38726 27048 38772 27850
rect 38726 27018 38732 27048
rect 37708 26756 37746 26828
rect 37664 26646 37746 26756
rect 38766 27018 38772 27048
rect 39782 31132 39790 31332
rect 39824 31332 39880 31424
rect 40962 31424 41088 31602
rect 39824 31132 39828 31332
rect 40962 31318 40990 31424
rect 39782 30330 39828 31132
rect 39782 30038 39790 30330
rect 39824 30038 39828 30330
rect 39782 29236 39828 30038
rect 40976 31132 40990 31318
rect 41024 31318 41088 31424
rect 42048 31424 42082 31440
rect 40976 31116 41024 31132
rect 42044 31132 42048 31330
rect 43080 31424 43148 31602
rect 43080 31336 43106 31424
rect 42082 31132 42090 31330
rect 40976 30346 41022 31116
rect 40976 30330 41024 30346
rect 40976 30038 40990 30330
rect 40976 30022 41024 30038
rect 42044 30330 42090 31132
rect 42044 30038 42048 30330
rect 42082 30038 42090 30330
rect 39782 28944 39790 29236
rect 39824 28944 39828 29236
rect 39782 28142 39828 28944
rect 40336 29890 40486 30016
rect 40336 28694 40358 29890
rect 40452 28694 40486 29890
rect 40336 28370 40486 28694
rect 40976 29252 41022 30022
rect 40976 29236 41024 29252
rect 40976 28944 40990 29236
rect 40976 28928 41024 28944
rect 42044 29236 42090 30038
rect 42044 28944 42048 29236
rect 42082 28944 42090 29236
rect 39782 27850 39790 28142
rect 39824 27850 39828 28142
rect 39782 27048 39828 27850
rect 39782 26990 39790 27048
rect 38732 26740 38766 26756
rect 39766 26756 39790 26850
rect 39824 26990 39828 27048
rect 40976 28158 41022 28928
rect 40976 28142 41024 28158
rect 40976 27850 40990 28142
rect 40976 27834 41024 27850
rect 42044 28142 42090 28944
rect 42044 27850 42048 28142
rect 42082 27850 42090 28142
rect 40976 27064 41022 27834
rect 40976 27048 41024 27064
rect 40976 26990 40990 27048
rect 39824 26756 39848 26850
rect 39766 26754 39848 26756
rect 40962 26756 40990 26836
rect 42044 27048 42090 27850
rect 42044 26968 42048 27048
rect 41024 26756 41088 26836
rect 39754 26646 39880 26754
rect 35538 26556 39988 26646
rect 35550 26550 39988 26556
rect 37664 26528 37746 26550
rect 36590 25866 36658 25882
rect 38714 25866 38782 25898
rect 34450 25856 38782 25866
rect 34348 25812 38782 25856
rect 34348 25776 38790 25812
rect 34348 25766 38638 25776
rect 32256 25290 32262 25490
rect 33258 25440 33280 25582
rect 32216 24488 32262 25290
rect 32216 24196 32222 24488
rect 32256 24196 32262 24488
rect 32216 23394 32262 24196
rect 32216 23102 32222 23394
rect 32256 23102 32262 23394
rect 32216 22300 32262 23102
rect 32216 22008 32222 22300
rect 32256 22008 32262 22300
rect 32216 21206 32262 22008
rect 32216 21176 32222 21206
rect 31198 20914 31236 20986
rect 31154 20804 31236 20914
rect 32256 21176 32262 21206
rect 33272 25290 33280 25440
rect 33314 25440 33384 25582
rect 34450 25588 34576 25766
rect 34450 25552 34500 25588
rect 33314 25290 33318 25440
rect 33272 24488 33318 25290
rect 33272 24196 33280 24488
rect 33314 24196 33318 24488
rect 33272 23394 33318 24196
rect 34486 25296 34500 25552
rect 34534 25552 34576 25588
rect 35558 25588 35592 25604
rect 34534 25486 34554 25552
rect 34486 25280 34534 25296
rect 35554 25296 35558 25494
rect 36590 25588 36658 25766
rect 36590 25500 36616 25588
rect 35592 25296 35600 25494
rect 34486 24510 34532 25280
rect 34486 24494 34534 24510
rect 34486 24202 34500 24494
rect 34486 24186 34534 24202
rect 35554 24494 35600 25296
rect 35554 24202 35558 24494
rect 35592 24202 35600 24494
rect 33272 23102 33280 23394
rect 33314 23102 33318 23394
rect 33272 22300 33318 23102
rect 33846 24054 33996 24180
rect 33846 22858 33868 24054
rect 33962 22858 33996 24054
rect 33846 22534 33996 22858
rect 34486 23416 34532 24186
rect 34486 23400 34534 23416
rect 34486 23108 34500 23400
rect 34486 23092 34534 23108
rect 35554 23400 35600 24202
rect 35554 23108 35558 23400
rect 35592 23108 35600 23400
rect 33272 22008 33280 22300
rect 33314 22008 33318 22300
rect 33272 21206 33318 22008
rect 33272 21148 33280 21206
rect 33256 20958 33280 21008
rect 32222 20898 32256 20914
rect 33244 20914 33280 20958
rect 33314 21148 33318 21206
rect 34486 22322 34532 23092
rect 34486 22306 34534 22322
rect 34486 22014 34500 22306
rect 34486 21998 34534 22014
rect 35554 22306 35600 23108
rect 35554 22014 35558 22306
rect 35592 22014 35600 22306
rect 34486 21228 34532 21998
rect 34486 21212 34534 21228
rect 34486 21170 34500 21212
rect 33314 20958 33338 21008
rect 33314 20914 33370 20958
rect 33244 20804 33370 20914
rect 34466 20920 34500 21170
rect 35554 21212 35600 22014
rect 34534 20920 34592 21170
rect 35554 21132 35558 21212
rect 29028 20714 33478 20804
rect 29040 20708 33478 20714
rect 31154 20686 31236 20708
rect 30080 19996 30148 20012
rect 32204 19996 32272 20028
rect 27926 19986 32272 19996
rect 27838 19942 32272 19986
rect 27838 19906 32280 19942
rect 27838 19896 32128 19906
rect 27926 19850 28058 19896
rect 25734 19410 25740 19610
rect 26688 19596 26758 19702
rect 25694 18608 25740 19410
rect 25694 18316 25700 18608
rect 25734 18316 25740 18608
rect 25694 17514 25740 18316
rect 25694 17222 25700 17514
rect 25734 17222 25740 17514
rect 25694 16420 25740 17222
rect 25694 16128 25700 16420
rect 25734 16128 25740 16420
rect 25694 15326 25740 16128
rect 25694 15296 25700 15326
rect 24676 15034 24714 15106
rect 24632 14924 24714 15034
rect 25734 15296 25740 15326
rect 26750 19410 26758 19596
rect 26792 19596 26820 19702
rect 27976 19718 28044 19850
rect 26792 19410 26796 19596
rect 26750 18608 26796 19410
rect 26750 18316 26758 18608
rect 26792 18316 26796 18608
rect 26750 17514 26796 18316
rect 27976 19426 27990 19718
rect 28024 19616 28044 19718
rect 29048 19718 29082 19734
rect 27976 19410 28024 19426
rect 29044 19426 29048 19624
rect 30080 19718 30148 19896
rect 30080 19630 30106 19718
rect 29082 19426 29090 19624
rect 27976 18640 28022 19410
rect 27976 18624 28024 18640
rect 27976 18332 27990 18624
rect 27976 18316 28024 18332
rect 29044 18624 29090 19426
rect 29044 18332 29048 18624
rect 29082 18332 29090 18624
rect 26750 17222 26758 17514
rect 26792 17222 26796 17514
rect 26750 16420 26796 17222
rect 27336 18184 27486 18310
rect 27336 16988 27358 18184
rect 27452 16988 27486 18184
rect 27336 16664 27486 16988
rect 27976 17546 28022 18316
rect 27976 17530 28024 17546
rect 27976 17238 27990 17530
rect 27976 17222 28024 17238
rect 29044 17530 29090 18332
rect 29044 17238 29048 17530
rect 29082 17238 29090 17530
rect 26750 16128 26758 16420
rect 26792 16128 26796 16420
rect 26750 15326 26796 16128
rect 27976 16452 28022 17222
rect 27976 16436 28024 16452
rect 27976 16144 27990 16436
rect 27976 16128 28024 16144
rect 29044 16436 29090 17238
rect 29044 16144 29048 16436
rect 29082 16144 29090 16436
rect 27976 15376 28022 16128
rect 26750 15268 26758 15326
rect 26748 15128 26758 15160
rect 25700 15018 25734 15034
rect 26734 15034 26758 15128
rect 26792 15268 26796 15326
rect 27970 15342 28102 15376
rect 26792 15034 26880 15160
rect 26734 14924 26880 15034
rect 27970 15050 27990 15342
rect 28024 15050 28102 15342
rect 29044 15342 29090 16144
rect 29044 15262 29048 15342
rect 22506 14834 26956 14924
rect 22518 14828 26956 14834
rect 24632 14806 24714 14828
rect 23568 14124 23636 14140
rect 25692 14124 25760 14156
rect 21440 14114 25760 14124
rect 21326 14070 25760 14114
rect 21326 14034 25768 14070
rect 21326 14024 25616 14034
rect 21440 13922 21572 14024
rect 19254 13570 19260 13770
rect 19214 12768 19260 13570
rect 19214 12476 19220 12768
rect 19254 12476 19260 12768
rect 19214 11674 19260 12476
rect 19214 11382 19220 11674
rect 19254 11382 19260 11674
rect 19214 10580 19260 11382
rect 19214 10288 19220 10580
rect 19254 10288 19260 10580
rect 19214 9486 19260 10288
rect 19214 9456 19220 9486
rect 18196 9194 18234 9266
rect 18152 9084 18234 9194
rect 19254 9456 19260 9486
rect 20242 13570 20278 13862
rect 20312 13570 20336 13862
rect 20242 12768 20336 13570
rect 20242 12476 20278 12768
rect 20312 12476 20336 12768
rect 20242 11674 20336 12476
rect 21464 13846 21532 13922
rect 21464 13554 21478 13846
rect 21512 13744 21532 13846
rect 22536 13846 22570 13862
rect 21464 13538 21512 13554
rect 22532 13554 22536 13752
rect 23568 13846 23636 14024
rect 23568 13758 23594 13846
rect 22570 13554 22578 13752
rect 21464 12768 21510 13538
rect 21464 12752 21512 12768
rect 21464 12460 21478 12752
rect 21464 12444 21512 12460
rect 22532 12752 22578 13554
rect 22532 12460 22536 12752
rect 22570 12460 22578 12752
rect 20242 11382 20278 11674
rect 20312 11382 20336 11674
rect 20242 10580 20336 11382
rect 20824 12312 20974 12438
rect 20824 11116 20846 12312
rect 20940 11116 20974 12312
rect 20824 10792 20974 11116
rect 21464 11674 21510 12444
rect 21464 11658 21512 11674
rect 21464 11366 21478 11658
rect 21464 11350 21512 11366
rect 22532 11658 22578 12460
rect 22532 11366 22536 11658
rect 22570 11366 22578 11658
rect 20242 10288 20278 10580
rect 20312 10288 20336 10580
rect 20242 9486 20336 10288
rect 19220 9178 19254 9194
rect 20242 9194 20278 9486
rect 20312 9226 20336 9486
rect 21464 10580 21510 11350
rect 21464 10564 21512 10580
rect 21464 10272 21478 10564
rect 21464 10256 21512 10272
rect 22532 10564 22578 11366
rect 22532 10272 22536 10564
rect 22570 10272 22578 10564
rect 21464 9486 21510 10256
rect 21464 9470 21512 9486
rect 21464 9416 21478 9470
rect 20312 9194 20380 9226
rect 20242 9084 20380 9194
rect 21454 9178 21478 9416
rect 22532 9470 22578 10272
rect 21512 9382 21524 9416
rect 22532 9390 22536 9470
rect 21512 9178 21586 9382
rect 16026 8994 20476 9084
rect 16038 8988 20476 8994
rect 18152 8966 18234 8988
rect 17096 8232 17164 8248
rect 19220 8232 19288 8264
rect 14940 8222 19288 8232
rect 14854 8178 19288 8222
rect 14854 8142 19296 8178
rect 14854 8132 19144 8142
rect 12766 7654 12772 7854
rect 13768 7840 13790 7946
rect 12726 6852 12772 7654
rect 12726 6560 12732 6852
rect 12766 6560 12772 6852
rect 12726 5758 12772 6560
rect 12726 5466 12732 5758
rect 12766 5466 12772 5758
rect 12726 4664 12772 5466
rect 12726 4372 12732 4664
rect 12766 4372 12772 4664
rect 12726 3570 12772 4372
rect 12726 3540 12732 3570
rect 11708 3278 11746 3350
rect 11664 3168 11746 3278
rect 12766 3540 12772 3570
rect 13782 7654 13790 7840
rect 13824 7840 13874 7946
rect 14940 7954 15072 8132
rect 13824 7654 13828 7840
rect 14940 7832 15006 7954
rect 13782 6852 13828 7654
rect 13782 6560 13790 6852
rect 13824 6560 13828 6852
rect 13782 5758 13828 6560
rect 14992 7662 15006 7832
rect 15040 7832 15072 7954
rect 16064 7954 16098 7970
rect 14992 7646 15040 7662
rect 16060 7662 16064 7860
rect 17096 7954 17164 8132
rect 17096 7866 17122 7954
rect 16098 7662 16106 7860
rect 14992 6876 15038 7646
rect 14992 6860 15040 6876
rect 14992 6568 15006 6860
rect 14992 6552 15040 6568
rect 16060 6860 16106 7662
rect 16060 6568 16064 6860
rect 16098 6568 16106 6860
rect 13782 5466 13790 5758
rect 13824 5466 13828 5758
rect 13782 4664 13828 5466
rect 14352 6420 14502 6546
rect 14352 5224 14374 6420
rect 14468 5224 14502 6420
rect 14352 4900 14502 5224
rect 14992 5782 15038 6552
rect 14992 5766 15040 5782
rect 14992 5474 15006 5766
rect 14992 5458 15040 5474
rect 16060 5766 16106 6568
rect 16060 5474 16064 5766
rect 16098 5474 16106 5766
rect 13782 4372 13790 4664
rect 13824 4372 13828 4664
rect 13782 3570 13828 4372
rect 13782 3512 13790 3570
rect 12732 3262 12766 3278
rect 13766 3278 13790 3372
rect 13824 3512 13828 3570
rect 14992 4688 15038 5458
rect 14992 4672 15040 4688
rect 14992 4380 15006 4672
rect 14992 4364 15040 4380
rect 16060 4672 16106 5474
rect 16060 4380 16064 4672
rect 16098 4380 16106 4672
rect 14992 3594 15038 4364
rect 14992 3578 15040 3594
rect 14992 3520 15006 3578
rect 13824 3278 13848 3372
rect 13766 3168 13848 3278
rect 16060 3578 16106 4380
rect 16060 3498 16064 3578
rect 15006 3270 15040 3286
rect 16044 3286 16064 3386
rect 16098 3498 16106 3578
rect 17112 7662 17122 7866
rect 17156 7918 17164 7954
rect 18180 7954 18214 7970
rect 17156 7866 17170 7918
rect 17156 7662 17158 7866
rect 17112 6860 17158 7662
rect 17112 6568 17122 6860
rect 17156 6568 17158 6860
rect 17112 5766 17158 6568
rect 17112 5474 17122 5766
rect 17156 5474 17158 5766
rect 17112 4672 17158 5474
rect 17112 4380 17122 4672
rect 17156 4380 17158 4672
rect 17112 3578 17158 4380
rect 17112 3520 17122 3578
rect 16098 3286 16126 3386
rect 16044 3176 16126 3286
rect 17156 3520 17158 3578
rect 19212 7954 19296 8142
rect 18214 7662 18226 7866
rect 19212 7862 19238 7954
rect 18180 6860 18226 7662
rect 18214 6568 18226 6860
rect 18180 5766 18226 6568
rect 18214 5474 18226 5766
rect 18180 4672 18226 5474
rect 18214 4380 18226 4672
rect 18180 3578 18226 4380
rect 17122 3270 17156 3286
rect 18170 3286 18180 3358
rect 18214 3504 18226 3578
rect 19232 7662 19238 7862
rect 19272 7862 19296 7954
rect 20242 7954 20380 8988
rect 21454 8216 21586 9178
rect 22516 9178 22536 9278
rect 22570 9390 22578 9470
rect 23584 13554 23594 13758
rect 23628 13810 23636 13846
rect 24652 13846 24686 13862
rect 23628 13758 23642 13810
rect 23628 13554 23630 13758
rect 23584 12752 23630 13554
rect 23584 12460 23594 12752
rect 23628 12460 23630 12752
rect 23584 11658 23630 12460
rect 23584 11366 23594 11658
rect 23628 11366 23630 11658
rect 23584 10564 23630 11366
rect 23584 10272 23594 10564
rect 23628 10272 23630 10564
rect 23584 9470 23630 10272
rect 23584 9412 23594 9470
rect 22570 9178 22598 9278
rect 22516 9068 22598 9178
rect 23628 9412 23630 9470
rect 25684 13846 25768 14034
rect 24686 13554 24698 13758
rect 25684 13754 25710 13846
rect 24652 12752 24698 13554
rect 24686 12460 24698 12752
rect 24652 11658 24698 12460
rect 24686 11366 24698 11658
rect 24652 10564 24698 11366
rect 24686 10272 24698 10564
rect 24652 9470 24698 10272
rect 23594 9162 23628 9178
rect 24642 9178 24652 9250
rect 24686 9396 24698 9470
rect 25704 13554 25710 13754
rect 25744 13754 25768 13846
rect 26748 13846 26880 14828
rect 27970 14140 28102 15050
rect 29028 15050 29048 15150
rect 29082 15262 29090 15342
rect 30096 19426 30106 19630
rect 30140 19682 30148 19718
rect 31164 19718 31198 19734
rect 30140 19630 30154 19682
rect 30140 19426 30142 19630
rect 30096 18624 30142 19426
rect 30096 18332 30106 18624
rect 30140 18332 30142 18624
rect 30096 17530 30142 18332
rect 30096 17238 30106 17530
rect 30140 17238 30142 17530
rect 30096 16436 30142 17238
rect 30096 16144 30106 16436
rect 30140 16144 30142 16436
rect 30096 15342 30142 16144
rect 30096 15284 30106 15342
rect 29082 15050 29110 15150
rect 29028 14940 29110 15050
rect 30140 15284 30142 15342
rect 32196 19718 32280 19906
rect 31198 19426 31210 19630
rect 32196 19626 32222 19718
rect 31164 18624 31210 19426
rect 31198 18332 31210 18624
rect 31164 17530 31210 18332
rect 31198 17238 31210 17530
rect 31164 16436 31210 17238
rect 31198 16144 31210 16436
rect 31164 15342 31210 16144
rect 30106 15034 30140 15050
rect 31154 15050 31164 15122
rect 31198 15268 31210 15342
rect 32216 19426 32222 19626
rect 32256 19626 32280 19718
rect 33244 19718 33370 20708
rect 34466 20002 34592 20920
rect 35538 20920 35558 21020
rect 35592 21132 35600 21212
rect 36606 25296 36616 25500
rect 36650 25552 36658 25588
rect 37674 25588 37708 25604
rect 36650 25500 36664 25552
rect 36650 25296 36652 25500
rect 36606 24494 36652 25296
rect 36606 24202 36616 24494
rect 36650 24202 36652 24494
rect 36606 23400 36652 24202
rect 36606 23108 36616 23400
rect 36650 23108 36652 23400
rect 36606 22306 36652 23108
rect 36606 22014 36616 22306
rect 36650 22014 36652 22306
rect 36606 21212 36652 22014
rect 36606 21154 36616 21212
rect 35592 20920 35620 21020
rect 35538 20810 35620 20920
rect 36650 21154 36652 21212
rect 38706 25588 38790 25776
rect 37708 25296 37720 25500
rect 38706 25496 38732 25588
rect 37674 24494 37720 25296
rect 37708 24202 37720 24494
rect 37674 23400 37720 24202
rect 37708 23108 37720 23400
rect 37674 22306 37720 23108
rect 37708 22014 37720 22306
rect 37674 21212 37720 22014
rect 36616 20904 36650 20920
rect 37664 20920 37674 20992
rect 37708 21138 37720 21212
rect 38726 25296 38732 25496
rect 38766 25496 38790 25588
rect 39754 25588 39880 26550
rect 40962 25866 41088 26756
rect 42028 26756 42048 26856
rect 42082 26968 42090 27048
rect 43096 31132 43106 31336
rect 43140 31388 43148 31424
rect 44164 31424 44198 31440
rect 43140 31336 43154 31388
rect 43140 31132 43142 31336
rect 43096 30330 43142 31132
rect 43096 30038 43106 30330
rect 43140 30038 43142 30330
rect 43096 29236 43142 30038
rect 43096 28944 43106 29236
rect 43140 28944 43142 29236
rect 43096 28142 43142 28944
rect 43096 27850 43106 28142
rect 43140 27850 43142 28142
rect 43096 27048 43142 27850
rect 43096 26990 43106 27048
rect 42082 26756 42110 26856
rect 42028 26646 42110 26756
rect 43140 26990 43142 27048
rect 45196 31424 45280 31612
rect 44198 31132 44210 31336
rect 45196 31332 45222 31424
rect 44164 30330 44210 31132
rect 44198 30038 44210 30330
rect 44164 29236 44210 30038
rect 44198 28944 44210 29236
rect 44164 28142 44210 28944
rect 44198 27850 44210 28142
rect 44164 27048 44210 27850
rect 43106 26740 43140 26756
rect 44154 26756 44164 26828
rect 44198 26974 44210 27048
rect 45216 31132 45222 31332
rect 45256 31332 45280 31424
rect 46242 31424 46368 32384
rect 47524 31724 47656 32612
rect 48616 32612 48636 32712
rect 48670 32824 48678 32904
rect 49684 36988 49694 37192
rect 49728 37244 49736 37280
rect 50752 37280 50786 37296
rect 49728 37192 49742 37244
rect 49728 36988 49730 37192
rect 49684 36186 49730 36988
rect 49684 35894 49694 36186
rect 49728 35894 49730 36186
rect 49684 35092 49730 35894
rect 49684 34800 49694 35092
rect 49728 34800 49730 35092
rect 49684 33998 49730 34800
rect 49684 33706 49694 33998
rect 49728 33706 49730 33998
rect 49684 32904 49730 33706
rect 49684 32846 49694 32904
rect 48670 32612 48698 32712
rect 48616 32502 48698 32612
rect 49728 32846 49730 32904
rect 51784 37280 51868 37468
rect 50786 36988 50798 37192
rect 51784 37188 51810 37280
rect 50752 36186 50798 36988
rect 50786 35894 50798 36186
rect 50752 35092 50798 35894
rect 50786 34800 50798 35092
rect 50752 33998 50798 34800
rect 50786 33706 50798 33998
rect 50752 32904 50798 33706
rect 49694 32596 49728 32612
rect 50742 32612 50752 32684
rect 50786 32830 50798 32904
rect 51804 36988 51810 37188
rect 51844 37188 51868 37280
rect 52850 37280 52946 38222
rect 54062 37572 54158 38442
rect 55130 38442 55150 38542
rect 55184 38654 55192 38734
rect 56198 42818 56208 43022
rect 56242 43074 56250 43110
rect 57266 43110 57300 43126
rect 56242 43022 56256 43074
rect 56242 42818 56244 43022
rect 56198 42016 56244 42818
rect 56198 41724 56208 42016
rect 56242 41724 56244 42016
rect 56198 40922 56244 41724
rect 56198 40630 56208 40922
rect 56242 40630 56244 40922
rect 56198 39828 56244 40630
rect 56198 39536 56208 39828
rect 56242 39536 56244 39828
rect 56198 38734 56244 39536
rect 56198 38676 56208 38734
rect 55184 38442 55212 38542
rect 55130 38332 55212 38442
rect 56242 38676 56244 38734
rect 58298 43110 58382 43198
rect 57300 42818 57312 43022
rect 58298 43018 58324 43110
rect 57266 42016 57312 42818
rect 57300 41724 57312 42016
rect 57266 40922 57312 41724
rect 57300 40630 57312 40922
rect 57266 39828 57312 40630
rect 57300 39536 57312 39828
rect 57266 38734 57312 39536
rect 56208 38426 56242 38442
rect 57256 38442 57266 38514
rect 57300 38660 57312 38734
rect 58318 42818 58324 43018
rect 58358 43018 58382 43110
rect 59348 43110 59446 43198
rect 58358 42818 58364 43018
rect 59348 42864 59382 43110
rect 58318 42016 58364 42818
rect 58318 41724 58324 42016
rect 58358 41724 58364 42016
rect 58318 40922 58364 41724
rect 58318 40630 58324 40922
rect 58358 40630 58364 40922
rect 58318 39828 58364 40630
rect 58318 39536 58324 39828
rect 58358 39536 58364 39828
rect 58318 38734 58364 39536
rect 58318 38704 58324 38734
rect 57300 38442 57338 38514
rect 57256 38332 57338 38442
rect 58358 38704 58364 38734
rect 59374 42818 59382 42864
rect 59416 42864 59446 43110
rect 62478 43268 62560 43284
rect 63842 43276 63992 43444
rect 66242 43426 66448 43532
rect 65776 43282 65850 43286
rect 63816 43272 63992 43276
rect 63808 43268 63992 43272
rect 65066 43268 65860 43282
rect 62478 43192 65860 43268
rect 62478 43108 62560 43192
rect 62478 42964 62508 43108
rect 62498 42936 62508 42964
rect 62542 42964 62560 43108
rect 63166 43108 63200 43124
rect 62542 42936 62556 42964
rect 59416 42818 59420 42864
rect 59374 42016 59420 42818
rect 59374 41724 59382 42016
rect 59416 41724 59420 42016
rect 62148 42630 62360 42700
rect 59374 40922 59420 41724
rect 59374 40630 59382 40922
rect 59416 40630 59420 40922
rect 59374 39828 59420 40630
rect 59530 41772 59934 41952
rect 59530 40204 59572 41772
rect 59836 40204 59934 41772
rect 62148 40876 62180 42630
rect 62328 40876 62360 42630
rect 62148 40790 62360 40876
rect 62498 42414 62556 42936
rect 62498 42242 62508 42414
rect 62542 42242 62556 42414
rect 62498 41720 62556 42242
rect 62498 41548 62508 41720
rect 62542 41548 62556 41720
rect 62498 41026 62556 41548
rect 62498 40854 62508 41026
rect 62542 40854 62556 41026
rect 62498 40332 62556 40854
rect 62498 40266 62508 40332
rect 59530 40066 59934 40204
rect 62542 40266 62556 40332
rect 63156 42936 63166 43036
rect 63808 43108 63878 43192
rect 65066 43164 65860 43192
rect 66268 43270 66448 43426
rect 67732 43438 67818 43584
rect 68110 43438 68228 43584
rect 67732 43396 68228 43438
rect 67610 43274 67672 43278
rect 67602 43270 67672 43274
rect 68904 43270 68998 43274
rect 66268 43194 68998 43270
rect 63200 42936 63214 43036
rect 63156 42414 63214 42936
rect 63156 42242 63166 42414
rect 63200 42242 63214 42414
rect 63156 41720 63214 42242
rect 63156 41548 63166 41720
rect 63200 41548 63214 41720
rect 63156 41026 63214 41548
rect 63156 40854 63166 41026
rect 63200 40854 63214 41026
rect 63156 40332 63214 40854
rect 63156 40270 63166 40332
rect 62508 40144 62542 40160
rect 63158 40160 63166 40270
rect 63200 40270 63214 40332
rect 63808 42936 63824 43108
rect 63858 42952 63878 43108
rect 64482 43108 64516 43124
rect 63858 42936 63866 42952
rect 63808 42414 63866 42936
rect 63808 42242 63824 42414
rect 63858 42242 63866 42414
rect 63808 41720 63866 42242
rect 63808 41548 63824 41720
rect 63858 41548 63866 41720
rect 63808 41026 63866 41548
rect 63808 40854 63824 41026
rect 63858 40854 63866 41026
rect 63808 40332 63866 40854
rect 63808 40270 63824 40332
rect 63200 40160 63212 40270
rect 63158 40072 63212 40160
rect 63858 40270 63866 40332
rect 64470 42936 64482 43072
rect 65110 43108 65204 43164
rect 64516 42936 64528 43072
rect 64470 42414 64528 42936
rect 65110 42936 65140 43108
rect 65174 42936 65204 43108
rect 65776 43108 65850 43164
rect 66268 43146 66448 43194
rect 65776 43054 65798 43108
rect 65774 43008 65798 43054
rect 65110 42890 65204 42936
rect 65788 42936 65798 43008
rect 65832 43054 65850 43108
rect 66272 43110 66354 43146
rect 65832 43008 65854 43054
rect 65832 42936 65846 43008
rect 66272 42966 66302 43110
rect 64470 42242 64482 42414
rect 64516 42242 64528 42414
rect 64470 41720 64528 42242
rect 64470 41548 64482 41720
rect 64516 41548 64528 41720
rect 64470 41026 64528 41548
rect 64470 40854 64482 41026
rect 64516 40854 64528 41026
rect 64470 40332 64528 40854
rect 64470 40306 64482 40332
rect 63824 40144 63858 40160
rect 64476 40160 64482 40268
rect 64516 40306 64528 40332
rect 65124 42414 65182 42890
rect 65124 42242 65140 42414
rect 65174 42242 65182 42414
rect 65124 41720 65182 42242
rect 65124 41548 65140 41720
rect 65174 41548 65182 41720
rect 65124 41026 65182 41548
rect 65124 40854 65140 41026
rect 65174 40854 65182 41026
rect 65124 40332 65182 40854
rect 65124 40274 65140 40332
rect 64516 40160 64530 40268
rect 64476 40072 64530 40160
rect 65174 40274 65182 40332
rect 65788 42664 65846 42936
rect 66292 42938 66302 42966
rect 66336 42966 66354 43110
rect 66960 43110 66994 43126
rect 66336 42938 66350 42966
rect 65886 42664 66202 42918
rect 65788 42632 66202 42664
rect 65788 42544 65974 42632
rect 65788 42414 65846 42544
rect 65886 42448 65974 42544
rect 65788 42242 65798 42414
rect 65832 42242 65846 42414
rect 65788 41720 65846 42242
rect 65788 41548 65798 41720
rect 65832 41548 65846 41720
rect 65788 41026 65846 41548
rect 65788 40854 65798 41026
rect 65832 40854 65846 41026
rect 65788 40332 65846 40854
rect 65942 40878 65974 42448
rect 66122 42448 66202 42632
rect 66122 40878 66154 42448
rect 65942 40792 66154 40878
rect 66292 42416 66350 42938
rect 66292 42244 66302 42416
rect 66336 42244 66350 42416
rect 66292 41722 66350 42244
rect 66292 41550 66302 41722
rect 66336 41550 66350 41722
rect 66292 41028 66350 41550
rect 66292 40856 66302 41028
rect 66336 40856 66350 41028
rect 65788 40272 65798 40332
rect 65140 40144 65174 40160
rect 65784 40160 65798 40272
rect 65832 40248 65846 40332
rect 66292 40334 66350 40856
rect 66292 40268 66302 40334
rect 65832 40160 65838 40248
rect 65784 40072 65838 40160
rect 66336 40268 66350 40334
rect 66950 42938 66960 43038
rect 67602 43110 67672 43194
rect 66994 42938 67008 43038
rect 66950 42416 67008 42938
rect 66950 42244 66960 42416
rect 66994 42244 67008 42416
rect 66950 41722 67008 42244
rect 66950 41550 66960 41722
rect 66994 41550 67008 41722
rect 66950 41028 67008 41550
rect 66950 40856 66960 41028
rect 66994 40856 67008 41028
rect 66950 40334 67008 40856
rect 66950 40272 66960 40334
rect 66302 40146 66336 40162
rect 66952 40162 66960 40272
rect 66994 40272 67008 40334
rect 67602 42938 67618 43110
rect 67652 42954 67672 43110
rect 68276 43110 68310 43126
rect 67652 42938 67660 42954
rect 67602 42416 67660 42938
rect 67602 42244 67618 42416
rect 67652 42244 67660 42416
rect 67602 41722 67660 42244
rect 67602 41550 67618 41722
rect 67652 41550 67660 41722
rect 67602 41028 67660 41550
rect 67602 40856 67618 41028
rect 67652 40856 67660 41028
rect 67602 40334 67660 40856
rect 67602 40272 67618 40334
rect 66994 40162 67006 40272
rect 66952 40074 67006 40162
rect 67652 40272 67660 40334
rect 68264 42938 68276 43074
rect 68904 43110 68998 43194
rect 68310 42938 68322 43074
rect 68264 42416 68322 42938
rect 68904 42938 68934 43110
rect 68968 42938 68998 43110
rect 68904 42892 68998 42938
rect 69578 43110 69748 43548
rect 71570 43444 71596 43614
rect 71844 43444 71878 43614
rect 71570 43426 71878 43444
rect 70100 43300 70162 43310
rect 69578 42938 69592 43110
rect 69626 42938 69748 43110
rect 70080 43284 70162 43300
rect 71418 43288 71480 43292
rect 71410 43284 71480 43288
rect 71656 43284 71788 43426
rect 72712 43286 72806 43288
rect 73364 43286 73456 43288
rect 72712 43284 73460 43286
rect 70080 43208 73460 43284
rect 70080 43124 70162 43208
rect 70080 42980 70110 43124
rect 69578 42916 69748 42938
rect 70100 42952 70110 42980
rect 70144 42980 70162 43124
rect 70768 43124 70802 43140
rect 70144 42952 70158 42980
rect 68264 42244 68276 42416
rect 68310 42244 68322 42416
rect 68264 41722 68322 42244
rect 68264 41550 68276 41722
rect 68310 41550 68322 41722
rect 68264 41028 68322 41550
rect 68264 40856 68276 41028
rect 68310 40856 68322 41028
rect 68264 40334 68322 40856
rect 68264 40308 68276 40334
rect 67618 40146 67652 40162
rect 68270 40162 68276 40270
rect 68310 40308 68322 40334
rect 68918 42416 68976 42892
rect 68918 42244 68934 42416
rect 68968 42244 68976 42416
rect 68918 41722 68976 42244
rect 69582 42416 69640 42916
rect 69582 42244 69592 42416
rect 69626 42244 69640 42416
rect 69582 41896 69640 42244
rect 69750 42646 69962 42716
rect 69750 41896 69782 42646
rect 69568 41790 69782 41896
rect 68918 41550 68934 41722
rect 68968 41550 68976 41722
rect 68918 41028 68976 41550
rect 68918 40856 68934 41028
rect 68968 40856 68976 41028
rect 68918 40334 68976 40856
rect 68918 40276 68934 40334
rect 68310 40162 68324 40270
rect 68270 40074 68324 40162
rect 68968 40276 68976 40334
rect 69582 41722 69640 41790
rect 69582 41550 69592 41722
rect 69626 41550 69640 41722
rect 69582 41028 69640 41550
rect 69582 40856 69592 41028
rect 69626 40856 69640 41028
rect 69582 40334 69640 40856
rect 69750 40892 69782 41790
rect 69930 40892 69962 42646
rect 69750 40806 69962 40892
rect 70100 42430 70158 42952
rect 70100 42258 70110 42430
rect 70144 42258 70158 42430
rect 70100 41736 70158 42258
rect 70100 41564 70110 41736
rect 70144 41564 70158 41736
rect 70100 41042 70158 41564
rect 70100 40870 70110 41042
rect 70144 40870 70158 41042
rect 69582 40274 69592 40334
rect 68934 40146 68968 40162
rect 69578 40162 69592 40274
rect 69626 40250 69640 40334
rect 70100 40348 70158 40870
rect 70100 40282 70110 40348
rect 69626 40162 69632 40250
rect 69578 40074 69632 40162
rect 70144 40282 70158 40348
rect 70758 42952 70768 43052
rect 71410 43124 71480 43208
rect 71656 43202 71788 43208
rect 72712 43192 73460 43208
rect 70802 42952 70816 43052
rect 70758 42430 70816 42952
rect 70758 42258 70768 42430
rect 70802 42258 70816 42430
rect 70758 41736 70816 42258
rect 70758 41564 70768 41736
rect 70802 41564 70816 41736
rect 70758 41042 70816 41564
rect 70758 40870 70768 41042
rect 70802 40870 70816 41042
rect 70758 40348 70816 40870
rect 70758 40286 70768 40348
rect 70110 40160 70144 40176
rect 70760 40176 70768 40286
rect 70802 40286 70816 40348
rect 71410 42952 71426 43124
rect 71460 42968 71480 43124
rect 72084 43124 72118 43140
rect 71460 42952 71468 42968
rect 71410 42430 71468 42952
rect 71410 42258 71426 42430
rect 71460 42258 71468 42430
rect 71410 41736 71468 42258
rect 71410 41564 71426 41736
rect 71460 41564 71468 41736
rect 71410 41042 71468 41564
rect 71410 40870 71426 41042
rect 71460 40870 71468 41042
rect 71410 40348 71468 40870
rect 71410 40286 71426 40348
rect 70802 40176 70814 40286
rect 70760 40088 70814 40176
rect 71460 40286 71468 40348
rect 72072 42952 72084 43088
rect 72712 43124 72806 43192
rect 72118 42952 72130 43088
rect 72072 42430 72130 42952
rect 72712 42952 72742 43124
rect 72776 42952 72806 43124
rect 73364 43124 73456 43192
rect 73364 43034 73400 43124
rect 72712 42906 72806 42952
rect 73374 42952 73400 43034
rect 73434 43080 73456 43124
rect 73434 42952 73460 43080
rect 73374 42942 73460 42952
rect 72072 42258 72084 42430
rect 72118 42258 72130 42430
rect 72072 41736 72130 42258
rect 72072 41564 72084 41736
rect 72118 41564 72130 41736
rect 72072 41042 72130 41564
rect 72072 40870 72084 41042
rect 72118 40870 72130 41042
rect 72072 40348 72130 40870
rect 72072 40322 72084 40348
rect 71426 40160 71460 40176
rect 72078 40176 72084 40284
rect 72118 40322 72130 40348
rect 72726 42430 72784 42906
rect 72726 42258 72742 42430
rect 72776 42258 72784 42430
rect 72726 41736 72784 42258
rect 72726 41564 72742 41736
rect 72776 41564 72784 41736
rect 72726 41042 72784 41564
rect 72726 40870 72742 41042
rect 72776 40870 72784 41042
rect 72726 40348 72784 40870
rect 72726 40290 72742 40348
rect 72118 40176 72132 40284
rect 72078 40088 72132 40176
rect 72776 40290 72784 40348
rect 73390 42896 73448 42942
rect 73610 42896 73950 43002
rect 73390 42876 73950 42896
rect 73390 42786 73646 42876
rect 73390 42430 73448 42786
rect 73390 42258 73400 42430
rect 73434 42258 73448 42430
rect 73390 41736 73448 42258
rect 73390 41564 73400 41736
rect 73434 41564 73448 41736
rect 73390 41042 73448 41564
rect 73390 40870 73400 41042
rect 73434 40870 73448 41042
rect 73390 40348 73448 40870
rect 73610 40970 73646 42786
rect 73876 40970 73950 42876
rect 73610 40668 73950 40970
rect 73390 40288 73400 40348
rect 72742 40160 72776 40176
rect 73386 40176 73400 40288
rect 73434 40264 73448 40348
rect 73434 40176 73440 40264
rect 73386 40088 73440 40176
rect 63142 39974 65846 40072
rect 66936 39976 69640 40074
rect 70744 39990 73448 40088
rect 72078 39986 72132 39990
rect 64476 39970 64530 39974
rect 68270 39972 68324 39976
rect 59374 39536 59382 39828
rect 59416 39536 59420 39828
rect 59374 38734 59420 39536
rect 80846 39538 81140 39582
rect 78496 39510 78834 39528
rect 78496 39406 78536 39510
rect 78796 39406 78834 39510
rect 77088 39254 77242 39398
rect 78496 39386 78834 39406
rect 80846 39410 80866 39538
rect 81116 39410 81140 39538
rect 78476 39254 78538 39264
rect 78574 39254 78706 39386
rect 79100 39254 79232 39294
rect 79776 39254 79838 39284
rect 77088 39200 79860 39254
rect 80414 39248 80568 39392
rect 80846 39390 81140 39410
rect 85028 39524 85372 39542
rect 85028 39412 85060 39524
rect 85316 39412 85372 39524
rect 85028 39402 85372 39412
rect 81802 39248 81864 39258
rect 83102 39248 83164 39278
rect 83724 39248 83878 39392
rect 85094 39248 85254 39402
rect 86696 39284 87008 39388
rect 85748 39248 85870 39260
rect 86412 39248 86474 39278
rect 77088 39160 77242 39200
rect 77144 39094 77206 39160
rect 59374 38676 59382 38734
rect 59358 38470 59382 38536
rect 58324 38426 58358 38442
rect 59342 38442 59382 38470
rect 59416 38676 59420 38734
rect 76634 38980 76978 39082
rect 77144 39006 77170 39094
rect 59416 38442 59440 38536
rect 59342 38332 59440 38442
rect 55130 38242 59580 38332
rect 55142 38236 59580 38242
rect 57256 38214 57338 38236
rect 56182 37572 56250 37588
rect 58306 37572 58374 37604
rect 54062 37562 58374 37572
rect 53940 37518 58374 37562
rect 53940 37482 58382 37518
rect 53940 37472 58230 37482
rect 52850 37198 52868 37280
rect 51844 36988 51850 37188
rect 51804 36186 51850 36988
rect 51804 35894 51810 36186
rect 51844 35894 51850 36186
rect 51804 35092 51850 35894
rect 51804 34800 51810 35092
rect 51844 34800 51850 35092
rect 51804 33998 51850 34800
rect 51804 33706 51810 33998
rect 51844 33706 51850 33998
rect 51804 32904 51850 33706
rect 51804 32874 51810 32904
rect 50786 32612 50824 32684
rect 50742 32502 50824 32612
rect 51844 32874 51850 32904
rect 52860 36988 52868 37198
rect 52902 37198 52946 37280
rect 54062 37294 54158 37472
rect 54062 37264 54092 37294
rect 52902 36988 52906 37198
rect 52860 36186 52906 36988
rect 52860 35894 52868 36186
rect 52902 35894 52906 36186
rect 52860 35092 52906 35894
rect 54078 37002 54092 37264
rect 54126 37264 54158 37294
rect 55150 37294 55184 37310
rect 54126 37192 54146 37264
rect 54078 36986 54126 37002
rect 55146 37002 55150 37200
rect 56182 37294 56250 37472
rect 56182 37206 56208 37294
rect 55184 37002 55192 37200
rect 54078 36216 54124 36986
rect 54078 36200 54126 36216
rect 54078 35908 54092 36200
rect 54078 35892 54126 35908
rect 55146 36200 55192 37002
rect 55146 35908 55150 36200
rect 55184 35908 55192 36200
rect 52860 34800 52868 35092
rect 52902 34800 52906 35092
rect 52860 33998 52906 34800
rect 53438 35760 53588 35886
rect 53438 34564 53460 35760
rect 53554 34564 53588 35760
rect 53438 34240 53588 34564
rect 54078 35122 54124 35892
rect 54078 35106 54126 35122
rect 54078 34814 54092 35106
rect 54078 34798 54126 34814
rect 55146 35106 55192 35908
rect 55146 34814 55150 35106
rect 55184 34814 55192 35106
rect 52860 33706 52868 33998
rect 52902 33706 52906 33998
rect 52860 32904 52906 33706
rect 52860 32846 52868 32904
rect 52844 32702 52868 32706
rect 51810 32596 51844 32612
rect 52842 32612 52868 32702
rect 52902 32846 52906 32904
rect 54078 34028 54124 34798
rect 54078 34012 54126 34028
rect 54078 33720 54092 34012
rect 54078 33704 54126 33720
rect 55146 34012 55192 34814
rect 55146 33720 55150 34012
rect 55184 33720 55192 34012
rect 54078 32934 54124 33704
rect 54078 32918 54126 32934
rect 54078 32860 54092 32918
rect 52902 32702 52926 32706
rect 52902 32612 52938 32702
rect 52842 32502 52938 32612
rect 54012 32626 54092 32806
rect 55146 32918 55192 33720
rect 55146 32838 55150 32918
rect 54126 32658 54144 32806
rect 54126 32626 54174 32658
rect 48616 32412 53066 32502
rect 48628 32406 53066 32412
rect 50742 32384 50824 32406
rect 49668 31724 49736 31740
rect 51792 31724 51860 31756
rect 47524 31714 51860 31724
rect 47426 31670 51860 31714
rect 47426 31634 51868 31670
rect 47426 31624 51716 31634
rect 45256 31132 45262 31332
rect 46242 31248 46280 31424
rect 45216 30330 45262 31132
rect 45216 30038 45222 30330
rect 45256 30038 45262 30330
rect 45216 29236 45262 30038
rect 45216 28944 45222 29236
rect 45256 28944 45262 29236
rect 45216 28142 45262 28944
rect 45216 27850 45222 28142
rect 45256 27850 45262 28142
rect 45216 27048 45262 27850
rect 45216 27018 45222 27048
rect 44198 26756 44236 26828
rect 44154 26646 44236 26756
rect 45256 27018 45262 27048
rect 46272 31132 46280 31248
rect 46314 31248 46368 31424
rect 47524 31446 47656 31624
rect 47524 31382 47578 31446
rect 46314 31132 46318 31248
rect 46272 30330 46318 31132
rect 46272 30038 46280 30330
rect 46314 30038 46318 30330
rect 47564 31154 47578 31382
rect 47612 31382 47656 31446
rect 48636 31446 48670 31462
rect 47612 31344 47632 31382
rect 47564 31138 47612 31154
rect 48632 31154 48636 31352
rect 49668 31446 49736 31624
rect 49668 31358 49694 31446
rect 48670 31154 48678 31352
rect 47564 30368 47610 31138
rect 47564 30352 47612 30368
rect 47564 30060 47578 30352
rect 47564 30044 47612 30060
rect 48632 30352 48678 31154
rect 48632 30060 48636 30352
rect 48670 30060 48678 30352
rect 46272 29236 46318 30038
rect 46272 28944 46280 29236
rect 46314 28944 46318 29236
rect 46272 28142 46318 28944
rect 46924 29912 47074 30038
rect 46924 28716 46946 29912
rect 47040 28716 47074 29912
rect 46924 28392 47074 28716
rect 47564 29274 47610 30044
rect 47564 29258 47612 29274
rect 47564 28966 47578 29258
rect 47564 28950 47612 28966
rect 48632 29258 48678 30060
rect 48632 28966 48636 29258
rect 48670 28966 48678 29258
rect 46272 27850 46280 28142
rect 46314 27850 46318 28142
rect 46272 27048 46318 27850
rect 47564 28180 47610 28950
rect 47564 28164 47612 28180
rect 47564 27872 47578 28164
rect 47564 27856 47612 27872
rect 48632 28164 48678 28966
rect 48632 27872 48636 28164
rect 48670 27872 48678 28164
rect 47564 27094 47610 27856
rect 46272 26990 46280 27048
rect 45222 26740 45256 26756
rect 46242 26756 46280 26864
rect 46314 26990 46318 27048
rect 47540 27070 47672 27094
rect 46314 26756 46368 26864
rect 46242 26646 46368 26756
rect 47540 26778 47578 27070
rect 47612 26778 47672 27070
rect 48632 27070 48678 27872
rect 48632 26990 48636 27070
rect 42028 26556 46478 26646
rect 42040 26550 46478 26556
rect 44154 26528 44236 26550
rect 43080 25866 43148 25882
rect 45204 25866 45272 25898
rect 40962 25856 45272 25866
rect 40838 25812 45272 25856
rect 40838 25776 45280 25812
rect 40838 25766 45128 25776
rect 38766 25296 38772 25496
rect 39754 25370 39790 25588
rect 38726 24494 38772 25296
rect 38726 24202 38732 24494
rect 38766 24202 38772 24494
rect 38726 23400 38772 24202
rect 38726 23108 38732 23400
rect 38766 23108 38772 23400
rect 38726 22306 38772 23108
rect 38726 22014 38732 22306
rect 38766 22014 38772 22306
rect 38726 21212 38772 22014
rect 38726 21182 38732 21212
rect 37708 20920 37746 20992
rect 37664 20810 37746 20920
rect 38766 21182 38772 21212
rect 39782 25296 39790 25370
rect 39824 25370 39880 25588
rect 40962 25588 41088 25766
rect 40962 25452 40990 25588
rect 39824 25296 39828 25370
rect 39782 24494 39828 25296
rect 39782 24202 39790 24494
rect 39824 24202 39828 24494
rect 39782 23400 39828 24202
rect 40976 25296 40990 25452
rect 41024 25452 41088 25588
rect 42048 25588 42082 25604
rect 40976 25280 41024 25296
rect 42044 25296 42048 25494
rect 43080 25588 43148 25766
rect 43080 25500 43106 25588
rect 42082 25296 42090 25494
rect 40976 24510 41022 25280
rect 40976 24494 41024 24510
rect 40976 24202 40990 24494
rect 40976 24186 41024 24202
rect 42044 24494 42090 25296
rect 42044 24202 42048 24494
rect 42082 24202 42090 24494
rect 39782 23108 39790 23400
rect 39824 23108 39828 23400
rect 39782 22306 39828 23108
rect 40336 24054 40486 24180
rect 40336 22858 40358 24054
rect 40452 22858 40486 24054
rect 40336 22534 40486 22858
rect 40976 23416 41022 24186
rect 40976 23400 41024 23416
rect 40976 23108 40990 23400
rect 40976 23092 41024 23108
rect 42044 23400 42090 24202
rect 42044 23108 42048 23400
rect 42082 23108 42090 23400
rect 39782 22014 39790 22306
rect 39824 22014 39828 22306
rect 39782 21212 39828 22014
rect 39782 21154 39790 21212
rect 39766 20958 39790 21014
rect 38732 20904 38766 20920
rect 39754 20920 39790 20958
rect 39824 21154 39828 21212
rect 40976 22322 41022 23092
rect 40976 22306 41024 22322
rect 40976 22014 40990 22306
rect 40976 21998 41024 22014
rect 42044 22306 42090 23108
rect 42044 22014 42048 22306
rect 42082 22014 42090 22306
rect 40976 21228 41022 21998
rect 40976 21212 41024 21228
rect 40976 21154 40990 21212
rect 39824 20958 39848 21014
rect 39824 20920 39880 20958
rect 39754 20810 39880 20920
rect 40948 20920 40990 21108
rect 42044 21212 42090 22014
rect 42044 21132 42048 21212
rect 41024 20920 41074 21108
rect 35538 20720 39988 20810
rect 35550 20714 39988 20720
rect 37664 20692 37746 20714
rect 36590 20002 36658 20018
rect 38714 20002 38782 20034
rect 34466 19992 38782 20002
rect 34348 19948 38782 19992
rect 34348 19912 38790 19948
rect 34348 19902 38638 19912
rect 34466 19786 34592 19902
rect 32256 19426 32262 19626
rect 33244 19574 33280 19718
rect 32216 18624 32262 19426
rect 32216 18332 32222 18624
rect 32256 18332 32262 18624
rect 32216 17530 32262 18332
rect 32216 17238 32222 17530
rect 32256 17238 32262 17530
rect 32216 16436 32262 17238
rect 32216 16144 32222 16436
rect 32256 16144 32262 16436
rect 32216 15342 32262 16144
rect 32216 15312 32222 15342
rect 31198 15050 31236 15122
rect 31154 14940 31236 15050
rect 32256 15312 32262 15342
rect 33272 19426 33280 19574
rect 33314 19574 33370 19718
rect 34486 19724 34554 19786
rect 33314 19426 33318 19574
rect 33272 18624 33318 19426
rect 33272 18332 33280 18624
rect 33314 18332 33318 18624
rect 33272 17530 33318 18332
rect 34486 19432 34500 19724
rect 34534 19622 34554 19724
rect 35558 19724 35592 19740
rect 34486 19416 34534 19432
rect 35554 19432 35558 19630
rect 36590 19724 36658 19902
rect 36590 19636 36616 19724
rect 35592 19432 35600 19630
rect 34486 18646 34532 19416
rect 34486 18630 34534 18646
rect 34486 18338 34500 18630
rect 34486 18322 34534 18338
rect 35554 18630 35600 19432
rect 35554 18338 35558 18630
rect 35592 18338 35600 18630
rect 33272 17238 33280 17530
rect 33314 17238 33318 17530
rect 33272 16436 33318 17238
rect 33846 18190 33996 18316
rect 33846 16994 33868 18190
rect 33962 16994 33996 18190
rect 33846 16670 33996 16994
rect 34486 17552 34532 18322
rect 34486 17536 34534 17552
rect 34486 17244 34500 17536
rect 34486 17228 34534 17244
rect 35554 17536 35600 18338
rect 35554 17244 35558 17536
rect 35592 17244 35600 17536
rect 33272 16144 33280 16436
rect 33314 16144 33318 16436
rect 33272 15342 33318 16144
rect 33272 15284 33280 15342
rect 32222 15034 32256 15050
rect 33256 15050 33280 15144
rect 33314 15284 33318 15342
rect 34486 16458 34532 17228
rect 34486 16442 34534 16458
rect 34486 16150 34500 16442
rect 34486 16134 34534 16150
rect 35554 16442 35600 17244
rect 35554 16150 35558 16442
rect 35592 16150 35600 16442
rect 34486 15364 34532 16134
rect 34486 15348 34534 15364
rect 34486 15290 34500 15348
rect 33314 15050 33338 15144
rect 33256 15038 33338 15050
rect 34450 15056 34500 15248
rect 35554 15348 35600 16150
rect 35554 15268 35558 15348
rect 34534 15056 34576 15248
rect 33244 14940 33370 15038
rect 29028 14850 33478 14940
rect 29040 14844 33478 14850
rect 31154 14822 31236 14844
rect 30090 14140 30158 14156
rect 32214 14140 32282 14172
rect 27970 14130 32282 14140
rect 27848 14086 32282 14130
rect 27848 14050 32290 14086
rect 27848 14040 32138 14050
rect 27970 13968 28102 14040
rect 25744 13554 25750 13754
rect 26748 13752 26768 13846
rect 25704 12752 25750 13554
rect 25704 12460 25710 12752
rect 25744 12460 25750 12752
rect 25704 11658 25750 12460
rect 25704 11366 25710 11658
rect 25744 11366 25750 11658
rect 25704 10564 25750 11366
rect 25704 10272 25710 10564
rect 25744 10272 25750 10564
rect 25704 9470 25750 10272
rect 25704 9440 25710 9470
rect 24686 9178 24724 9250
rect 24642 9068 24724 9178
rect 25744 9440 25750 9470
rect 26760 13554 26768 13752
rect 26802 13752 26880 13846
rect 27986 13862 28054 13968
rect 26802 13554 26806 13752
rect 26760 12752 26806 13554
rect 26760 12460 26768 12752
rect 26802 12460 26806 12752
rect 26760 11658 26806 12460
rect 27986 13570 28000 13862
rect 28034 13760 28054 13862
rect 29058 13862 29092 13878
rect 27986 13554 28034 13570
rect 29054 13570 29058 13768
rect 30090 13862 30158 14040
rect 30090 13774 30116 13862
rect 29092 13570 29100 13768
rect 27986 12784 28032 13554
rect 27986 12768 28034 12784
rect 27986 12476 28000 12768
rect 27986 12460 28034 12476
rect 29054 12768 29100 13570
rect 29054 12476 29058 12768
rect 29092 12476 29100 12768
rect 26760 11366 26768 11658
rect 26802 11366 26806 11658
rect 26760 10564 26806 11366
rect 27346 12328 27496 12454
rect 27346 11132 27368 12328
rect 27462 11132 27496 12328
rect 27346 10808 27496 11132
rect 27986 11690 28032 12460
rect 27986 11674 28034 11690
rect 27986 11382 28000 11674
rect 27986 11366 28034 11382
rect 29054 11674 29100 12476
rect 29054 11382 29058 11674
rect 29092 11382 29100 11674
rect 26760 10272 26768 10564
rect 26802 10272 26806 10564
rect 26760 9470 26806 10272
rect 27986 10596 28032 11366
rect 27986 10580 28034 10596
rect 27986 10288 28000 10580
rect 27986 10272 28034 10288
rect 29054 10580 29100 11382
rect 29054 10288 29058 10580
rect 29092 10288 29100 10580
rect 27986 9502 28032 10272
rect 27986 9500 28034 9502
rect 26760 9412 26768 9470
rect 26744 9218 26768 9272
rect 25710 9162 25744 9178
rect 26710 9178 26768 9218
rect 26802 9412 26806 9470
rect 27974 9486 28068 9500
rect 27974 9390 28000 9486
rect 26802 9218 26826 9272
rect 26802 9178 26842 9218
rect 26710 9068 26842 9178
rect 27964 9194 28000 9390
rect 28034 9390 28068 9486
rect 29054 9486 29100 10288
rect 29054 9406 29058 9486
rect 28034 9194 28096 9390
rect 22516 8978 26966 9068
rect 22528 8972 26966 8978
rect 24642 8950 24724 8972
rect 23586 8216 23654 8232
rect 25710 8216 25778 8248
rect 21454 8206 25778 8216
rect 21344 8162 25778 8206
rect 21344 8126 25786 8162
rect 21344 8116 25634 8126
rect 21454 7974 21586 8116
rect 19272 7662 19278 7862
rect 20242 7834 20296 7954
rect 20248 7818 20296 7834
rect 19232 6860 19278 7662
rect 19232 6568 19238 6860
rect 19272 6568 19278 6860
rect 19232 5766 19278 6568
rect 19232 5474 19238 5766
rect 19272 5474 19278 5766
rect 19232 4672 19278 5474
rect 19232 4380 19238 4672
rect 19272 4380 19278 4672
rect 19232 3578 19278 4380
rect 19232 3548 19238 3578
rect 18214 3286 18252 3358
rect 18170 3176 18252 3286
rect 19272 3548 19278 3578
rect 20288 7662 20296 7818
rect 20330 7818 20380 7954
rect 21482 7938 21550 7974
rect 20330 7662 20334 7818
rect 20288 6860 20334 7662
rect 20288 6568 20296 6860
rect 20330 6568 20334 6860
rect 20288 5766 20334 6568
rect 21482 7646 21496 7938
rect 21530 7836 21550 7938
rect 22554 7938 22588 7954
rect 21482 7630 21530 7646
rect 22550 7646 22554 7844
rect 23586 7938 23654 8116
rect 23586 7850 23612 7938
rect 22588 7646 22596 7844
rect 21482 6860 21528 7630
rect 21482 6844 21530 6860
rect 21482 6552 21496 6844
rect 21482 6536 21530 6552
rect 22550 6844 22596 7646
rect 22550 6552 22554 6844
rect 22588 6552 22596 6844
rect 20288 5474 20296 5766
rect 20330 5474 20334 5766
rect 20288 4672 20334 5474
rect 20842 6404 20992 6530
rect 20842 5208 20864 6404
rect 20958 5208 20992 6404
rect 20842 4884 20992 5208
rect 21482 5766 21528 6536
rect 21482 5750 21530 5766
rect 21482 5458 21496 5750
rect 21482 5442 21530 5458
rect 22550 5750 22596 6552
rect 22550 5458 22554 5750
rect 22588 5458 22596 5750
rect 20288 4380 20296 4672
rect 20330 4380 20334 4672
rect 20288 3578 20334 4380
rect 20288 3520 20296 3578
rect 19238 3270 19272 3286
rect 20272 3286 20296 3380
rect 20330 3520 20334 3578
rect 21482 4672 21528 5442
rect 21482 4656 21530 4672
rect 21482 4364 21496 4656
rect 21482 4348 21530 4364
rect 22550 4656 22596 5458
rect 22550 4364 22554 4656
rect 22588 4364 22596 4656
rect 21482 3578 21528 4348
rect 21482 3562 21530 3578
rect 21482 3504 21496 3562
rect 20330 3286 20354 3380
rect 20272 3176 20354 3286
rect 22550 3562 22596 4364
rect 22550 3482 22554 3562
rect 21496 3254 21530 3270
rect 22534 3270 22554 3370
rect 22588 3482 22596 3562
rect 23602 7646 23612 7850
rect 23646 7902 23654 7938
rect 24670 7938 24704 7954
rect 23646 7850 23660 7902
rect 23646 7646 23648 7850
rect 23602 6844 23648 7646
rect 23602 6552 23612 6844
rect 23646 6552 23648 6844
rect 23602 5750 23648 6552
rect 23602 5458 23612 5750
rect 23646 5458 23648 5750
rect 23602 4656 23648 5458
rect 23602 4364 23612 4656
rect 23646 4364 23648 4656
rect 23602 3562 23648 4364
rect 23602 3504 23612 3562
rect 22588 3270 22616 3370
rect 3024 3070 7474 3160
rect 9538 3078 13988 3168
rect 16044 3086 20494 3176
rect 16056 3080 20494 3086
rect 22534 3160 22616 3270
rect 23646 3504 23648 3562
rect 25702 7938 25786 8126
rect 24704 7646 24716 7850
rect 25702 7846 25728 7938
rect 24670 6844 24716 7646
rect 24704 6552 24716 6844
rect 24670 5750 24716 6552
rect 24704 5458 24716 5750
rect 24670 4656 24716 5458
rect 24704 4364 24716 4656
rect 24670 3562 24716 4364
rect 23612 3254 23646 3270
rect 24660 3270 24670 3342
rect 24704 3488 24716 3562
rect 25722 7646 25728 7846
rect 25762 7846 25786 7938
rect 26710 7938 26842 8972
rect 27964 8232 28096 9194
rect 29038 9194 29058 9294
rect 29092 9406 29100 9486
rect 30106 13570 30116 13774
rect 30150 13826 30158 13862
rect 31174 13862 31208 13878
rect 30150 13774 30164 13826
rect 30150 13570 30152 13774
rect 30106 12768 30152 13570
rect 30106 12476 30116 12768
rect 30150 12476 30152 12768
rect 30106 11674 30152 12476
rect 30106 11382 30116 11674
rect 30150 11382 30152 11674
rect 30106 10580 30152 11382
rect 30106 10288 30116 10580
rect 30150 10288 30152 10580
rect 30106 9486 30152 10288
rect 30106 9428 30116 9486
rect 29092 9194 29120 9294
rect 29038 9084 29120 9194
rect 30150 9428 30152 9486
rect 32206 13862 32290 14050
rect 31208 13570 31220 13774
rect 32206 13770 32232 13862
rect 31174 12768 31220 13570
rect 31208 12476 31220 12768
rect 31174 11674 31220 12476
rect 31208 11382 31220 11674
rect 31174 10580 31220 11382
rect 31208 10288 31220 10580
rect 31174 9486 31220 10288
rect 30116 9178 30150 9194
rect 31164 9194 31174 9266
rect 31208 9412 31220 9486
rect 32226 13570 32232 13770
rect 32266 13770 32290 13862
rect 33244 13862 33370 14844
rect 34450 14146 34576 15056
rect 35538 15056 35558 15156
rect 35592 15268 35600 15348
rect 36606 19432 36616 19636
rect 36650 19688 36658 19724
rect 37674 19724 37708 19740
rect 36650 19636 36664 19688
rect 36650 19432 36652 19636
rect 36606 18630 36652 19432
rect 36606 18338 36616 18630
rect 36650 18338 36652 18630
rect 36606 17536 36652 18338
rect 36606 17244 36616 17536
rect 36650 17244 36652 17536
rect 36606 16442 36652 17244
rect 36606 16150 36616 16442
rect 36650 16150 36652 16442
rect 36606 15348 36652 16150
rect 36606 15290 36616 15348
rect 35592 15056 35620 15156
rect 35538 14946 35620 15056
rect 36650 15290 36652 15348
rect 38706 19724 38790 19912
rect 37708 19432 37720 19636
rect 38706 19632 38732 19724
rect 37674 18630 37720 19432
rect 37708 18338 37720 18630
rect 37674 17536 37720 18338
rect 37708 17244 37720 17536
rect 37674 16442 37720 17244
rect 37708 16150 37720 16442
rect 37674 15348 37720 16150
rect 36616 15040 36650 15056
rect 37664 15056 37674 15128
rect 37708 15274 37720 15348
rect 38726 19432 38732 19632
rect 38766 19632 38790 19724
rect 39754 19724 39880 20714
rect 40948 20002 41074 20920
rect 42028 20920 42048 21020
rect 42082 21132 42090 21212
rect 43096 25296 43106 25500
rect 43140 25552 43148 25588
rect 44164 25588 44198 25604
rect 43140 25500 43154 25552
rect 43140 25296 43142 25500
rect 43096 24494 43142 25296
rect 43096 24202 43106 24494
rect 43140 24202 43142 24494
rect 43096 23400 43142 24202
rect 43096 23108 43106 23400
rect 43140 23108 43142 23400
rect 43096 22306 43142 23108
rect 43096 22014 43106 22306
rect 43140 22014 43142 22306
rect 43096 21212 43142 22014
rect 43096 21154 43106 21212
rect 42082 20920 42110 21020
rect 42028 20810 42110 20920
rect 43140 21154 43142 21212
rect 45196 25588 45280 25776
rect 44198 25296 44210 25500
rect 45196 25496 45222 25588
rect 44164 24494 44210 25296
rect 44198 24202 44210 24494
rect 44164 23400 44210 24202
rect 44198 23108 44210 23400
rect 44164 22306 44210 23108
rect 44198 22014 44210 22306
rect 44164 21212 44210 22014
rect 43106 20904 43140 20920
rect 44154 20920 44164 20992
rect 44198 21138 44210 21212
rect 45216 25296 45222 25496
rect 45256 25496 45280 25588
rect 46242 25588 46368 26550
rect 47540 25888 47672 26778
rect 48616 26778 48636 26878
rect 48670 26990 48678 27070
rect 49684 31154 49694 31358
rect 49728 31410 49736 31446
rect 50752 31446 50786 31462
rect 49728 31358 49742 31410
rect 49728 31154 49730 31358
rect 49684 30352 49730 31154
rect 49684 30060 49694 30352
rect 49728 30060 49730 30352
rect 49684 29258 49730 30060
rect 49684 28966 49694 29258
rect 49728 28966 49730 29258
rect 49684 28164 49730 28966
rect 49684 27872 49694 28164
rect 49728 27872 49730 28164
rect 49684 27070 49730 27872
rect 49684 27012 49694 27070
rect 48670 26778 48698 26878
rect 48616 26668 48698 26778
rect 49728 27012 49730 27070
rect 51784 31446 51868 31634
rect 50786 31154 50798 31358
rect 51784 31354 51810 31446
rect 50752 30352 50798 31154
rect 50786 30060 50798 30352
rect 50752 29258 50798 30060
rect 50786 28966 50798 29258
rect 50752 28164 50798 28966
rect 50786 27872 50798 28164
rect 50752 27070 50798 27872
rect 49694 26762 49728 26778
rect 50742 26778 50752 26850
rect 50786 26996 50798 27070
rect 51804 31154 51810 31354
rect 51844 31354 51868 31446
rect 52842 31446 52938 32406
rect 54012 31738 54174 32626
rect 55130 32626 55150 32726
rect 55184 32838 55192 32918
rect 56198 37002 56208 37206
rect 56242 37258 56250 37294
rect 57266 37294 57300 37310
rect 56242 37206 56256 37258
rect 56242 37002 56244 37206
rect 56198 36200 56244 37002
rect 56198 35908 56208 36200
rect 56242 35908 56244 36200
rect 56198 35106 56244 35908
rect 56198 34814 56208 35106
rect 56242 34814 56244 35106
rect 56198 34012 56244 34814
rect 56198 33720 56208 34012
rect 56242 33720 56244 34012
rect 56198 32918 56244 33720
rect 56198 32860 56208 32918
rect 55184 32626 55212 32726
rect 55130 32516 55212 32626
rect 56242 32860 56244 32918
rect 58298 37294 58382 37482
rect 57300 37002 57312 37206
rect 58298 37202 58324 37294
rect 57266 36200 57312 37002
rect 57300 35908 57312 36200
rect 57266 35106 57312 35908
rect 57300 34814 57312 35106
rect 57266 34012 57312 34814
rect 57300 33720 57312 34012
rect 57266 32918 57312 33720
rect 56208 32610 56242 32626
rect 57256 32626 57266 32698
rect 57300 32844 57312 32918
rect 58318 37002 58324 37202
rect 58358 37202 58382 37294
rect 59342 37294 59438 38236
rect 58358 37002 58364 37202
rect 59342 37132 59382 37294
rect 58318 36200 58364 37002
rect 58318 35908 58324 36200
rect 58358 35908 58364 36200
rect 58318 35106 58364 35908
rect 58318 34814 58324 35106
rect 58358 34814 58364 35106
rect 58318 34012 58364 34814
rect 58318 33720 58324 34012
rect 58358 33720 58364 34012
rect 58318 32918 58364 33720
rect 58318 32888 58324 32918
rect 57300 32626 57338 32698
rect 57256 32516 57338 32626
rect 58358 32888 58364 32918
rect 59374 37002 59382 37132
rect 59416 37132 59438 37294
rect 59416 37002 59420 37132
rect 59374 36200 59420 37002
rect 59374 35908 59382 36200
rect 59416 35908 59420 36200
rect 59374 35106 59420 35908
rect 59374 34814 59382 35106
rect 59416 34814 59420 35106
rect 59374 34012 59420 34814
rect 59600 35834 60002 36084
rect 59600 34446 59684 35834
rect 59892 34446 60002 35834
rect 76634 35632 76712 38980
rect 76940 35632 76978 38980
rect 76634 35530 76978 35632
rect 77160 38922 77170 39006
rect 77204 39052 77206 39094
rect 77828 39094 77862 39110
rect 77204 39006 77210 39052
rect 77204 38922 77206 39006
rect 77160 38400 77206 38922
rect 77160 38228 77170 38400
rect 77204 38228 77206 38400
rect 77160 37706 77206 38228
rect 77160 37534 77170 37706
rect 77204 37534 77206 37706
rect 77160 37012 77206 37534
rect 77160 36840 77170 37012
rect 77204 36840 77206 37012
rect 77160 36318 77206 36840
rect 77160 36146 77170 36318
rect 77204 36146 77206 36318
rect 77160 35624 77206 36146
rect 77160 35524 77170 35624
rect 77204 35524 77206 35624
rect 77820 38922 77828 39032
rect 78476 39094 78538 39200
rect 78574 39194 78706 39200
rect 77862 38922 77866 39032
rect 78476 39030 78486 39094
rect 77820 38400 77866 38922
rect 77820 38228 77828 38400
rect 77862 38228 77866 38400
rect 77820 37706 77866 38228
rect 77820 37534 77828 37706
rect 77862 37534 77866 37706
rect 77820 37012 77866 37534
rect 77820 36840 77828 37012
rect 77862 36840 77866 37012
rect 77820 36318 77866 36840
rect 77820 36146 77828 36318
rect 77862 36146 77866 36318
rect 77820 35624 77866 36146
rect 77820 35540 77828 35624
rect 77170 35436 77204 35452
rect 77808 35452 77828 35504
rect 77862 35540 77866 35624
rect 78478 38922 78486 39030
rect 78520 39030 78538 39094
rect 79100 39094 79232 39200
rect 78520 38922 78524 39030
rect 79100 38998 79144 39094
rect 78478 38400 78524 38922
rect 78478 38228 78486 38400
rect 78520 38228 78524 38400
rect 78478 37706 78524 38228
rect 78478 37534 78486 37706
rect 78520 37534 78524 37706
rect 78478 37012 78524 37534
rect 78478 36840 78486 37012
rect 78520 36840 78524 37012
rect 78478 36318 78524 36840
rect 78478 36146 78486 36318
rect 78520 36146 78524 36318
rect 78478 35624 78524 36146
rect 78478 35540 78486 35624
rect 77862 35452 77870 35504
rect 77808 35332 77870 35452
rect 78520 35540 78524 35624
rect 79138 38922 79144 38998
rect 79178 38998 79232 39094
rect 79776 39094 79838 39200
rect 80414 39194 83186 39248
rect 83724 39194 86496 39248
rect 80414 39154 80568 39194
rect 79776 39014 79802 39094
rect 79178 38922 79184 38998
rect 79138 38400 79184 38922
rect 79798 38922 79802 39014
rect 79836 39086 79838 39094
rect 80470 39088 80532 39154
rect 79836 38922 79844 39086
rect 79798 38766 79844 38922
rect 79960 38974 80304 39076
rect 80470 39000 80496 39088
rect 79960 38766 80038 38974
rect 79794 38670 80038 38766
rect 79138 38228 79144 38400
rect 79178 38228 79184 38400
rect 79138 37706 79184 38228
rect 79138 37534 79144 37706
rect 79178 37534 79184 37706
rect 79138 37012 79184 37534
rect 79138 36840 79144 37012
rect 79178 36840 79184 37012
rect 79138 36318 79184 36840
rect 79138 36146 79144 36318
rect 79178 36146 79184 36318
rect 79138 35624 79184 36146
rect 79138 35552 79144 35624
rect 78486 35436 78520 35452
rect 79120 35452 79144 35496
rect 79178 35552 79184 35624
rect 79798 38400 79844 38670
rect 79798 38228 79802 38400
rect 79836 38228 79844 38400
rect 79798 37706 79844 38228
rect 79798 37534 79802 37706
rect 79836 37534 79844 37706
rect 79798 37012 79844 37534
rect 79798 36840 79802 37012
rect 79836 36840 79844 37012
rect 79798 36318 79844 36840
rect 79798 36146 79802 36318
rect 79836 36146 79844 36318
rect 79798 35624 79844 36146
rect 79798 35556 79802 35624
rect 79178 35452 79182 35496
rect 79120 35332 79182 35452
rect 79836 35556 79844 35624
rect 79960 35626 80038 38670
rect 80266 35626 80304 38974
rect 79960 35524 80304 35626
rect 80486 38916 80496 39000
rect 80530 39046 80532 39088
rect 81154 39088 81188 39104
rect 80530 39000 80536 39046
rect 80530 38916 80532 39000
rect 80486 38394 80532 38916
rect 80486 38222 80496 38394
rect 80530 38222 80532 38394
rect 80486 37700 80532 38222
rect 80486 37528 80496 37700
rect 80530 37528 80532 37700
rect 80486 37006 80532 37528
rect 80486 36834 80496 37006
rect 80530 36834 80532 37006
rect 80486 36312 80532 36834
rect 80486 36140 80496 36312
rect 80530 36140 80532 36312
rect 80486 35618 80532 36140
rect 80486 35518 80496 35618
rect 79802 35436 79836 35452
rect 80530 35518 80532 35618
rect 81146 38916 81154 39026
rect 81802 39088 81864 39194
rect 81188 38916 81192 39026
rect 81802 39024 81812 39088
rect 81146 38394 81192 38916
rect 81146 38222 81154 38394
rect 81188 38222 81192 38394
rect 81146 37700 81192 38222
rect 81146 37528 81154 37700
rect 81188 37528 81192 37700
rect 81146 37006 81192 37528
rect 81146 36834 81154 37006
rect 81188 36834 81192 37006
rect 81146 36312 81192 36834
rect 81146 36140 81154 36312
rect 81188 36140 81192 36312
rect 81146 35618 81192 36140
rect 81146 35534 81154 35618
rect 80496 35430 80530 35446
rect 81134 35446 81154 35498
rect 81188 35534 81192 35618
rect 81804 38916 81812 39024
rect 81846 39024 81864 39088
rect 82470 39088 82504 39104
rect 81846 38916 81850 39024
rect 81804 38394 81850 38916
rect 81804 38222 81812 38394
rect 81846 38222 81850 38394
rect 81804 37700 81850 38222
rect 81804 37528 81812 37700
rect 81846 37528 81850 37700
rect 81804 37006 81850 37528
rect 81804 36834 81812 37006
rect 81846 36834 81850 37006
rect 81804 36312 81850 36834
rect 81804 36140 81812 36312
rect 81846 36140 81850 36312
rect 81804 35618 81850 36140
rect 81804 35534 81812 35618
rect 81188 35446 81196 35498
rect 77808 35270 79192 35332
rect 77820 35266 79192 35270
rect 81134 35326 81196 35446
rect 81846 35534 81850 35618
rect 82464 38916 82470 39038
rect 83102 39088 83164 39194
rect 83724 39154 83878 39194
rect 85094 39186 85254 39194
rect 82504 38916 82510 39038
rect 83102 39008 83128 39088
rect 82464 38394 82510 38916
rect 82464 38222 82470 38394
rect 82504 38222 82510 38394
rect 82464 37700 82510 38222
rect 82464 37528 82470 37700
rect 82504 37528 82510 37700
rect 82464 37006 82510 37528
rect 82464 36834 82470 37006
rect 82504 36834 82510 37006
rect 82464 36312 82510 36834
rect 82464 36140 82470 36312
rect 82504 36140 82510 36312
rect 82464 35618 82510 36140
rect 82464 35546 82470 35618
rect 81812 35430 81846 35446
rect 82446 35446 82470 35490
rect 82504 35546 82510 35618
rect 83124 38916 83128 39008
rect 83162 39080 83164 39088
rect 83780 39088 83842 39154
rect 83162 38916 83170 39080
rect 83124 38394 83170 38916
rect 83124 38222 83128 38394
rect 83162 38222 83170 38394
rect 83124 37700 83170 38222
rect 83124 37528 83128 37700
rect 83162 37528 83170 37700
rect 83124 37006 83170 37528
rect 83124 36834 83128 37006
rect 83162 36834 83170 37006
rect 83124 36312 83170 36834
rect 83124 36140 83128 36312
rect 83162 36140 83170 36312
rect 83124 35618 83170 36140
rect 83124 35550 83128 35618
rect 82504 35446 82508 35490
rect 82446 35326 82508 35446
rect 83162 35550 83170 35618
rect 83270 38974 83614 39076
rect 83780 39000 83806 39088
rect 83270 35626 83348 38974
rect 83576 35626 83614 38974
rect 83270 35524 83614 35626
rect 83796 38916 83806 39000
rect 83840 39046 83842 39088
rect 84464 39088 84498 39104
rect 83840 39000 83846 39046
rect 83840 38916 83842 39000
rect 83796 38394 83842 38916
rect 83796 38222 83806 38394
rect 83840 38222 83842 38394
rect 83796 37700 83842 38222
rect 83796 37528 83806 37700
rect 83840 37528 83842 37700
rect 83796 37006 83842 37528
rect 83796 36834 83806 37006
rect 83840 36834 83842 37006
rect 83796 36312 83842 36834
rect 83796 36140 83806 36312
rect 83840 36140 83842 36312
rect 83796 35618 83842 36140
rect 83796 35518 83806 35618
rect 83128 35430 83162 35446
rect 83840 35518 83842 35618
rect 84456 38916 84464 39026
rect 85112 39088 85174 39186
rect 84498 38916 84502 39026
rect 85112 39024 85122 39088
rect 84456 38394 84502 38916
rect 84456 38222 84464 38394
rect 84498 38222 84502 38394
rect 84456 37700 84502 38222
rect 84456 37528 84464 37700
rect 84498 37528 84502 37700
rect 84456 37006 84502 37528
rect 84456 36834 84464 37006
rect 84498 36834 84502 37006
rect 84456 36312 84502 36834
rect 84456 36140 84464 36312
rect 84498 36140 84502 36312
rect 84456 35618 84502 36140
rect 84456 35534 84464 35618
rect 83806 35430 83840 35446
rect 84444 35446 84464 35498
rect 84498 35534 84502 35618
rect 85114 38916 85122 39024
rect 85156 39024 85174 39088
rect 85748 39088 85870 39194
rect 85156 38916 85160 39024
rect 85748 39016 85780 39088
rect 85114 38394 85160 38916
rect 85114 38222 85122 38394
rect 85156 38222 85160 38394
rect 85114 37700 85160 38222
rect 85114 37528 85122 37700
rect 85156 37528 85160 37700
rect 85114 37006 85160 37528
rect 85114 36834 85122 37006
rect 85156 36834 85160 37006
rect 85114 36312 85160 36834
rect 85114 36140 85122 36312
rect 85156 36140 85160 36312
rect 85114 35618 85160 36140
rect 85114 35534 85122 35618
rect 84498 35446 84506 35498
rect 84444 35326 84506 35446
rect 85156 35534 85160 35618
rect 85774 38916 85780 39016
rect 85814 39016 85870 39088
rect 86412 39088 86474 39194
rect 85814 38916 85820 39016
rect 86412 39008 86438 39088
rect 86434 38916 86438 39008
rect 86472 39080 86474 39088
rect 86472 38916 86480 39080
rect 86696 38916 86742 39284
rect 85774 38394 85820 38916
rect 86430 38844 86742 38916
rect 85774 38222 85780 38394
rect 85814 38222 85820 38394
rect 85774 37700 85820 38222
rect 85774 37528 85780 37700
rect 85814 37528 85820 37700
rect 85774 37006 85820 37528
rect 85774 36834 85780 37006
rect 85814 36834 85820 37006
rect 85774 36312 85820 36834
rect 85774 36140 85780 36312
rect 85814 36140 85820 36312
rect 85774 35618 85820 36140
rect 85774 35546 85780 35618
rect 85122 35430 85156 35446
rect 85756 35446 85780 35490
rect 85814 35546 85820 35618
rect 86434 38394 86480 38844
rect 86434 38222 86438 38394
rect 86472 38222 86480 38394
rect 86434 37700 86480 38222
rect 86434 37528 86438 37700
rect 86472 37528 86480 37700
rect 86434 37006 86480 37528
rect 86434 36834 86438 37006
rect 86472 36834 86480 37006
rect 86434 36312 86480 36834
rect 86434 36140 86438 36312
rect 86472 36140 86480 36312
rect 86434 35618 86480 36140
rect 86434 35550 86438 35618
rect 85814 35446 85818 35490
rect 85756 35326 85818 35446
rect 86472 35550 86480 35618
rect 86438 35430 86472 35446
rect 86696 35360 86742 38844
rect 86978 35360 87008 39284
rect 78196 35100 78270 35266
rect 79120 35262 79182 35266
rect 81134 35264 82518 35326
rect 84444 35264 85828 35326
rect 81146 35260 82518 35264
rect 84456 35260 85828 35264
rect 81522 35094 81596 35260
rect 82446 35256 82508 35260
rect 84832 35094 84906 35260
rect 85756 35256 85818 35260
rect 86696 35242 87008 35360
rect 59600 34156 60002 34446
rect 59374 33720 59382 34012
rect 59416 33720 59420 34012
rect 59374 32918 59420 33720
rect 59374 32860 59382 32918
rect 59358 32702 59382 32720
rect 58324 32610 58358 32626
rect 59350 32626 59382 32702
rect 59416 32860 59420 32918
rect 59416 32702 59440 32720
rect 59416 32626 59446 32702
rect 59350 32516 59446 32626
rect 55130 32426 59580 32516
rect 55142 32420 59580 32426
rect 57256 32398 57338 32420
rect 56182 31738 56250 31754
rect 58306 31738 58374 31770
rect 54012 31728 58374 31738
rect 53940 31684 58374 31728
rect 53940 31648 58382 31684
rect 53940 31638 58230 31648
rect 52842 31364 52868 31446
rect 51844 31154 51850 31354
rect 51804 30352 51850 31154
rect 51804 30060 51810 30352
rect 51844 30060 51850 30352
rect 51804 29258 51850 30060
rect 51804 28966 51810 29258
rect 51844 28966 51850 29258
rect 51804 28164 51850 28966
rect 51804 27872 51810 28164
rect 51844 27872 51850 28164
rect 51804 27070 51850 27872
rect 51804 27040 51810 27070
rect 50786 26778 50824 26850
rect 50742 26668 50824 26778
rect 51844 27040 51850 27070
rect 52860 31154 52868 31364
rect 52902 31364 52938 31446
rect 54012 31460 54174 31638
rect 54012 31398 54092 31460
rect 52902 31154 52906 31364
rect 52860 30352 52906 31154
rect 52860 30060 52868 30352
rect 52902 30060 52906 30352
rect 52860 29258 52906 30060
rect 54078 31168 54092 31398
rect 54126 31398 54174 31460
rect 55150 31460 55184 31476
rect 54126 31358 54146 31398
rect 54078 31152 54126 31168
rect 55146 31168 55150 31366
rect 56182 31460 56250 31638
rect 56182 31372 56208 31460
rect 55184 31168 55192 31366
rect 54078 30382 54124 31152
rect 54078 30366 54126 30382
rect 54078 30074 54092 30366
rect 54078 30058 54126 30074
rect 55146 30366 55192 31168
rect 55146 30074 55150 30366
rect 55184 30074 55192 30366
rect 52860 28966 52868 29258
rect 52902 28966 52906 29258
rect 52860 28164 52906 28966
rect 53438 29926 53588 30052
rect 53438 28730 53460 29926
rect 53554 28730 53588 29926
rect 53438 28406 53588 28730
rect 54078 29288 54124 30058
rect 54078 29272 54126 29288
rect 54078 28980 54092 29272
rect 54078 28964 54126 28980
rect 55146 29272 55192 30074
rect 55146 28980 55150 29272
rect 55184 28980 55192 29272
rect 52860 27872 52868 28164
rect 52902 27872 52906 28164
rect 52860 27070 52906 27872
rect 52860 27012 52868 27070
rect 52844 26840 52868 26872
rect 51810 26762 51844 26778
rect 52836 26778 52868 26840
rect 52902 27012 52906 27070
rect 54078 28194 54124 28964
rect 54078 28178 54126 28194
rect 54078 27886 54092 28178
rect 54078 27870 54126 27886
rect 55146 28178 55192 28980
rect 55146 27886 55150 28178
rect 55184 27886 55192 28178
rect 54078 27106 54124 27870
rect 54078 27084 54174 27106
rect 52902 26840 52926 26872
rect 52902 26778 52932 26840
rect 52836 26668 52932 26778
rect 54078 26792 54092 27084
rect 54126 26792 54174 27084
rect 55146 27084 55192 27886
rect 55146 27004 55150 27084
rect 48616 26578 53066 26668
rect 48628 26572 53066 26578
rect 50742 26550 50824 26572
rect 49668 25888 49736 25904
rect 51792 25888 51860 25920
rect 47540 25878 51860 25888
rect 47426 25834 51860 25878
rect 47426 25798 51868 25834
rect 47426 25788 51716 25798
rect 47540 25686 47672 25788
rect 45256 25296 45262 25496
rect 46242 25480 46280 25588
rect 45216 24494 45262 25296
rect 45216 24202 45222 24494
rect 45256 24202 45262 24494
rect 45216 23400 45262 24202
rect 45216 23108 45222 23400
rect 45256 23108 45262 23400
rect 45216 22306 45262 23108
rect 45216 22014 45222 22306
rect 45256 22014 45262 22306
rect 45216 21212 45262 22014
rect 45216 21182 45222 21212
rect 44198 20920 44236 20992
rect 44154 20810 44236 20920
rect 45256 21182 45262 21212
rect 46272 25296 46280 25480
rect 46314 25480 46368 25588
rect 47564 25610 47632 25686
rect 46314 25296 46318 25480
rect 46272 24494 46318 25296
rect 46272 24202 46280 24494
rect 46314 24202 46318 24494
rect 47564 25318 47578 25610
rect 47612 25508 47632 25610
rect 48636 25610 48670 25626
rect 47564 25302 47612 25318
rect 48632 25318 48636 25516
rect 49668 25610 49736 25788
rect 49668 25522 49694 25610
rect 48670 25318 48678 25516
rect 47564 24532 47610 25302
rect 47564 24516 47612 24532
rect 47564 24224 47578 24516
rect 47564 24208 47612 24224
rect 48632 24516 48678 25318
rect 48632 24224 48636 24516
rect 48670 24224 48678 24516
rect 46272 23400 46318 24202
rect 46272 23108 46280 23400
rect 46314 23108 46318 23400
rect 46272 22306 46318 23108
rect 46924 24076 47074 24202
rect 46924 22880 46946 24076
rect 47040 22880 47074 24076
rect 46924 22556 47074 22880
rect 47564 23438 47610 24208
rect 47564 23422 47612 23438
rect 47564 23130 47578 23422
rect 47564 23114 47612 23130
rect 48632 23422 48678 24224
rect 48632 23130 48636 23422
rect 48670 23130 48678 23422
rect 46272 22014 46280 22306
rect 46314 22014 46318 22306
rect 46272 21212 46318 22014
rect 46272 21154 46280 21212
rect 46256 20998 46280 21014
rect 45222 20904 45256 20920
rect 46242 20920 46280 20998
rect 46314 21154 46318 21212
rect 47564 22344 47610 23114
rect 47564 22328 47612 22344
rect 47564 22036 47578 22328
rect 47564 22020 47612 22036
rect 48632 22328 48678 23130
rect 48632 22036 48636 22328
rect 48670 22036 48678 22328
rect 47564 21250 47610 22020
rect 47564 21234 47612 21250
rect 47564 21176 47578 21234
rect 46314 20998 46338 21014
rect 46314 20920 46368 20998
rect 46242 20810 46368 20920
rect 47548 20942 47578 21094
rect 48632 21234 48678 22036
rect 48632 21154 48636 21234
rect 47612 20942 47680 21094
rect 42028 20720 46478 20810
rect 42040 20714 46478 20720
rect 44154 20692 44236 20714
rect 43080 20002 43148 20018
rect 45204 20002 45272 20034
rect 40948 19992 45272 20002
rect 40838 19948 45272 19992
rect 40838 19912 45280 19948
rect 40838 19902 45128 19912
rect 40948 19724 41074 19902
rect 42048 19724 42082 19740
rect 38766 19432 38772 19632
rect 39754 19574 39790 19724
rect 38726 18630 38772 19432
rect 38726 18338 38732 18630
rect 38766 18338 38772 18630
rect 38726 17536 38772 18338
rect 38726 17244 38732 17536
rect 38766 17244 38772 17536
rect 38726 16442 38772 17244
rect 38726 16150 38732 16442
rect 38766 16150 38772 16442
rect 38726 15348 38772 16150
rect 38726 15318 38732 15348
rect 37708 15056 37746 15128
rect 37664 14946 37746 15056
rect 38766 15318 38772 15348
rect 39782 19432 39790 19574
rect 39824 19574 39880 19724
rect 39824 19432 39828 19574
rect 39782 18630 39828 19432
rect 39782 18338 39790 18630
rect 39824 18338 39828 18630
rect 39782 17536 39828 18338
rect 40976 19432 40990 19724
rect 41024 19622 41044 19724
rect 40976 19416 41024 19432
rect 42044 19432 42048 19630
rect 43080 19724 43148 19902
rect 43080 19636 43106 19724
rect 42082 19432 42090 19630
rect 40976 18646 41022 19416
rect 40976 18630 41024 18646
rect 40976 18338 40990 18630
rect 40976 18322 41024 18338
rect 42044 18630 42090 19432
rect 42044 18338 42048 18630
rect 42082 18338 42090 18630
rect 39782 17244 39790 17536
rect 39824 17244 39828 17536
rect 39782 16442 39828 17244
rect 40336 18190 40486 18316
rect 40336 16994 40358 18190
rect 40452 16994 40486 18190
rect 40336 16670 40486 16994
rect 40976 17552 41022 18322
rect 40976 17536 41024 17552
rect 40976 17244 40990 17536
rect 40976 17228 41024 17244
rect 42044 17536 42090 18338
rect 42044 17244 42048 17536
rect 42082 17244 42090 17536
rect 39782 16150 39790 16442
rect 39824 16150 39828 16442
rect 39782 15348 39828 16150
rect 39782 15290 39790 15348
rect 38732 15040 38766 15056
rect 39766 15056 39790 15150
rect 39824 15290 39828 15348
rect 40976 16458 41022 17228
rect 40976 16442 41024 16458
rect 40976 16150 40990 16442
rect 40976 16134 41024 16150
rect 42044 16442 42090 17244
rect 42044 16150 42048 16442
rect 42082 16150 42090 16442
rect 40976 15364 41022 16134
rect 40976 15348 41024 15364
rect 40976 15290 40990 15348
rect 39824 15080 39848 15150
rect 39824 15056 39894 15080
rect 39766 14946 39894 15056
rect 40976 15056 40990 15256
rect 42044 15348 42090 16150
rect 42044 15268 42048 15348
rect 41024 15056 41102 15256
rect 35538 14856 39988 14946
rect 35550 14850 39988 14856
rect 37664 14828 37746 14850
rect 36600 14146 36668 14162
rect 38724 14146 38792 14178
rect 34450 14136 38792 14146
rect 34358 14092 38792 14136
rect 34358 14056 38800 14092
rect 34358 14046 38648 14056
rect 34450 13868 34576 14046
rect 34450 13864 34510 13868
rect 32266 13570 32272 13770
rect 33244 13654 33290 13862
rect 32226 12768 32272 13570
rect 32226 12476 32232 12768
rect 32266 12476 32272 12768
rect 32226 11674 32272 12476
rect 32226 11382 32232 11674
rect 32266 11382 32272 11674
rect 32226 10580 32272 11382
rect 32226 10288 32232 10580
rect 32266 10288 32272 10580
rect 32226 9486 32272 10288
rect 32226 9456 32232 9486
rect 31208 9194 31246 9266
rect 31164 9084 31246 9194
rect 32266 9456 32272 9486
rect 33282 13570 33290 13654
rect 33324 13654 33370 13862
rect 33324 13570 33328 13654
rect 33282 12768 33328 13570
rect 33282 12476 33290 12768
rect 33324 12476 33328 12768
rect 33282 11674 33328 12476
rect 34496 13576 34510 13864
rect 34544 13864 34576 13868
rect 35568 13868 35602 13884
rect 34544 13766 34564 13864
rect 34496 13560 34544 13576
rect 35564 13576 35568 13774
rect 36600 13868 36668 14046
rect 36600 13780 36626 13868
rect 35602 13576 35610 13774
rect 34496 12790 34542 13560
rect 34496 12774 34544 12790
rect 34496 12482 34510 12774
rect 34496 12466 34544 12482
rect 35564 12774 35610 13576
rect 35564 12482 35568 12774
rect 35602 12482 35610 12774
rect 33282 11382 33290 11674
rect 33324 11382 33328 11674
rect 33282 10580 33328 11382
rect 33856 12334 34006 12460
rect 33856 11138 33878 12334
rect 33972 11138 34006 12334
rect 33856 10814 34006 11138
rect 34496 11696 34542 12466
rect 34496 11680 34544 11696
rect 34496 11388 34510 11680
rect 34496 11372 34544 11388
rect 35564 11680 35610 12482
rect 35564 11388 35568 11680
rect 35602 11388 35610 11680
rect 33282 10288 33290 10580
rect 33324 10288 33328 10580
rect 33282 9486 33328 10288
rect 33282 9428 33290 9486
rect 33266 9202 33290 9288
rect 32232 9178 32266 9194
rect 33258 9194 33290 9202
rect 33324 9428 33328 9486
rect 34496 10602 34542 11372
rect 34496 10586 34544 10602
rect 34496 10294 34510 10586
rect 34496 10278 34544 10294
rect 35564 10586 35610 11388
rect 35564 10294 35568 10586
rect 35602 10294 35610 10586
rect 34496 9508 34542 10278
rect 34496 9492 34544 9508
rect 34496 9434 34510 9492
rect 33324 9202 33348 9288
rect 33324 9194 33384 9202
rect 33258 9084 33384 9194
rect 34466 9200 34510 9342
rect 35564 9492 35610 10294
rect 35564 9412 35568 9492
rect 34544 9200 34592 9342
rect 29038 8994 33488 9084
rect 29050 8988 33488 8994
rect 31164 8966 31246 8988
rect 30108 8232 30176 8248
rect 32232 8232 32300 8264
rect 27964 8222 32300 8232
rect 27866 8178 32300 8222
rect 27866 8142 32308 8178
rect 27866 8132 32156 8142
rect 27964 7982 28096 8132
rect 25762 7646 25768 7846
rect 26710 7810 26786 7938
rect 25722 6844 25768 7646
rect 25722 6552 25728 6844
rect 25762 6552 25768 6844
rect 25722 5750 25768 6552
rect 25722 5458 25728 5750
rect 25762 5458 25768 5750
rect 25722 4656 25768 5458
rect 25722 4364 25728 4656
rect 25762 4364 25768 4656
rect 25722 3562 25768 4364
rect 25722 3532 25728 3562
rect 24704 3270 24742 3342
rect 24660 3160 24742 3270
rect 25762 3532 25768 3562
rect 26778 7646 26786 7810
rect 26820 7810 26842 7938
rect 28004 7954 28072 7982
rect 26820 7646 26824 7810
rect 26778 6844 26824 7646
rect 26778 6552 26786 6844
rect 26820 6552 26824 6844
rect 26778 5750 26824 6552
rect 28004 7662 28018 7954
rect 28052 7852 28072 7954
rect 29076 7954 29110 7970
rect 28004 7646 28052 7662
rect 29072 7662 29076 7860
rect 30108 7954 30176 8132
rect 30108 7866 30134 7954
rect 29110 7662 29118 7860
rect 28004 6876 28050 7646
rect 28004 6860 28052 6876
rect 28004 6568 28018 6860
rect 28004 6552 28052 6568
rect 29072 6860 29118 7662
rect 29072 6568 29076 6860
rect 29110 6568 29118 6860
rect 26778 5458 26786 5750
rect 26820 5458 26824 5750
rect 26778 4656 26824 5458
rect 27364 6420 27514 6546
rect 27364 5224 27386 6420
rect 27480 5224 27514 6420
rect 27364 4900 27514 5224
rect 28004 5782 28050 6552
rect 28004 5766 28052 5782
rect 28004 5474 28018 5766
rect 28004 5458 28052 5474
rect 29072 5766 29118 6568
rect 29072 5474 29076 5766
rect 29110 5474 29118 5766
rect 26778 4364 26786 4656
rect 26820 4364 26824 4656
rect 26778 3562 26824 4364
rect 26778 3504 26786 3562
rect 25728 3254 25762 3270
rect 26762 3270 26786 3364
rect 26820 3504 26824 3562
rect 28004 4688 28050 5458
rect 28004 4672 28052 4688
rect 28004 4380 28018 4672
rect 28004 4364 28052 4380
rect 29072 4672 29118 5474
rect 29072 4380 29076 4672
rect 29110 4380 29118 4672
rect 28004 3594 28050 4364
rect 28004 3578 28052 3594
rect 28004 3520 28018 3578
rect 26820 3270 26844 3364
rect 29072 3578 29118 4380
rect 29072 3498 29076 3578
rect 28018 3270 28052 3286
rect 29056 3286 29076 3386
rect 29110 3498 29118 3578
rect 30124 7662 30134 7866
rect 30168 7918 30176 7954
rect 31192 7954 31226 7970
rect 30168 7866 30182 7918
rect 30168 7662 30170 7866
rect 30124 6860 30170 7662
rect 30124 6568 30134 6860
rect 30168 6568 30170 6860
rect 30124 5766 30170 6568
rect 30124 5474 30134 5766
rect 30168 5474 30170 5766
rect 30124 4672 30170 5474
rect 30124 4380 30134 4672
rect 30168 4380 30170 4672
rect 30124 3578 30170 4380
rect 30124 3520 30134 3578
rect 29110 3286 29138 3386
rect 26762 3164 26844 3270
rect 29056 3176 29138 3286
rect 30168 3520 30170 3578
rect 32224 7954 32308 8142
rect 31226 7662 31238 7866
rect 32224 7862 32250 7954
rect 31192 6860 31238 7662
rect 31226 6568 31238 6860
rect 31192 5766 31238 6568
rect 31226 5474 31238 5766
rect 31192 4672 31238 5474
rect 31226 4380 31238 4672
rect 31192 3578 31238 4380
rect 30134 3270 30168 3286
rect 31182 3286 31192 3358
rect 31226 3504 31238 3578
rect 32244 7662 32250 7862
rect 32284 7862 32308 7954
rect 33258 7954 33384 8988
rect 34466 8238 34592 9200
rect 35548 9200 35568 9300
rect 35602 9412 35610 9492
rect 36616 13576 36626 13780
rect 36660 13832 36668 13868
rect 37684 13868 37718 13884
rect 36660 13780 36674 13832
rect 36660 13576 36662 13780
rect 36616 12774 36662 13576
rect 36616 12482 36626 12774
rect 36660 12482 36662 12774
rect 36616 11680 36662 12482
rect 36616 11388 36626 11680
rect 36660 11388 36662 11680
rect 36616 10586 36662 11388
rect 36616 10294 36626 10586
rect 36660 10294 36662 10586
rect 36616 9492 36662 10294
rect 36616 9434 36626 9492
rect 35602 9200 35630 9300
rect 35548 9090 35630 9200
rect 36660 9434 36662 9492
rect 38716 13868 38800 14056
rect 37718 13576 37730 13780
rect 38716 13776 38742 13868
rect 37684 12774 37730 13576
rect 37718 12482 37730 12774
rect 37684 11680 37730 12482
rect 37718 11388 37730 11680
rect 37684 10586 37730 11388
rect 37718 10294 37730 10586
rect 37684 9492 37730 10294
rect 36626 9184 36660 9200
rect 37674 9200 37684 9272
rect 37718 9418 37730 9492
rect 38736 13576 38742 13776
rect 38776 13776 38800 13868
rect 39768 13868 39894 14850
rect 40976 14146 41102 15056
rect 42028 15056 42048 15156
rect 42082 15268 42090 15348
rect 43096 19432 43106 19636
rect 43140 19688 43148 19724
rect 44164 19724 44198 19740
rect 43140 19636 43154 19688
rect 43140 19432 43142 19636
rect 43096 18630 43142 19432
rect 43096 18338 43106 18630
rect 43140 18338 43142 18630
rect 43096 17536 43142 18338
rect 43096 17244 43106 17536
rect 43140 17244 43142 17536
rect 43096 16442 43142 17244
rect 43096 16150 43106 16442
rect 43140 16150 43142 16442
rect 43096 15348 43142 16150
rect 43096 15290 43106 15348
rect 42082 15056 42110 15156
rect 42028 14946 42110 15056
rect 43140 15290 43142 15348
rect 45196 19724 45280 19912
rect 44198 19432 44210 19636
rect 45196 19632 45222 19724
rect 44164 18630 44210 19432
rect 44198 18338 44210 18630
rect 44164 17536 44210 18338
rect 44198 17244 44210 17536
rect 44164 16442 44210 17244
rect 44198 16150 44210 16442
rect 44164 15348 44210 16150
rect 43106 15040 43140 15056
rect 44154 15056 44164 15128
rect 44198 15274 44210 15348
rect 45216 19432 45222 19632
rect 45256 19632 45280 19724
rect 46242 19724 46368 20714
rect 47548 20024 47680 20942
rect 48616 20942 48636 21042
rect 48670 21154 48678 21234
rect 49684 25318 49694 25522
rect 49728 25574 49736 25610
rect 50752 25610 50786 25626
rect 49728 25522 49742 25574
rect 49728 25318 49730 25522
rect 49684 24516 49730 25318
rect 49684 24224 49694 24516
rect 49728 24224 49730 24516
rect 49684 23422 49730 24224
rect 49684 23130 49694 23422
rect 49728 23130 49730 23422
rect 49684 22328 49730 23130
rect 49684 22036 49694 22328
rect 49728 22036 49730 22328
rect 49684 21234 49730 22036
rect 49684 21176 49694 21234
rect 48670 20942 48698 21042
rect 48616 20832 48698 20942
rect 49728 21176 49730 21234
rect 51784 25610 51868 25798
rect 50786 25318 50798 25522
rect 51784 25518 51810 25610
rect 50752 24516 50798 25318
rect 50786 24224 50798 24516
rect 50752 23422 50798 24224
rect 50786 23130 50798 23422
rect 50752 22328 50798 23130
rect 50786 22036 50798 22328
rect 50752 21234 50798 22036
rect 49694 20926 49728 20942
rect 50742 20942 50752 21014
rect 50786 21160 50798 21234
rect 51804 25318 51810 25518
rect 51844 25518 51868 25610
rect 52836 25610 52932 26572
rect 54078 25902 54174 26792
rect 55130 26792 55150 26892
rect 55184 27004 55192 27084
rect 56198 31168 56208 31372
rect 56242 31424 56250 31460
rect 57266 31460 57300 31476
rect 56242 31372 56256 31424
rect 56242 31168 56244 31372
rect 56198 30366 56244 31168
rect 56198 30074 56208 30366
rect 56242 30074 56244 30366
rect 56198 29272 56244 30074
rect 56198 28980 56208 29272
rect 56242 28980 56244 29272
rect 56198 28178 56244 28980
rect 56198 27886 56208 28178
rect 56242 27886 56244 28178
rect 56198 27084 56244 27886
rect 56198 27026 56208 27084
rect 55184 26792 55212 26892
rect 55130 26682 55212 26792
rect 56242 27026 56244 27084
rect 58298 31460 58382 31648
rect 57300 31168 57312 31372
rect 58298 31368 58324 31460
rect 57266 30366 57312 31168
rect 57300 30074 57312 30366
rect 57266 29272 57312 30074
rect 57300 28980 57312 29272
rect 57266 28178 57312 28980
rect 57300 27886 57312 28178
rect 57266 27084 57312 27886
rect 56208 26776 56242 26792
rect 57256 26792 57266 26864
rect 57300 27010 57312 27084
rect 58318 31168 58324 31368
rect 58358 31368 58382 31460
rect 59350 31460 59446 32420
rect 58358 31168 58364 31368
rect 59350 31364 59382 31460
rect 58318 30366 58364 31168
rect 58318 30074 58324 30366
rect 58358 30074 58364 30366
rect 58318 29272 58364 30074
rect 58318 28980 58324 29272
rect 58358 28980 58364 29272
rect 58318 28178 58364 28980
rect 58318 27886 58324 28178
rect 58358 27886 58364 28178
rect 58318 27084 58364 27886
rect 58318 27054 58324 27084
rect 57300 26792 57338 26864
rect 57256 26682 57338 26792
rect 58358 27054 58364 27084
rect 59374 31168 59382 31364
rect 59416 31364 59446 31460
rect 59416 31168 59420 31364
rect 59374 30366 59420 31168
rect 59374 30074 59382 30366
rect 59416 30074 59420 30366
rect 59374 29272 59420 30074
rect 59374 28980 59382 29272
rect 59416 28980 59420 29272
rect 59374 28178 59420 28980
rect 59374 27886 59382 28178
rect 59416 27886 59420 28178
rect 59586 29896 60030 30090
rect 59586 28426 59642 29896
rect 59974 28426 60030 29896
rect 59586 28134 60030 28426
rect 59374 27084 59420 27886
rect 59374 27026 59382 27084
rect 59358 26884 59382 26886
rect 58324 26776 58358 26792
rect 59356 26792 59382 26884
rect 59416 27026 59420 27084
rect 59416 26884 59440 26886
rect 59416 26792 59452 26884
rect 59356 26682 59452 26792
rect 55130 26592 59580 26682
rect 55142 26586 59580 26592
rect 57256 26564 57338 26586
rect 56182 25902 56250 25918
rect 58306 25902 58374 25934
rect 54078 25892 58374 25902
rect 53940 25848 58374 25892
rect 53940 25812 58382 25848
rect 53940 25802 58230 25812
rect 51844 25318 51850 25518
rect 52836 25502 52868 25610
rect 51804 24516 51850 25318
rect 51804 24224 51810 24516
rect 51844 24224 51850 24516
rect 51804 23422 51850 24224
rect 51804 23130 51810 23422
rect 51844 23130 51850 23422
rect 51804 22328 51850 23130
rect 51804 22036 51810 22328
rect 51844 22036 51850 22328
rect 51804 21234 51850 22036
rect 51804 21204 51810 21234
rect 50786 20942 50824 21014
rect 50742 20832 50824 20942
rect 51844 21204 51850 21234
rect 52860 25318 52868 25502
rect 52902 25502 52932 25610
rect 54078 25768 54174 25802
rect 54078 25624 54146 25768
rect 52902 25318 52906 25502
rect 52860 24516 52906 25318
rect 52860 24224 52868 24516
rect 52902 24224 52906 24516
rect 52860 23422 52906 24224
rect 54078 25332 54092 25624
rect 54126 25522 54146 25624
rect 55150 25624 55184 25640
rect 54078 25316 54126 25332
rect 55146 25332 55150 25530
rect 56182 25624 56250 25802
rect 56182 25536 56208 25624
rect 55184 25332 55192 25530
rect 54078 24546 54124 25316
rect 54078 24530 54126 24546
rect 54078 24238 54092 24530
rect 54078 24222 54126 24238
rect 55146 24530 55192 25332
rect 55146 24238 55150 24530
rect 55184 24238 55192 24530
rect 52860 23130 52868 23422
rect 52902 23130 52906 23422
rect 52860 22328 52906 23130
rect 53438 24090 53588 24216
rect 53438 22894 53460 24090
rect 53554 22894 53588 24090
rect 53438 22570 53588 22894
rect 54078 23452 54124 24222
rect 54078 23436 54126 23452
rect 54078 23144 54092 23436
rect 54078 23128 54126 23144
rect 55146 23436 55192 24238
rect 55146 23144 55150 23436
rect 55184 23144 55192 23436
rect 52860 22036 52868 22328
rect 52902 22036 52906 22328
rect 52860 21234 52906 22036
rect 52860 21176 52868 21234
rect 51810 20926 51844 20942
rect 52844 20942 52868 21036
rect 52902 21176 52906 21234
rect 54078 22358 54124 23128
rect 54078 22342 54126 22358
rect 54078 22050 54092 22342
rect 54078 22034 54126 22050
rect 55146 22342 55192 23144
rect 55146 22050 55150 22342
rect 55184 22050 55192 22342
rect 54078 21264 54124 22034
rect 54078 21248 54126 21264
rect 54078 21190 54092 21248
rect 52902 20970 52926 21036
rect 52902 20942 52954 20970
rect 52844 20832 52954 20942
rect 54024 20956 54092 21070
rect 55146 21248 55192 22050
rect 55146 21168 55150 21248
rect 54126 20956 54150 21070
rect 48616 20742 53066 20832
rect 48628 20736 53066 20742
rect 50742 20714 50824 20736
rect 49668 20024 49736 20040
rect 51792 20024 51860 20056
rect 47548 20014 51860 20024
rect 47426 19970 51860 20014
rect 47426 19934 51868 19970
rect 47426 19924 51716 19934
rect 45256 19432 45262 19632
rect 46242 19614 46280 19724
rect 45216 18630 45262 19432
rect 45216 18338 45222 18630
rect 45256 18338 45262 18630
rect 45216 17536 45262 18338
rect 45216 17244 45222 17536
rect 45256 17244 45262 17536
rect 45216 16442 45262 17244
rect 45216 16150 45222 16442
rect 45256 16150 45262 16442
rect 45216 15348 45262 16150
rect 45216 15318 45222 15348
rect 44198 15056 44236 15128
rect 44154 14946 44236 15056
rect 45256 15318 45262 15348
rect 46272 19432 46280 19614
rect 46314 19614 46368 19724
rect 47548 19746 47680 19924
rect 47548 19686 47578 19746
rect 46314 19432 46318 19614
rect 46272 18630 46318 19432
rect 46272 18338 46280 18630
rect 46314 18338 46318 18630
rect 47564 19454 47578 19686
rect 47612 19686 47680 19746
rect 48636 19746 48670 19762
rect 47612 19644 47632 19686
rect 47564 19438 47612 19454
rect 48632 19454 48636 19652
rect 49668 19746 49736 19924
rect 49668 19658 49694 19746
rect 48670 19454 48678 19652
rect 47564 18668 47610 19438
rect 47564 18652 47612 18668
rect 47564 18360 47578 18652
rect 47564 18344 47612 18360
rect 48632 18652 48678 19454
rect 48632 18360 48636 18652
rect 48670 18360 48678 18652
rect 46272 17536 46318 18338
rect 46272 17244 46280 17536
rect 46314 17244 46318 17536
rect 46272 16442 46318 17244
rect 46924 18212 47074 18338
rect 46924 17016 46946 18212
rect 47040 17016 47074 18212
rect 46924 16692 47074 17016
rect 47564 17574 47610 18344
rect 47564 17558 47612 17574
rect 47564 17266 47578 17558
rect 47564 17250 47612 17266
rect 48632 17558 48678 18360
rect 48632 17266 48636 17558
rect 48670 17266 48678 17558
rect 46272 16150 46280 16442
rect 46314 16150 46318 16442
rect 46272 15348 46318 16150
rect 46272 15290 46280 15348
rect 45222 15040 45256 15056
rect 46256 15056 46280 15150
rect 46314 15290 46318 15348
rect 47564 16480 47610 17250
rect 47564 16464 47612 16480
rect 47564 16172 47578 16464
rect 47564 16156 47612 16172
rect 48632 16464 48678 17266
rect 48632 16172 48636 16464
rect 48670 16172 48678 16464
rect 47564 15386 47610 16156
rect 47564 15370 47612 15386
rect 47564 15312 47578 15370
rect 46314 15056 46338 15150
rect 46256 15032 46338 15056
rect 47528 15078 47578 15276
rect 48632 15370 48678 16172
rect 48632 15290 48636 15370
rect 47612 15078 47654 15276
rect 46256 14946 46382 15032
rect 42028 14856 46478 14946
rect 42040 14850 46478 14856
rect 44154 14828 44236 14850
rect 43090 14146 43158 14162
rect 45214 14146 45282 14178
rect 40976 14136 45282 14146
rect 40848 14092 45282 14136
rect 40848 14056 45290 14092
rect 40848 14046 45138 14056
rect 40976 13872 41102 14046
rect 38776 13576 38782 13776
rect 39768 13696 39800 13868
rect 38736 12774 38782 13576
rect 38736 12482 38742 12774
rect 38776 12482 38782 12774
rect 38736 11680 38782 12482
rect 38736 11388 38742 11680
rect 38776 11388 38782 11680
rect 38736 10586 38782 11388
rect 38736 10294 38742 10586
rect 38776 10294 38782 10586
rect 38736 9492 38782 10294
rect 38736 9462 38742 9492
rect 37718 9200 37756 9272
rect 37674 9090 37756 9200
rect 38776 9462 38782 9492
rect 39792 13576 39800 13696
rect 39834 13696 39894 13868
rect 40986 13868 41054 13872
rect 39834 13576 39838 13696
rect 39792 12774 39838 13576
rect 39792 12482 39800 12774
rect 39834 12482 39838 12774
rect 39792 11680 39838 12482
rect 40986 13576 41000 13868
rect 41034 13766 41054 13868
rect 42058 13868 42092 13884
rect 40986 13560 41034 13576
rect 42054 13576 42058 13774
rect 43090 13868 43158 14046
rect 43090 13780 43116 13868
rect 42092 13576 42100 13774
rect 40986 12790 41032 13560
rect 40986 12774 41034 12790
rect 40986 12482 41000 12774
rect 40986 12466 41034 12482
rect 42054 12774 42100 13576
rect 42054 12482 42058 12774
rect 42092 12482 42100 12774
rect 39792 11388 39800 11680
rect 39834 11388 39838 11680
rect 39792 10586 39838 11388
rect 40346 12334 40496 12460
rect 40346 11138 40368 12334
rect 40462 11138 40496 12334
rect 40346 10814 40496 11138
rect 40986 11696 41032 12466
rect 40986 11680 41034 11696
rect 40986 11388 41000 11680
rect 40986 11372 41034 11388
rect 42054 11680 42100 12482
rect 42054 11388 42058 11680
rect 42092 11388 42100 11680
rect 39792 10294 39800 10586
rect 39834 10294 39838 10586
rect 39792 9492 39838 10294
rect 39792 9434 39800 9492
rect 38742 9184 38776 9200
rect 39776 9200 39800 9294
rect 39834 9434 39838 9492
rect 40986 10602 41032 11372
rect 40986 10586 41034 10602
rect 40986 10294 41000 10586
rect 40986 10278 41034 10294
rect 42054 10586 42100 11388
rect 42054 10294 42058 10586
rect 42092 10294 42100 10586
rect 40986 9508 41032 10278
rect 40986 9492 41034 9508
rect 40986 9434 41000 9492
rect 39834 9258 39858 9294
rect 39834 9200 39908 9258
rect 39776 9090 39908 9200
rect 40948 9200 41000 9390
rect 42054 9492 42100 10294
rect 42054 9412 42058 9492
rect 41034 9200 41074 9390
rect 35548 9000 39998 9090
rect 35560 8994 39998 9000
rect 37674 8972 37756 8994
rect 36618 8238 36686 8254
rect 38742 8238 38810 8270
rect 34466 8228 38810 8238
rect 34376 8184 38810 8228
rect 34376 8148 38818 8184
rect 34376 8138 38666 8148
rect 34466 7960 34592 8138
rect 34466 7958 34528 7960
rect 32284 7662 32290 7862
rect 33258 7818 33308 7954
rect 32244 6860 32290 7662
rect 32244 6568 32250 6860
rect 32284 6568 32290 6860
rect 32244 5766 32290 6568
rect 32244 5474 32250 5766
rect 32284 5474 32290 5766
rect 32244 4672 32290 5474
rect 32244 4380 32250 4672
rect 32284 4380 32290 4672
rect 32244 3578 32290 4380
rect 32244 3548 32250 3578
rect 31226 3286 31264 3358
rect 31182 3176 31264 3286
rect 32284 3548 32290 3578
rect 33300 7662 33308 7818
rect 33342 7818 33384 7954
rect 33342 7662 33346 7818
rect 33300 6860 33346 7662
rect 33300 6568 33308 6860
rect 33342 6568 33346 6860
rect 33300 5766 33346 6568
rect 34514 7668 34528 7958
rect 34562 7958 34592 7960
rect 35586 7960 35620 7976
rect 34562 7858 34582 7958
rect 34514 7652 34562 7668
rect 35582 7668 35586 7866
rect 36618 7960 36686 8138
rect 36618 7872 36644 7960
rect 35620 7668 35628 7866
rect 34514 6882 34560 7652
rect 34514 6866 34562 6882
rect 34514 6574 34528 6866
rect 34514 6558 34562 6574
rect 35582 6866 35628 7668
rect 35582 6574 35586 6866
rect 35620 6574 35628 6866
rect 33300 5474 33308 5766
rect 33342 5474 33346 5766
rect 33300 4672 33346 5474
rect 33874 6426 34024 6552
rect 33874 5230 33896 6426
rect 33990 5230 34024 6426
rect 33874 4906 34024 5230
rect 34514 5788 34560 6558
rect 34514 5772 34562 5788
rect 34514 5480 34528 5772
rect 34514 5464 34562 5480
rect 35582 5772 35628 6574
rect 35582 5480 35586 5772
rect 35620 5480 35628 5772
rect 33300 4380 33308 4672
rect 33342 4380 33346 4672
rect 33300 3578 33346 4380
rect 33300 3520 33308 3578
rect 32250 3270 32284 3286
rect 33284 3286 33308 3380
rect 33342 3520 33346 3578
rect 34514 4694 34560 5464
rect 34514 4678 34562 4694
rect 34514 4386 34528 4678
rect 34514 4370 34562 4386
rect 35582 4678 35628 5480
rect 35582 4386 35586 4678
rect 35620 4386 35628 4678
rect 34514 3600 34560 4370
rect 34514 3584 34562 3600
rect 34514 3526 34528 3584
rect 33342 3286 33366 3380
rect 33284 3228 33366 3286
rect 35582 3584 35628 4386
rect 35582 3504 35586 3584
rect 34528 3276 34562 3292
rect 35566 3292 35586 3392
rect 35620 3504 35628 3584
rect 36634 7668 36644 7872
rect 36678 7924 36686 7960
rect 37702 7960 37736 7976
rect 36678 7872 36692 7924
rect 36678 7668 36680 7872
rect 36634 6866 36680 7668
rect 36634 6574 36644 6866
rect 36678 6574 36680 6866
rect 36634 5772 36680 6574
rect 36634 5480 36644 5772
rect 36678 5480 36680 5772
rect 36634 4678 36680 5480
rect 36634 4386 36644 4678
rect 36678 4386 36680 4678
rect 36634 3584 36680 4386
rect 36634 3526 36644 3584
rect 35620 3292 35648 3392
rect 35566 3228 35648 3292
rect 36678 3526 36680 3584
rect 38734 7960 38818 8148
rect 37736 7668 37748 7872
rect 38734 7868 38760 7960
rect 37702 6866 37748 7668
rect 37736 6574 37748 6866
rect 37702 5772 37748 6574
rect 37736 5480 37748 5772
rect 37702 4678 37748 5480
rect 37736 4386 37748 4678
rect 37702 3584 37748 4386
rect 36644 3276 36678 3292
rect 37692 3292 37702 3364
rect 37736 3510 37748 3584
rect 38754 7668 38760 7868
rect 38794 7868 38818 7960
rect 39782 7960 39908 8994
rect 40948 8238 41074 9200
rect 42038 9200 42058 9300
rect 42092 9412 42100 9492
rect 43106 13576 43116 13780
rect 43150 13832 43158 13868
rect 44174 13868 44208 13884
rect 43150 13780 43164 13832
rect 43150 13576 43152 13780
rect 43106 12774 43152 13576
rect 43106 12482 43116 12774
rect 43150 12482 43152 12774
rect 43106 11680 43152 12482
rect 43106 11388 43116 11680
rect 43150 11388 43152 11680
rect 43106 10586 43152 11388
rect 43106 10294 43116 10586
rect 43150 10294 43152 10586
rect 43106 9492 43152 10294
rect 43106 9434 43116 9492
rect 42092 9200 42120 9300
rect 42038 9090 42120 9200
rect 43150 9434 43152 9492
rect 45206 13868 45290 14056
rect 44208 13576 44220 13780
rect 45206 13776 45232 13868
rect 44174 12774 44220 13576
rect 44208 12482 44220 12774
rect 44174 11680 44220 12482
rect 44208 11388 44220 11680
rect 44174 10586 44220 11388
rect 44208 10294 44220 10586
rect 44174 9492 44220 10294
rect 43116 9184 43150 9200
rect 44164 9200 44174 9272
rect 44208 9418 44220 9492
rect 45226 13576 45232 13776
rect 45266 13776 45290 13868
rect 46256 13868 46382 14850
rect 47528 14168 47654 15078
rect 48616 15078 48636 15178
rect 48670 15290 48678 15370
rect 49684 19454 49694 19658
rect 49728 19710 49736 19746
rect 50752 19746 50786 19762
rect 49728 19658 49742 19710
rect 49728 19454 49730 19658
rect 49684 18652 49730 19454
rect 49684 18360 49694 18652
rect 49728 18360 49730 18652
rect 49684 17558 49730 18360
rect 49684 17266 49694 17558
rect 49728 17266 49730 17558
rect 49684 16464 49730 17266
rect 49684 16172 49694 16464
rect 49728 16172 49730 16464
rect 49684 15370 49730 16172
rect 49684 15312 49694 15370
rect 48670 15078 48698 15178
rect 48616 14968 48698 15078
rect 49728 15312 49730 15370
rect 51784 19746 51868 19934
rect 50786 19454 50798 19658
rect 51784 19654 51810 19746
rect 50752 18652 50798 19454
rect 50786 18360 50798 18652
rect 50752 17558 50798 18360
rect 50786 17266 50798 17558
rect 50752 16464 50798 17266
rect 50786 16172 50798 16464
rect 50752 15370 50798 16172
rect 49694 15062 49728 15078
rect 50742 15078 50752 15150
rect 50786 15296 50798 15370
rect 51804 19454 51810 19654
rect 51844 19654 51868 19746
rect 52858 19746 52954 20736
rect 54024 20038 54150 20956
rect 55130 20956 55150 21056
rect 55184 21168 55192 21248
rect 56198 25332 56208 25536
rect 56242 25588 56250 25624
rect 57266 25624 57300 25640
rect 56242 25536 56256 25588
rect 56242 25332 56244 25536
rect 56198 24530 56244 25332
rect 56198 24238 56208 24530
rect 56242 24238 56244 24530
rect 56198 23436 56244 24238
rect 56198 23144 56208 23436
rect 56242 23144 56244 23436
rect 56198 22342 56244 23144
rect 56198 22050 56208 22342
rect 56242 22050 56244 22342
rect 56198 21248 56244 22050
rect 56198 21190 56208 21248
rect 55184 20956 55212 21056
rect 55130 20846 55212 20956
rect 56242 21190 56244 21248
rect 58298 25624 58382 25812
rect 57300 25332 57312 25536
rect 58298 25532 58324 25624
rect 57266 24530 57312 25332
rect 57300 24238 57312 24530
rect 57266 23436 57312 24238
rect 57300 23144 57312 23436
rect 57266 22342 57312 23144
rect 57300 22050 57312 22342
rect 57266 21248 57312 22050
rect 56208 20940 56242 20956
rect 57256 20956 57266 21028
rect 57300 21174 57312 21248
rect 58318 25332 58324 25532
rect 58358 25532 58382 25624
rect 59356 25624 59452 26586
rect 67546 26320 68312 26348
rect 67546 26188 67586 26320
rect 68284 26188 68312 26320
rect 67546 26160 68312 26188
rect 93948 26288 94478 26316
rect 66326 25864 66394 25878
rect 67860 25864 68078 26160
rect 93948 26156 93994 26288
rect 94426 26156 94478 26288
rect 93948 26134 94478 26156
rect 62098 25846 62166 25856
rect 64202 25846 64270 25862
rect 66306 25846 68924 25864
rect 62098 25844 68924 25846
rect 70664 25844 70732 25860
rect 72788 25844 72856 25876
rect 62098 25836 72856 25844
rect 79482 25836 79550 25850
rect 61960 25828 72856 25836
rect 73852 25828 73926 25834
rect 61960 25756 73926 25828
rect 75254 25818 75322 25828
rect 77358 25818 77426 25834
rect 79462 25818 82080 25836
rect 75254 25816 82080 25818
rect 83820 25816 83888 25832
rect 85944 25816 86012 25848
rect 92716 25828 92784 25842
rect 94142 25828 94370 26134
rect 99178 25838 99246 25840
rect 75254 25808 86012 25816
rect 61960 25746 66250 25756
rect 66306 25754 73926 25756
rect 59356 25546 59382 25624
rect 58358 25332 58364 25532
rect 58318 24530 58364 25332
rect 58318 24238 58324 24530
rect 58358 24238 58364 24530
rect 58318 23436 58364 24238
rect 58318 23144 58324 23436
rect 58358 23144 58364 23436
rect 58318 22342 58364 23144
rect 58318 22050 58324 22342
rect 58358 22050 58364 22342
rect 58318 21248 58364 22050
rect 58318 21218 58324 21248
rect 57300 20956 57338 21028
rect 57256 20846 57338 20956
rect 58358 21218 58364 21248
rect 59374 25332 59382 25546
rect 59416 25546 59452 25624
rect 62098 25568 62166 25746
rect 59416 25332 59420 25546
rect 59374 24530 59420 25332
rect 59374 24238 59382 24530
rect 59416 24238 59420 24530
rect 62098 25276 62112 25568
rect 62146 25466 62166 25568
rect 63170 25568 63204 25584
rect 62098 25260 62146 25276
rect 63166 25276 63170 25474
rect 64202 25568 64270 25746
rect 66306 25744 72712 25754
rect 66306 25710 68924 25744
rect 64202 25480 64228 25568
rect 63204 25276 63212 25474
rect 59374 23436 59420 24238
rect 59374 23144 59382 23436
rect 59416 23144 59420 23436
rect 59374 22342 59420 23144
rect 59572 24250 59934 24514
rect 59572 22696 59614 24250
rect 59864 22696 59934 24250
rect 62098 24490 62144 25260
rect 62098 24474 62146 24490
rect 62098 24182 62112 24474
rect 62098 24166 62146 24182
rect 63166 24474 63212 25276
rect 63166 24182 63170 24474
rect 63204 24182 63212 24474
rect 59572 22418 59934 22696
rect 61458 24034 61608 24160
rect 61458 22838 61480 24034
rect 61574 22838 61608 24034
rect 61458 22514 61608 22838
rect 62098 23396 62144 24166
rect 62098 23380 62146 23396
rect 62098 23088 62112 23380
rect 62098 23072 62146 23088
rect 63166 23380 63212 24182
rect 63166 23088 63170 23380
rect 63204 23088 63212 23380
rect 59374 22050 59382 22342
rect 59416 22050 59420 22342
rect 59374 21248 59420 22050
rect 59374 21190 59382 21248
rect 58324 20940 58358 20956
rect 59358 20956 59382 21050
rect 59416 21190 59420 21248
rect 62098 22302 62144 23072
rect 62098 22286 62146 22302
rect 62098 21994 62112 22286
rect 62098 21978 62146 21994
rect 63166 22286 63212 23088
rect 63166 21994 63170 22286
rect 63204 21994 63212 22286
rect 62098 21208 62144 21978
rect 62098 21192 62146 21208
rect 62098 21134 62112 21192
rect 59416 21014 59440 21050
rect 59416 20956 59460 21014
rect 59358 20846 59460 20956
rect 63166 21192 63212 21994
rect 63166 21112 63170 21192
rect 62112 20884 62146 20900
rect 63150 20900 63170 21000
rect 63204 21112 63212 21192
rect 64218 25276 64228 25480
rect 64262 25532 64270 25568
rect 65286 25568 65320 25584
rect 64262 25480 64276 25532
rect 64262 25276 64264 25480
rect 64218 24474 64264 25276
rect 64218 24182 64228 24474
rect 64262 24182 64264 24474
rect 64218 23380 64264 24182
rect 64218 23088 64228 23380
rect 64262 23088 64264 23380
rect 64218 22286 64264 23088
rect 64218 21994 64228 22286
rect 64262 21994 64264 22286
rect 64218 21192 64264 21994
rect 64218 21134 64228 21192
rect 63204 20900 63232 21000
rect 55130 20756 59580 20846
rect 55142 20750 59580 20756
rect 63150 20790 63232 20900
rect 64262 21134 64264 21192
rect 66318 25568 66402 25710
rect 67860 25702 68078 25710
rect 65320 25276 65332 25480
rect 66318 25476 66344 25568
rect 65286 24474 65332 25276
rect 65320 24182 65332 24474
rect 65286 23380 65332 24182
rect 65320 23088 65332 23380
rect 65286 22286 65332 23088
rect 65320 21994 65332 22286
rect 65286 21192 65332 21994
rect 64228 20884 64262 20900
rect 65276 20900 65286 20972
rect 65320 21118 65332 21192
rect 66338 25276 66344 25476
rect 66378 25476 66402 25568
rect 67402 25568 67436 25584
rect 66378 25276 66384 25476
rect 66338 24474 66384 25276
rect 66338 24182 66344 24474
rect 66378 24182 66384 24474
rect 66338 23380 66384 24182
rect 66338 23088 66344 23380
rect 66378 23088 66384 23380
rect 66338 22286 66384 23088
rect 66338 21994 66344 22286
rect 66378 21994 66384 22286
rect 66338 21192 66384 21994
rect 66338 21162 66344 21192
rect 65320 20900 65358 20972
rect 65276 20790 65358 20900
rect 66378 21162 66384 21192
rect 67394 25276 67402 25496
rect 68560 25566 68628 25710
rect 67436 25276 67440 25496
rect 67394 24474 67440 25276
rect 67394 24182 67402 24474
rect 67436 24182 67440 24474
rect 67394 23380 67440 24182
rect 68560 25274 68574 25566
rect 68608 25464 68628 25566
rect 69632 25566 69666 25582
rect 68560 25258 68608 25274
rect 69628 25274 69632 25472
rect 70664 25566 70732 25744
rect 72780 25726 73926 25754
rect 70664 25478 70690 25566
rect 69666 25274 69674 25472
rect 68560 24488 68606 25258
rect 68560 24472 68608 24488
rect 68560 24180 68574 24472
rect 68560 24164 68608 24180
rect 69628 24472 69674 25274
rect 69628 24180 69632 24472
rect 69666 24180 69674 24472
rect 67394 23088 67402 23380
rect 67436 23088 67440 23380
rect 67394 22286 67440 23088
rect 67920 24032 68070 24158
rect 67920 22836 67942 24032
rect 68036 22836 68070 24032
rect 67920 22512 68070 22836
rect 68560 23394 68606 24164
rect 68560 23378 68608 23394
rect 68560 23086 68574 23378
rect 68560 23070 68608 23086
rect 69628 23378 69674 24180
rect 69628 23086 69632 23378
rect 69666 23086 69674 23378
rect 67394 21994 67402 22286
rect 67436 21994 67440 22286
rect 67394 21192 67440 21994
rect 67394 21134 67402 21192
rect 66344 20884 66378 20900
rect 67378 20900 67402 20994
rect 67436 21134 67440 21192
rect 68560 22300 68606 23070
rect 68560 22284 68608 22300
rect 68560 21992 68574 22284
rect 68560 21976 68608 21992
rect 69628 22284 69674 23086
rect 69628 21992 69632 22284
rect 69666 21992 69674 22284
rect 68560 21206 68606 21976
rect 68560 21190 68608 21206
rect 68560 21132 68574 21190
rect 67436 20900 67460 20994
rect 67378 20790 67460 20900
rect 69628 21190 69674 21992
rect 69628 21110 69632 21190
rect 68574 20882 68608 20898
rect 69612 20898 69632 20998
rect 69666 21110 69674 21190
rect 70680 25274 70690 25478
rect 70724 25530 70732 25566
rect 71748 25566 71782 25582
rect 70724 25478 70738 25530
rect 70724 25274 70726 25478
rect 70680 24472 70726 25274
rect 70680 24180 70690 24472
rect 70724 24180 70726 24472
rect 70680 23378 70726 24180
rect 70680 23086 70690 23378
rect 70724 23086 70726 23378
rect 70680 22284 70726 23086
rect 70680 21992 70690 22284
rect 70724 21992 70726 22284
rect 70680 21190 70726 21992
rect 70680 21132 70690 21190
rect 69666 20898 69694 20998
rect 57256 20728 57338 20750
rect 56182 20038 56250 20054
rect 58306 20038 58374 20070
rect 54024 20028 58374 20038
rect 53940 19984 58374 20028
rect 53940 19948 58382 19984
rect 53940 19938 58230 19948
rect 51844 19454 51850 19654
rect 52858 19632 52868 19746
rect 51804 18652 51850 19454
rect 51804 18360 51810 18652
rect 51844 18360 51850 18652
rect 51804 17558 51850 18360
rect 51804 17266 51810 17558
rect 51844 17266 51850 17558
rect 51804 16464 51850 17266
rect 51804 16172 51810 16464
rect 51844 16172 51850 16464
rect 51804 15370 51850 16172
rect 51804 15340 51810 15370
rect 50786 15078 50824 15150
rect 50742 14968 50824 15078
rect 51844 15340 51850 15370
rect 52860 19454 52868 19632
rect 52902 19632 52954 19746
rect 54024 19760 54150 19938
rect 54024 19686 54092 19760
rect 52902 19454 52906 19632
rect 52860 18652 52906 19454
rect 52860 18360 52868 18652
rect 52902 18360 52906 18652
rect 52860 17558 52906 18360
rect 54078 19468 54092 19686
rect 54126 19686 54150 19760
rect 55150 19760 55184 19776
rect 54126 19658 54146 19686
rect 54078 19452 54126 19468
rect 55146 19468 55150 19666
rect 56182 19760 56250 19938
rect 56182 19672 56208 19760
rect 55184 19468 55192 19666
rect 54078 18682 54124 19452
rect 54078 18666 54126 18682
rect 54078 18374 54092 18666
rect 54078 18358 54126 18374
rect 55146 18666 55192 19468
rect 55146 18374 55150 18666
rect 55184 18374 55192 18666
rect 52860 17266 52868 17558
rect 52902 17266 52906 17558
rect 52860 16464 52906 17266
rect 53438 18226 53588 18352
rect 53438 17030 53460 18226
rect 53554 17030 53588 18226
rect 53438 16706 53588 17030
rect 54078 17588 54124 18358
rect 54078 17572 54126 17588
rect 54078 17280 54092 17572
rect 54078 17264 54126 17280
rect 55146 17572 55192 18374
rect 55146 17280 55150 17572
rect 55184 17280 55192 17572
rect 52860 16172 52868 16464
rect 52902 16172 52906 16464
rect 52860 15370 52906 16172
rect 52860 15332 52868 15370
rect 51810 15062 51844 15078
rect 52830 15078 52868 15332
rect 52902 15332 52906 15370
rect 54078 16494 54124 17264
rect 54078 16478 54126 16494
rect 54078 16186 54092 16478
rect 54078 16170 54126 16186
rect 55146 16478 55192 17280
rect 55146 16186 55150 16478
rect 55184 16186 55192 16478
rect 54078 15400 54124 16170
rect 54078 15384 54126 15400
rect 54078 15360 54092 15384
rect 52902 15078 52956 15332
rect 52830 14968 52956 15078
rect 54038 15092 54092 15360
rect 55146 15384 55192 16186
rect 54126 15092 54164 15360
rect 55146 15304 55150 15384
rect 48616 14878 53066 14968
rect 48628 14872 53066 14878
rect 50742 14850 50824 14872
rect 49678 14168 49746 14184
rect 51802 14168 51870 14200
rect 47528 14158 51870 14168
rect 47436 14114 51870 14158
rect 47436 14078 51878 14114
rect 47436 14068 51726 14078
rect 47528 13892 47654 14068
rect 45266 13576 45272 13776
rect 46256 13648 46290 13868
rect 45226 12774 45272 13576
rect 45226 12482 45232 12774
rect 45266 12482 45272 12774
rect 45226 11680 45272 12482
rect 45226 11388 45232 11680
rect 45266 11388 45272 11680
rect 45226 10586 45272 11388
rect 45226 10294 45232 10586
rect 45266 10294 45272 10586
rect 45226 9492 45272 10294
rect 45226 9462 45232 9492
rect 44208 9200 44246 9272
rect 44164 9090 44246 9200
rect 45266 9462 45272 9492
rect 46282 13576 46290 13648
rect 46324 13648 46382 13868
rect 47574 13890 47642 13892
rect 46324 13576 46328 13648
rect 46282 12774 46328 13576
rect 46282 12482 46290 12774
rect 46324 12482 46328 12774
rect 47574 13598 47588 13890
rect 47622 13788 47642 13890
rect 48646 13890 48680 13906
rect 47574 13582 47622 13598
rect 48642 13598 48646 13796
rect 49678 13890 49746 14068
rect 49678 13802 49704 13890
rect 48680 13598 48688 13796
rect 47574 12812 47620 13582
rect 47574 12796 47622 12812
rect 47574 12504 47588 12796
rect 47574 12488 47622 12504
rect 48642 12796 48688 13598
rect 48642 12504 48646 12796
rect 48680 12504 48688 12796
rect 46282 11680 46328 12482
rect 46282 11388 46290 11680
rect 46324 11388 46328 11680
rect 46282 10586 46328 11388
rect 46934 12356 47084 12482
rect 46934 11160 46956 12356
rect 47050 11160 47084 12356
rect 46934 10836 47084 11160
rect 47574 11718 47620 12488
rect 47574 11702 47622 11718
rect 47574 11410 47588 11702
rect 47574 11394 47622 11410
rect 48642 11702 48688 12504
rect 48642 11410 48646 11702
rect 48680 11410 48688 11702
rect 46282 10294 46290 10586
rect 46324 10294 46328 10586
rect 46282 9492 46328 10294
rect 46282 9434 46290 9492
rect 45232 9184 45266 9200
rect 46266 9200 46290 9294
rect 46324 9434 46328 9492
rect 47574 10624 47620 11394
rect 47574 10608 47622 10624
rect 47574 10316 47588 10608
rect 47574 10300 47622 10316
rect 48642 10608 48688 11410
rect 48642 10316 48646 10608
rect 48680 10316 48688 10608
rect 47574 9530 47620 10300
rect 47574 9514 47622 9530
rect 47574 9456 47588 9514
rect 46324 9200 46348 9294
rect 46266 9110 46348 9200
rect 47542 9222 47588 9398
rect 48642 9514 48688 10316
rect 48642 9434 48646 9514
rect 47622 9222 47668 9398
rect 46256 9090 46382 9110
rect 42038 9000 46488 9090
rect 42050 8994 46488 9000
rect 44164 8972 44246 8994
rect 43108 8238 43176 8254
rect 45232 8238 45300 8270
rect 40948 8228 45300 8238
rect 40866 8184 45300 8228
rect 40866 8148 45308 8184
rect 40866 8138 45156 8148
rect 40948 8006 41074 8138
rect 39782 7874 39818 7960
rect 38794 7668 38800 7868
rect 38754 6866 38800 7668
rect 38754 6574 38760 6866
rect 38794 6574 38800 6866
rect 38754 5772 38800 6574
rect 38754 5480 38760 5772
rect 38794 5480 38800 5772
rect 38754 4678 38800 5480
rect 38754 4386 38760 4678
rect 38794 4386 38800 4678
rect 38754 3584 38800 4386
rect 38754 3554 38760 3584
rect 37736 3292 37774 3364
rect 33026 3182 36022 3228
rect 37692 3182 37774 3292
rect 38794 3554 38800 3584
rect 39810 7668 39818 7874
rect 39852 7874 39908 7960
rect 41004 7960 41072 8006
rect 39852 7668 39856 7874
rect 39810 6866 39856 7668
rect 39810 6574 39818 6866
rect 39852 6574 39856 6866
rect 39810 5772 39856 6574
rect 41004 7668 41018 7960
rect 41052 7858 41072 7960
rect 42076 7960 42110 7976
rect 41004 7652 41052 7668
rect 42072 7668 42076 7866
rect 43108 7960 43176 8138
rect 43108 7872 43134 7960
rect 42110 7668 42118 7866
rect 41004 6882 41050 7652
rect 41004 6866 41052 6882
rect 41004 6574 41018 6866
rect 41004 6558 41052 6574
rect 42072 6866 42118 7668
rect 42072 6574 42076 6866
rect 42110 6574 42118 6866
rect 40364 6426 40514 6552
rect 40364 5796 40386 6426
rect 39810 5480 39818 5772
rect 39852 5480 39856 5772
rect 39810 4678 39856 5480
rect 39810 4386 39818 4678
rect 39852 4386 39856 4678
rect 39810 3584 39856 4386
rect 39810 3526 39818 3584
rect 38760 3276 38794 3292
rect 39794 3292 39818 3386
rect 39852 3526 39856 3584
rect 40322 5230 40386 5796
rect 40480 5796 40514 6426
rect 40480 5230 40566 5796
rect 39852 3292 39876 3386
rect 39794 3182 39876 3292
rect 33026 3176 40016 3182
rect 29056 3164 40016 3176
rect 26502 3160 40016 3164
rect 22534 3086 40016 3160
rect 22534 3080 36022 3086
rect 9550 3072 13988 3078
rect 3036 3064 7474 3070
rect 5150 3042 5232 3064
rect 11664 3050 11746 3072
rect 18170 3058 18252 3080
rect 22534 3070 29524 3080
rect 22546 3064 29524 3070
rect 24660 3042 24742 3064
rect 26502 2960 29524 3064
rect 31182 3058 31264 3080
rect 33026 2970 36022 3080
rect 37692 3064 37774 3086
rect 40322 -496 40566 5230
rect 41004 5788 41050 6558
rect 41004 5772 41052 5788
rect 41004 5480 41018 5772
rect 41004 5464 41052 5480
rect 42072 5772 42118 6574
rect 42072 5480 42076 5772
rect 42110 5480 42118 5772
rect 41004 4694 41050 5464
rect 41004 4678 41052 4694
rect 41004 4386 41018 4678
rect 41004 4370 41052 4386
rect 42072 4678 42118 5480
rect 42072 4386 42076 4678
rect 42110 4386 42118 4678
rect 41004 3600 41050 4370
rect 41004 3584 41052 3600
rect 41004 3526 41018 3584
rect 42072 3584 42118 4386
rect 42072 3504 42076 3584
rect 41018 3276 41052 3292
rect 42056 3292 42076 3392
rect 42110 3504 42118 3584
rect 43124 7668 43134 7872
rect 43168 7924 43176 7960
rect 44192 7960 44226 7976
rect 43168 7872 43182 7924
rect 43168 7668 43170 7872
rect 43124 6866 43170 7668
rect 43124 6574 43134 6866
rect 43168 6574 43170 6866
rect 43124 5772 43170 6574
rect 43124 5480 43134 5772
rect 43168 5480 43170 5772
rect 43124 4678 43170 5480
rect 43124 4386 43134 4678
rect 43168 4386 43170 4678
rect 43124 3584 43170 4386
rect 43124 3526 43134 3584
rect 42110 3292 42138 3392
rect 42056 3182 42138 3292
rect 43168 3526 43170 3584
rect 45224 7960 45308 8148
rect 44226 7668 44238 7872
rect 45224 7868 45250 7960
rect 44192 6866 44238 7668
rect 44226 6574 44238 6866
rect 44192 5772 44238 6574
rect 44226 5480 44238 5772
rect 44192 4678 44238 5480
rect 44226 4386 44238 4678
rect 44192 3584 44238 4386
rect 43134 3276 43168 3292
rect 44182 3292 44192 3364
rect 44226 3510 44238 3584
rect 45244 7668 45250 7868
rect 45284 7868 45308 7960
rect 46256 7960 46382 8994
rect 47542 8260 47668 9222
rect 48626 9222 48646 9322
rect 48680 9434 48688 9514
rect 49694 13598 49704 13802
rect 49738 13854 49746 13890
rect 50762 13890 50796 13906
rect 49738 13802 49752 13854
rect 49738 13598 49740 13802
rect 49694 12796 49740 13598
rect 49694 12504 49704 12796
rect 49738 12504 49740 12796
rect 49694 11702 49740 12504
rect 49694 11410 49704 11702
rect 49738 11410 49740 11702
rect 49694 10608 49740 11410
rect 49694 10316 49704 10608
rect 49738 10316 49740 10608
rect 49694 9514 49740 10316
rect 49694 9456 49704 9514
rect 48680 9222 48708 9322
rect 48626 9112 48708 9222
rect 49738 9456 49740 9514
rect 51794 13890 51878 14078
rect 52830 13948 52956 14872
rect 54038 14182 54164 15092
rect 55130 15092 55150 15192
rect 55184 15304 55192 15384
rect 56198 19468 56208 19672
rect 56242 19724 56250 19760
rect 57266 19760 57300 19776
rect 56242 19672 56256 19724
rect 56242 19468 56244 19672
rect 56198 18666 56244 19468
rect 56198 18374 56208 18666
rect 56242 18374 56244 18666
rect 56198 17572 56244 18374
rect 56198 17280 56208 17572
rect 56242 17280 56244 17572
rect 56198 16478 56244 17280
rect 56198 16186 56208 16478
rect 56242 16186 56244 16478
rect 56198 15384 56244 16186
rect 56198 15326 56208 15384
rect 55184 15092 55212 15192
rect 55130 14982 55212 15092
rect 56242 15326 56244 15384
rect 58298 19760 58382 19948
rect 57300 19468 57312 19672
rect 58298 19668 58324 19760
rect 57266 18666 57312 19468
rect 57300 18374 57312 18666
rect 57266 17572 57312 18374
rect 57300 17280 57312 17572
rect 57266 16478 57312 17280
rect 57300 16186 57312 16478
rect 57266 15384 57312 16186
rect 56208 15076 56242 15092
rect 57256 15092 57266 15164
rect 57300 15310 57312 15384
rect 58318 19468 58324 19668
rect 58358 19668 58382 19760
rect 59364 19760 59460 20750
rect 63150 20700 67600 20790
rect 63162 20694 67600 20700
rect 69612 20788 69694 20898
rect 70724 21132 70726 21190
rect 72780 25566 72864 25726
rect 71782 25274 71794 25478
rect 72780 25474 72806 25566
rect 71748 24472 71794 25274
rect 71782 24180 71794 24472
rect 71748 23378 71794 24180
rect 71782 23086 71794 23378
rect 71748 22284 71794 23086
rect 71782 21992 71794 22284
rect 71748 21190 71794 21992
rect 70690 20882 70724 20898
rect 71738 20898 71748 20970
rect 71782 21116 71794 21190
rect 72800 25274 72806 25474
rect 72840 25474 72864 25566
rect 73852 25566 73926 25726
rect 75116 25762 86012 25808
rect 88488 25810 88556 25820
rect 90592 25810 90660 25826
rect 92696 25810 95314 25828
rect 99138 25826 100334 25838
rect 88488 25808 95314 25810
rect 97054 25808 97122 25824
rect 99138 25808 100356 25826
rect 88488 25800 100356 25808
rect 75116 25728 86020 25762
rect 75116 25718 79406 25728
rect 79462 25726 86020 25728
rect 72840 25274 72846 25474
rect 73852 25452 73864 25566
rect 72800 24472 72846 25274
rect 72800 24180 72806 24472
rect 72840 24180 72846 24472
rect 72800 23378 72846 24180
rect 72800 23086 72806 23378
rect 72840 23086 72846 23378
rect 72800 22284 72846 23086
rect 72800 21992 72806 22284
rect 72840 21992 72846 22284
rect 72800 21190 72846 21992
rect 72800 21160 72806 21190
rect 71782 20898 71820 20970
rect 71738 20788 71820 20898
rect 72840 21160 72846 21190
rect 73856 25274 73864 25452
rect 73898 25452 73926 25566
rect 75254 25540 75322 25718
rect 73898 25274 73902 25452
rect 73856 24472 73902 25274
rect 73856 24180 73864 24472
rect 73898 24180 73902 24472
rect 73856 23378 73902 24180
rect 75254 25248 75268 25540
rect 75302 25438 75322 25540
rect 76326 25540 76360 25556
rect 75254 25232 75302 25248
rect 76322 25248 76326 25446
rect 77358 25540 77426 25718
rect 79462 25716 85868 25726
rect 79462 25682 82080 25716
rect 77358 25452 77384 25540
rect 76360 25248 76368 25446
rect 75254 24462 75300 25232
rect 75254 24446 75302 24462
rect 75254 24154 75268 24446
rect 75254 24138 75302 24154
rect 76322 24446 76368 25248
rect 76322 24154 76326 24446
rect 76360 24154 76368 24446
rect 73856 23086 73864 23378
rect 73898 23086 73902 23378
rect 73856 22284 73902 23086
rect 74614 24006 74764 24132
rect 74614 22810 74636 24006
rect 74730 22810 74764 24006
rect 74614 22486 74764 22810
rect 75254 23368 75300 24138
rect 75254 23352 75302 23368
rect 75254 23060 75268 23352
rect 75254 23044 75302 23060
rect 76322 23352 76368 24154
rect 76322 23060 76326 23352
rect 76360 23060 76368 23352
rect 73856 21992 73864 22284
rect 73898 21992 73902 22284
rect 73856 21190 73902 21992
rect 73856 21132 73864 21190
rect 72806 20882 72840 20898
rect 73840 20898 73864 20992
rect 73898 21132 73902 21190
rect 75254 22274 75300 23044
rect 75254 22258 75302 22274
rect 75254 21966 75268 22258
rect 75254 21950 75302 21966
rect 76322 22258 76368 23060
rect 76322 21966 76326 22258
rect 76360 21966 76368 22258
rect 75254 21180 75300 21950
rect 75254 21164 75302 21180
rect 75254 21106 75268 21164
rect 73898 20898 73922 20992
rect 73840 20788 73922 20898
rect 76322 21164 76368 21966
rect 76322 21084 76326 21164
rect 75268 20856 75302 20872
rect 76306 20872 76326 20972
rect 76360 21084 76368 21164
rect 77374 25248 77384 25452
rect 77418 25504 77426 25540
rect 78442 25540 78476 25556
rect 77418 25452 77432 25504
rect 77418 25248 77420 25452
rect 77374 24446 77420 25248
rect 77374 24154 77384 24446
rect 77418 24154 77420 24446
rect 77374 23352 77420 24154
rect 77374 23060 77384 23352
rect 77418 23060 77420 23352
rect 77374 22258 77420 23060
rect 77374 21966 77384 22258
rect 77418 21966 77420 22258
rect 77374 21164 77420 21966
rect 77374 21106 77384 21164
rect 76360 20872 76388 20972
rect 69612 20698 74062 20788
rect 65276 20672 65358 20694
rect 69624 20692 74062 20698
rect 76306 20762 76388 20872
rect 77418 21106 77420 21164
rect 79474 25540 79558 25682
rect 78476 25248 78488 25452
rect 79474 25448 79500 25540
rect 78442 24446 78488 25248
rect 78476 24154 78488 24446
rect 78442 23352 78488 24154
rect 78476 23060 78488 23352
rect 78442 22258 78488 23060
rect 78476 21966 78488 22258
rect 78442 21164 78488 21966
rect 77384 20856 77418 20872
rect 78432 20872 78442 20944
rect 78476 21090 78488 21164
rect 79494 25248 79500 25448
rect 79534 25448 79558 25540
rect 80558 25540 80592 25556
rect 79534 25248 79540 25448
rect 79494 24446 79540 25248
rect 79494 24154 79500 24446
rect 79534 24154 79540 24446
rect 79494 23352 79540 24154
rect 79494 23060 79500 23352
rect 79534 23060 79540 23352
rect 79494 22258 79540 23060
rect 79494 21966 79500 22258
rect 79534 21966 79540 22258
rect 79494 21164 79540 21966
rect 79494 21134 79500 21164
rect 78476 20872 78514 20944
rect 78432 20762 78514 20872
rect 79534 21134 79540 21164
rect 80550 25248 80558 25468
rect 81716 25538 81784 25682
rect 80592 25248 80596 25468
rect 80550 24446 80596 25248
rect 80550 24154 80558 24446
rect 80592 24154 80596 24446
rect 80550 23352 80596 24154
rect 81716 25246 81730 25538
rect 81764 25436 81784 25538
rect 82788 25538 82822 25554
rect 81716 25230 81764 25246
rect 82784 25246 82788 25444
rect 83820 25538 83888 25716
rect 83820 25450 83846 25538
rect 82822 25246 82830 25444
rect 81716 24460 81762 25230
rect 81716 24444 81764 24460
rect 81716 24152 81730 24444
rect 81716 24136 81764 24152
rect 82784 24444 82830 25246
rect 82784 24152 82788 24444
rect 82822 24152 82830 24444
rect 80550 23060 80558 23352
rect 80592 23060 80596 23352
rect 80550 22258 80596 23060
rect 81076 24004 81226 24130
rect 81076 22808 81098 24004
rect 81192 22808 81226 24004
rect 81076 22484 81226 22808
rect 81716 23366 81762 24136
rect 81716 23350 81764 23366
rect 81716 23058 81730 23350
rect 81716 23042 81764 23058
rect 82784 23350 82830 24152
rect 82784 23058 82788 23350
rect 82822 23058 82830 23350
rect 80550 21966 80558 22258
rect 80592 21966 80596 22258
rect 80550 21164 80596 21966
rect 80550 21106 80558 21164
rect 79500 20856 79534 20872
rect 80534 20872 80558 20966
rect 80592 21106 80596 21164
rect 81716 22272 81762 23042
rect 81716 22256 81764 22272
rect 81716 21964 81730 22256
rect 81716 21948 81764 21964
rect 82784 22256 82830 23058
rect 82784 21964 82788 22256
rect 82822 21964 82830 22256
rect 81716 21178 81762 21948
rect 81716 21162 81764 21178
rect 81716 21104 81730 21162
rect 80592 20872 80616 20966
rect 80534 20762 80616 20872
rect 82784 21162 82830 21964
rect 82784 21082 82788 21162
rect 81730 20854 81764 20870
rect 82768 20870 82788 20970
rect 82822 21082 82830 21162
rect 83836 25246 83846 25450
rect 83880 25502 83888 25538
rect 84904 25538 84938 25554
rect 83880 25450 83894 25502
rect 83880 25246 83882 25450
rect 83836 24444 83882 25246
rect 83836 24152 83846 24444
rect 83880 24152 83882 24444
rect 83836 23350 83882 24152
rect 83836 23058 83846 23350
rect 83880 23058 83882 23350
rect 83836 22256 83882 23058
rect 83836 21964 83846 22256
rect 83880 21964 83882 22256
rect 83836 21162 83882 21964
rect 83836 21104 83846 21162
rect 82822 20870 82850 20970
rect 71738 20670 71820 20692
rect 76306 20672 80756 20762
rect 76318 20666 80756 20672
rect 82768 20760 82850 20870
rect 83880 21104 83882 21162
rect 85936 25538 86020 25726
rect 88350 25720 100356 25800
rect 88350 25710 92640 25720
rect 92696 25718 100356 25720
rect 84938 25246 84950 25450
rect 85936 25446 85962 25538
rect 84904 24444 84950 25246
rect 84938 24152 84950 24444
rect 84904 23350 84950 24152
rect 84938 23058 84950 23350
rect 84904 22256 84950 23058
rect 84938 21964 84950 22256
rect 84904 21162 84950 21964
rect 83846 20854 83880 20870
rect 84894 20870 84904 20942
rect 84938 21088 84950 21162
rect 85956 25246 85962 25446
rect 85996 25446 86020 25538
rect 87020 25538 87054 25554
rect 85996 25246 86002 25446
rect 85956 24444 86002 25246
rect 85956 24152 85962 24444
rect 85996 24152 86002 24444
rect 85956 23350 86002 24152
rect 85956 23058 85962 23350
rect 85996 23058 86002 23350
rect 85956 22256 86002 23058
rect 85956 21964 85962 22256
rect 85996 21964 86002 22256
rect 85956 21162 86002 21964
rect 85956 21132 85962 21162
rect 84938 20870 84976 20942
rect 84894 20760 84976 20870
rect 85996 21132 86002 21162
rect 87012 25246 87020 25466
rect 88488 25532 88556 25710
rect 87054 25246 87058 25466
rect 87012 24444 87058 25246
rect 87012 24152 87020 24444
rect 87054 24152 87058 24444
rect 87012 23350 87058 24152
rect 88488 25240 88502 25532
rect 88536 25430 88556 25532
rect 89560 25532 89594 25548
rect 88488 25224 88536 25240
rect 89556 25240 89560 25438
rect 90592 25532 90660 25710
rect 92696 25708 99102 25718
rect 92696 25674 95314 25708
rect 90592 25444 90618 25532
rect 89594 25240 89602 25438
rect 88488 24454 88534 25224
rect 88488 24438 88536 24454
rect 88488 24146 88502 24438
rect 88488 24130 88536 24146
rect 89556 24438 89602 25240
rect 89556 24146 89560 24438
rect 89594 24146 89602 24438
rect 87012 23058 87020 23350
rect 87054 23058 87058 23350
rect 87012 22256 87058 23058
rect 87848 23998 87998 24124
rect 87848 22802 87870 23998
rect 87964 22802 87998 23998
rect 87848 22478 87998 22802
rect 88488 23360 88534 24130
rect 88488 23344 88536 23360
rect 88488 23052 88502 23344
rect 88488 23036 88536 23052
rect 89556 23344 89602 24146
rect 89556 23052 89560 23344
rect 89594 23052 89602 23344
rect 87012 21964 87020 22256
rect 87054 21964 87058 22256
rect 87012 21162 87058 21964
rect 87012 21104 87020 21162
rect 85962 20854 85996 20870
rect 86996 20870 87020 20964
rect 87054 21104 87058 21162
rect 88488 22266 88534 23036
rect 88488 22250 88536 22266
rect 88488 21958 88502 22250
rect 88488 21942 88536 21958
rect 89556 22250 89602 23052
rect 89556 21958 89560 22250
rect 89594 21958 89602 22250
rect 88488 21172 88534 21942
rect 88488 21156 88536 21172
rect 88488 21098 88502 21156
rect 87054 20870 87078 20964
rect 86996 20760 87078 20870
rect 89556 21156 89602 21958
rect 89556 21076 89560 21156
rect 88502 20848 88536 20864
rect 89540 20864 89560 20964
rect 89594 21076 89602 21156
rect 90608 25240 90618 25444
rect 90652 25496 90660 25532
rect 91676 25532 91710 25548
rect 90652 25444 90666 25496
rect 90652 25240 90654 25444
rect 90608 24438 90654 25240
rect 90608 24146 90618 24438
rect 90652 24146 90654 24438
rect 90608 23344 90654 24146
rect 90608 23052 90618 23344
rect 90652 23052 90654 23344
rect 90608 22250 90654 23052
rect 90608 21958 90618 22250
rect 90652 21958 90654 22250
rect 90608 21156 90654 21958
rect 90608 21098 90618 21156
rect 89594 20864 89622 20964
rect 82768 20670 87218 20760
rect 78432 20644 78514 20666
rect 82780 20664 87218 20670
rect 89540 20754 89622 20864
rect 90652 21098 90654 21156
rect 92708 25532 92792 25674
rect 91710 25240 91722 25444
rect 92708 25440 92734 25532
rect 91676 24438 91722 25240
rect 91710 24146 91722 24438
rect 91676 23344 91722 24146
rect 91710 23052 91722 23344
rect 91676 22250 91722 23052
rect 91710 21958 91722 22250
rect 91676 21156 91722 21958
rect 90618 20848 90652 20864
rect 91666 20864 91676 20936
rect 91710 21082 91722 21156
rect 92728 25240 92734 25440
rect 92768 25440 92792 25532
rect 93792 25532 93826 25548
rect 92768 25240 92774 25440
rect 92728 24438 92774 25240
rect 92728 24146 92734 24438
rect 92768 24146 92774 24438
rect 92728 23344 92774 24146
rect 92728 23052 92734 23344
rect 92768 23052 92774 23344
rect 92728 22250 92774 23052
rect 92728 21958 92734 22250
rect 92768 21958 92774 22250
rect 92728 21156 92774 21958
rect 92728 21126 92734 21156
rect 91710 20864 91748 20936
rect 91666 20754 91748 20864
rect 92768 21126 92774 21156
rect 93784 25240 93792 25460
rect 94950 25530 95018 25674
rect 93826 25240 93830 25460
rect 93784 24438 93830 25240
rect 93784 24146 93792 24438
rect 93826 24146 93830 24438
rect 93784 23344 93830 24146
rect 94950 25238 94964 25530
rect 94998 25428 95018 25530
rect 96022 25530 96056 25546
rect 94950 25222 94998 25238
rect 96018 25238 96022 25436
rect 97054 25530 97122 25708
rect 99138 25678 100356 25718
rect 97054 25442 97080 25530
rect 96056 25238 96064 25436
rect 94950 24452 94996 25222
rect 94950 24436 94998 24452
rect 94950 24144 94964 24436
rect 94950 24128 94998 24144
rect 96018 24436 96064 25238
rect 96018 24144 96022 24436
rect 96056 24144 96064 24436
rect 93784 23052 93792 23344
rect 93826 23052 93830 23344
rect 93784 22250 93830 23052
rect 94310 23996 94460 24122
rect 94310 22800 94332 23996
rect 94426 22800 94460 23996
rect 94310 22476 94460 22800
rect 94950 23358 94996 24128
rect 94950 23342 94998 23358
rect 94950 23050 94964 23342
rect 94950 23034 94998 23050
rect 96018 23342 96064 24144
rect 96018 23050 96022 23342
rect 96056 23050 96064 23342
rect 93784 21958 93792 22250
rect 93826 21958 93830 22250
rect 93784 21156 93830 21958
rect 93784 21098 93792 21156
rect 92734 20848 92768 20864
rect 93768 20864 93792 20958
rect 93826 21098 93830 21156
rect 94950 22264 94996 23034
rect 94950 22248 94998 22264
rect 94950 21956 94964 22248
rect 94950 21940 94998 21956
rect 96018 22248 96064 23050
rect 96018 21956 96022 22248
rect 96056 21956 96064 22248
rect 94950 21170 94996 21940
rect 94950 21154 94998 21170
rect 94950 21096 94964 21154
rect 93826 20864 93850 20958
rect 93768 20754 93850 20864
rect 96018 21154 96064 21956
rect 96018 21074 96022 21154
rect 94964 20846 94998 20862
rect 96002 20862 96022 20962
rect 96056 21074 96064 21154
rect 97070 25238 97080 25442
rect 97114 25494 97122 25530
rect 98138 25530 98172 25546
rect 97114 25442 97128 25494
rect 97114 25238 97116 25442
rect 97070 24436 97116 25238
rect 97070 24144 97080 24436
rect 97114 24144 97116 24436
rect 97070 23342 97116 24144
rect 97070 23050 97080 23342
rect 97114 23050 97116 23342
rect 97070 22248 97116 23050
rect 97070 21956 97080 22248
rect 97114 21956 97116 22248
rect 97070 21154 97116 21956
rect 97070 21096 97080 21154
rect 96056 20862 96084 20962
rect 89540 20664 93990 20754
rect 84894 20642 84976 20664
rect 89552 20658 93990 20664
rect 96002 20752 96084 20862
rect 97114 21096 97116 21154
rect 99170 25530 99254 25678
rect 98172 25238 98184 25442
rect 99170 25438 99196 25530
rect 98138 24436 98184 25238
rect 98172 24144 98184 24436
rect 98138 23342 98184 24144
rect 98172 23050 98184 23342
rect 98138 22248 98184 23050
rect 98172 21956 98184 22248
rect 98138 21154 98184 21956
rect 97080 20846 97114 20862
rect 98128 20862 98138 20934
rect 98172 21080 98184 21154
rect 99190 25238 99196 25438
rect 99230 25438 99254 25530
rect 100198 25530 100356 25678
rect 99230 25238 99236 25438
rect 100198 25370 100254 25530
rect 99190 24436 99236 25238
rect 99190 24144 99196 24436
rect 99230 24144 99236 24436
rect 99190 23342 99236 24144
rect 99190 23050 99196 23342
rect 99230 23050 99236 23342
rect 99190 22248 99236 23050
rect 99190 21956 99196 22248
rect 99230 21956 99236 22248
rect 99190 21154 99236 21956
rect 99190 21124 99196 21154
rect 98172 20862 98210 20934
rect 98128 20752 98210 20862
rect 99230 21124 99236 21154
rect 100246 25238 100254 25370
rect 100288 25370 100356 25530
rect 100288 25238 100292 25370
rect 100246 24436 100292 25238
rect 100246 24144 100254 24436
rect 100288 24144 100292 24436
rect 100246 23342 100292 24144
rect 100246 23050 100254 23342
rect 100288 23050 100292 23342
rect 100246 22248 100292 23050
rect 100246 21956 100254 22248
rect 100288 21956 100292 22248
rect 100246 21154 100292 21956
rect 100246 21096 100254 21154
rect 99196 20846 99230 20862
rect 100230 20862 100254 20956
rect 100288 21096 100292 21154
rect 100676 25188 101320 25566
rect 100676 21336 100720 25188
rect 101232 25032 101320 25188
rect 101276 21760 101320 25032
rect 101232 21336 101320 21760
rect 100676 21046 101320 21336
rect 100288 20862 100312 20956
rect 100230 20752 100312 20862
rect 96002 20662 100452 20752
rect 91666 20636 91748 20658
rect 96014 20656 100452 20662
rect 98128 20634 98210 20656
rect 62104 20008 62172 20018
rect 64208 20008 64276 20024
rect 66332 20008 66400 20040
rect 68568 20020 68636 20030
rect 70672 20020 70740 20036
rect 72796 20020 72864 20052
rect 68568 20010 72864 20020
rect 62104 19998 66400 20008
rect 61966 19954 66400 19998
rect 68430 19966 72864 20010
rect 75260 19980 75328 19990
rect 77364 19980 77432 19996
rect 79488 19980 79556 20012
rect 81724 19992 81792 20002
rect 83828 19992 83896 20008
rect 85952 19992 86020 20024
rect 81724 19982 86020 19992
rect 75260 19970 79556 19980
rect 61966 19918 66408 19954
rect 68430 19930 72872 19966
rect 68430 19920 72720 19930
rect 61966 19908 66256 19918
rect 59364 19676 59382 19760
rect 58358 19468 58364 19668
rect 58318 18666 58364 19468
rect 58318 18374 58324 18666
rect 58358 18374 58364 18666
rect 58318 17572 58364 18374
rect 58318 17280 58324 17572
rect 58358 17280 58364 17572
rect 58318 16478 58364 17280
rect 58318 16186 58324 16478
rect 58358 16186 58364 16478
rect 58318 15384 58364 16186
rect 58318 15354 58324 15384
rect 57300 15092 57338 15164
rect 57256 14982 57338 15092
rect 58358 15354 58364 15384
rect 59374 19468 59382 19676
rect 59416 19676 59460 19760
rect 62104 19730 62172 19908
rect 59416 19468 59420 19676
rect 59374 18666 59420 19468
rect 62104 19438 62118 19730
rect 62152 19628 62172 19730
rect 63176 19730 63210 19746
rect 62104 19422 62152 19438
rect 63172 19438 63176 19636
rect 64208 19730 64276 19908
rect 64208 19642 64234 19730
rect 63210 19438 63218 19636
rect 59374 18374 59382 18666
rect 59416 18374 59420 18666
rect 59374 17572 59420 18374
rect 59374 17280 59382 17572
rect 59416 17280 59420 17572
rect 59374 16478 59420 17280
rect 59628 18464 60002 18686
rect 59628 16980 59698 18464
rect 59892 16980 60002 18464
rect 62104 18652 62150 19422
rect 62104 18636 62152 18652
rect 62104 18344 62118 18636
rect 62104 18328 62152 18344
rect 63172 18636 63218 19438
rect 63172 18344 63176 18636
rect 63210 18344 63218 18636
rect 59628 16702 60002 16980
rect 61464 18196 61614 18322
rect 61464 17000 61486 18196
rect 61580 17000 61614 18196
rect 61464 16676 61614 17000
rect 62104 17558 62150 18328
rect 62104 17542 62152 17558
rect 62104 17250 62118 17542
rect 62104 17234 62152 17250
rect 63172 17542 63218 18344
rect 63172 17250 63176 17542
rect 63210 17250 63218 17542
rect 59374 16186 59382 16478
rect 59416 16186 59420 16478
rect 59374 15384 59420 16186
rect 59374 15326 59382 15384
rect 58324 15076 58358 15092
rect 59358 15092 59382 15186
rect 59416 15326 59420 15384
rect 62104 16464 62150 17234
rect 62104 16448 62152 16464
rect 62104 16156 62118 16448
rect 62104 16140 62152 16156
rect 63172 16448 63218 17250
rect 63172 16156 63176 16448
rect 63210 16156 63218 16448
rect 62104 15370 62150 16140
rect 62104 15354 62152 15370
rect 62104 15296 62118 15354
rect 59416 15092 59508 15192
rect 59358 14982 59508 15092
rect 63172 15354 63218 16156
rect 63172 15274 63176 15354
rect 62118 15046 62152 15062
rect 63156 15062 63176 15162
rect 63210 15274 63218 15354
rect 64224 19438 64234 19642
rect 64268 19694 64276 19730
rect 65292 19730 65326 19746
rect 64268 19642 64282 19694
rect 64268 19438 64270 19642
rect 64224 18636 64270 19438
rect 64224 18344 64234 18636
rect 64268 18344 64270 18636
rect 64224 17542 64270 18344
rect 64224 17250 64234 17542
rect 64268 17250 64270 17542
rect 64224 16448 64270 17250
rect 64224 16156 64234 16448
rect 64268 16156 64270 16448
rect 64224 15354 64270 16156
rect 64224 15296 64234 15354
rect 63210 15062 63238 15162
rect 55130 14892 59580 14982
rect 55142 14886 59580 14892
rect 63156 14952 63238 15062
rect 64268 15296 64270 15354
rect 66324 19730 66408 19918
rect 65326 19438 65338 19642
rect 66324 19638 66350 19730
rect 65292 18636 65338 19438
rect 65326 18344 65338 18636
rect 65292 17542 65338 18344
rect 65326 17250 65338 17542
rect 65292 16448 65338 17250
rect 65326 16156 65338 16448
rect 65292 15354 65338 16156
rect 64234 15046 64268 15062
rect 65282 15062 65292 15134
rect 65326 15280 65338 15354
rect 66344 19438 66350 19638
rect 66384 19638 66408 19730
rect 67408 19730 67442 19746
rect 66384 19438 66390 19638
rect 66344 18636 66390 19438
rect 66344 18344 66350 18636
rect 66384 18344 66390 18636
rect 66344 17542 66390 18344
rect 66344 17250 66350 17542
rect 66384 17250 66390 17542
rect 66344 16448 66390 17250
rect 66344 16156 66350 16448
rect 66384 16156 66390 16448
rect 66344 15354 66390 16156
rect 66344 15324 66350 15354
rect 65326 15062 65364 15134
rect 65282 14952 65364 15062
rect 66384 15324 66390 15354
rect 67400 19438 67408 19658
rect 68568 19742 68636 19920
rect 67442 19438 67446 19658
rect 67400 18636 67446 19438
rect 67400 18344 67408 18636
rect 67442 18344 67446 18636
rect 67400 17542 67446 18344
rect 68568 19450 68582 19742
rect 68616 19640 68636 19742
rect 69640 19742 69674 19758
rect 68568 19434 68616 19450
rect 69636 19450 69640 19648
rect 70672 19742 70740 19920
rect 70672 19654 70698 19742
rect 69674 19450 69682 19648
rect 68568 18664 68614 19434
rect 68568 18648 68616 18664
rect 68568 18356 68582 18648
rect 68568 18340 68616 18356
rect 69636 18648 69682 19450
rect 69636 18356 69640 18648
rect 69674 18356 69682 18648
rect 67400 17250 67408 17542
rect 67442 17250 67446 17542
rect 67400 16448 67446 17250
rect 67928 18208 68078 18334
rect 67928 17012 67950 18208
rect 68044 17012 68078 18208
rect 67928 16688 68078 17012
rect 68568 17570 68614 18340
rect 68568 17554 68616 17570
rect 68568 17262 68582 17554
rect 68568 17246 68616 17262
rect 69636 17554 69682 18356
rect 69636 17262 69640 17554
rect 69674 17262 69682 17554
rect 67400 16156 67408 16448
rect 67442 16156 67446 16448
rect 67400 15354 67446 16156
rect 67400 15296 67408 15354
rect 66350 15046 66384 15062
rect 67384 15062 67408 15156
rect 67442 15296 67446 15354
rect 68568 16476 68614 17246
rect 68568 16460 68616 16476
rect 68568 16168 68582 16460
rect 68568 16152 68616 16168
rect 69636 16460 69682 17262
rect 69636 16168 69640 16460
rect 69674 16168 69682 16460
rect 68568 15382 68614 16152
rect 68568 15366 68616 15382
rect 68568 15308 68582 15366
rect 67442 15062 67466 15156
rect 67384 14952 67466 15062
rect 69636 15366 69682 16168
rect 69636 15286 69640 15366
rect 68582 15058 68616 15074
rect 69620 15074 69640 15174
rect 69674 15286 69682 15366
rect 70688 19450 70698 19654
rect 70732 19706 70740 19742
rect 71756 19742 71790 19758
rect 70732 19654 70746 19706
rect 70732 19450 70734 19654
rect 70688 18648 70734 19450
rect 70688 18356 70698 18648
rect 70732 18356 70734 18648
rect 70688 17554 70734 18356
rect 70688 17262 70698 17554
rect 70732 17262 70734 17554
rect 70688 16460 70734 17262
rect 70688 16168 70698 16460
rect 70732 16168 70734 16460
rect 70688 15366 70734 16168
rect 70688 15308 70698 15366
rect 69674 15074 69702 15174
rect 69620 14964 69702 15074
rect 70732 15308 70734 15366
rect 72788 19742 72872 19930
rect 75122 19926 79556 19970
rect 81586 19938 86020 19982
rect 88494 19972 88562 19982
rect 90598 19972 90666 19988
rect 92722 19972 92790 20004
rect 94958 19984 95026 19994
rect 97062 19984 97130 20000
rect 99186 19984 99254 20016
rect 94958 19974 99254 19984
rect 88494 19962 92790 19972
rect 75122 19890 79564 19926
rect 81586 19902 86028 19938
rect 81586 19892 85876 19902
rect 75122 19880 79412 19890
rect 71790 19450 71802 19654
rect 72788 19650 72814 19742
rect 71756 18648 71802 19450
rect 71790 18356 71802 18648
rect 71756 17554 71802 18356
rect 71790 17262 71802 17554
rect 71756 16460 71802 17262
rect 71790 16168 71802 16460
rect 71756 15366 71802 16168
rect 70698 15058 70732 15074
rect 71746 15074 71756 15146
rect 71790 15292 71802 15366
rect 72808 19450 72814 19650
rect 72848 19650 72872 19742
rect 73872 19742 73906 19758
rect 72848 19450 72854 19650
rect 72808 18648 72854 19450
rect 72808 18356 72814 18648
rect 72848 18356 72854 18648
rect 72808 17554 72854 18356
rect 72808 17262 72814 17554
rect 72848 17262 72854 17554
rect 72808 16460 72854 17262
rect 72808 16168 72814 16460
rect 72848 16168 72854 16460
rect 72808 15366 72854 16168
rect 72808 15336 72814 15366
rect 71790 15074 71828 15146
rect 71746 14964 71828 15074
rect 72848 15336 72854 15366
rect 73864 19450 73872 19670
rect 75260 19702 75328 19880
rect 73906 19450 73910 19670
rect 73864 18648 73910 19450
rect 73864 18356 73872 18648
rect 73906 18356 73910 18648
rect 73864 17554 73910 18356
rect 75260 19410 75274 19702
rect 75308 19600 75328 19702
rect 76332 19702 76366 19718
rect 75260 19394 75308 19410
rect 76328 19410 76332 19608
rect 77364 19702 77432 19880
rect 77364 19614 77390 19702
rect 76366 19410 76374 19608
rect 75260 18624 75306 19394
rect 75260 18608 75308 18624
rect 75260 18316 75274 18608
rect 75260 18300 75308 18316
rect 76328 18608 76374 19410
rect 76328 18316 76332 18608
rect 76366 18316 76374 18608
rect 73864 17262 73872 17554
rect 73906 17262 73910 17554
rect 73864 16460 73910 17262
rect 74620 18168 74770 18294
rect 74620 16972 74642 18168
rect 74736 16972 74770 18168
rect 74620 16648 74770 16972
rect 75260 17530 75306 18300
rect 75260 17514 75308 17530
rect 75260 17222 75274 17514
rect 75260 17206 75308 17222
rect 76328 17514 76374 18316
rect 76328 17222 76332 17514
rect 76366 17222 76374 17514
rect 73864 16168 73872 16460
rect 73906 16168 73910 16460
rect 73864 15366 73910 16168
rect 73864 15308 73872 15366
rect 72814 15058 72848 15074
rect 73848 15074 73872 15168
rect 73906 15308 73910 15366
rect 75260 16436 75306 17206
rect 75260 16420 75308 16436
rect 75260 16128 75274 16420
rect 75260 16112 75308 16128
rect 76328 16420 76374 17222
rect 76328 16128 76332 16420
rect 76366 16128 76374 16420
rect 75260 15342 75306 16112
rect 75260 15326 75308 15342
rect 75260 15268 75274 15326
rect 73906 15074 73930 15168
rect 73848 14964 73930 15074
rect 76328 15326 76374 16128
rect 76328 15246 76332 15326
rect 75274 15018 75308 15034
rect 76312 15034 76332 15134
rect 76366 15246 76374 15326
rect 77380 19410 77390 19614
rect 77424 19666 77432 19702
rect 78448 19702 78482 19718
rect 77424 19614 77438 19666
rect 77424 19410 77426 19614
rect 77380 18608 77426 19410
rect 77380 18316 77390 18608
rect 77424 18316 77426 18608
rect 77380 17514 77426 18316
rect 77380 17222 77390 17514
rect 77424 17222 77426 17514
rect 77380 16420 77426 17222
rect 77380 16128 77390 16420
rect 77424 16128 77426 16420
rect 77380 15326 77426 16128
rect 77380 15268 77390 15326
rect 76366 15034 76394 15134
rect 57256 14864 57338 14886
rect 56192 14182 56260 14198
rect 58316 14182 58384 14214
rect 54038 14172 58384 14182
rect 53950 14128 58384 14172
rect 53950 14092 58392 14128
rect 53950 14082 58240 14092
rect 54038 13976 54164 14082
rect 50796 13598 50808 13802
rect 51794 13798 51820 13890
rect 50762 12796 50808 13598
rect 50796 12504 50808 12796
rect 50762 11702 50808 12504
rect 50796 11410 50808 11702
rect 50762 10608 50808 11410
rect 50796 10316 50808 10608
rect 50762 9514 50808 10316
rect 49704 9206 49738 9222
rect 50752 9222 50762 9294
rect 50796 9440 50808 9514
rect 51814 13598 51820 13798
rect 51854 13798 51878 13890
rect 52878 13890 52912 13906
rect 51854 13598 51860 13798
rect 51814 12796 51860 13598
rect 51814 12504 51820 12796
rect 51854 12504 51860 12796
rect 51814 11702 51860 12504
rect 51814 11410 51820 11702
rect 51854 11410 51860 11702
rect 51814 10608 51860 11410
rect 51814 10316 51820 10608
rect 51854 10316 51860 10608
rect 51814 9514 51860 10316
rect 51814 9484 51820 9514
rect 50796 9222 50834 9294
rect 50752 9112 50834 9222
rect 51854 9484 51860 9514
rect 52870 13598 52878 13818
rect 54088 13904 54156 13976
rect 52912 13598 52916 13818
rect 52870 12796 52916 13598
rect 52870 12504 52878 12796
rect 52912 12504 52916 12796
rect 52870 11702 52916 12504
rect 54088 13612 54102 13904
rect 54136 13802 54156 13904
rect 55160 13904 55194 13920
rect 54088 13596 54136 13612
rect 55156 13612 55160 13810
rect 56192 13904 56260 14082
rect 56192 13816 56218 13904
rect 55194 13612 55202 13810
rect 54088 12826 54134 13596
rect 54088 12810 54136 12826
rect 54088 12518 54102 12810
rect 54088 12502 54136 12518
rect 55156 12810 55202 13612
rect 55156 12518 55160 12810
rect 55194 12518 55202 12810
rect 52870 11410 52878 11702
rect 52912 11410 52916 11702
rect 52870 10608 52916 11410
rect 53448 12370 53598 12496
rect 53448 11174 53470 12370
rect 53564 11174 53598 12370
rect 53448 10850 53598 11174
rect 54088 11732 54134 12502
rect 54088 11716 54136 11732
rect 54088 11424 54102 11716
rect 54088 11408 54136 11424
rect 55156 11716 55202 12518
rect 55156 11424 55160 11716
rect 55194 11424 55202 11716
rect 52870 10316 52878 10608
rect 52912 10316 52916 10608
rect 52870 9514 52916 10316
rect 52870 9456 52878 9514
rect 51820 9206 51854 9222
rect 52854 9222 52878 9316
rect 52912 9456 52916 9514
rect 54088 10638 54134 11408
rect 54088 10622 54136 10638
rect 54088 10330 54102 10622
rect 54088 10314 54136 10330
rect 55156 10622 55202 11424
rect 55156 10330 55160 10622
rect 55194 10330 55202 10622
rect 54088 9544 54134 10314
rect 54088 9528 54136 9544
rect 54088 9488 54102 9528
rect 52912 9222 52936 9316
rect 52854 9174 52936 9222
rect 54052 9236 54102 9488
rect 55156 9528 55202 10330
rect 54136 9454 54176 9488
rect 54136 9236 54178 9454
rect 55156 9448 55160 9528
rect 52854 9112 52998 9174
rect 48626 9022 53076 9112
rect 48638 9016 53076 9022
rect 50752 8994 50834 9016
rect 49696 8260 49764 8276
rect 51820 8260 51888 8292
rect 47542 8250 51888 8260
rect 47454 8206 51888 8250
rect 47454 8170 51896 8206
rect 47454 8160 51744 8170
rect 47542 8014 47668 8160
rect 45284 7668 45290 7868
rect 46256 7726 46308 7960
rect 45244 6866 45290 7668
rect 45244 6574 45250 6866
rect 45284 6574 45290 6866
rect 45244 5772 45290 6574
rect 45244 5480 45250 5772
rect 45284 5480 45290 5772
rect 45244 4678 45290 5480
rect 45244 4386 45250 4678
rect 45284 4386 45290 4678
rect 45244 3584 45290 4386
rect 45244 3554 45250 3584
rect 44226 3292 44264 3364
rect 44182 3182 44264 3292
rect 45284 3554 45290 3584
rect 46300 7668 46308 7726
rect 46342 7726 46382 7960
rect 47592 7982 47660 8014
rect 46342 7668 46346 7726
rect 46300 6866 46346 7668
rect 46300 6574 46308 6866
rect 46342 6574 46346 6866
rect 47592 7690 47606 7982
rect 47640 7880 47660 7982
rect 48664 7982 48698 7998
rect 47592 7674 47640 7690
rect 48660 7690 48664 7888
rect 49696 7982 49764 8160
rect 49696 7894 49722 7982
rect 48698 7690 48706 7888
rect 47592 6904 47638 7674
rect 47592 6888 47640 6904
rect 47592 6596 47606 6888
rect 47592 6580 47640 6596
rect 48660 6888 48706 7690
rect 48660 6596 48664 6888
rect 48698 6596 48706 6888
rect 46300 5772 46346 6574
rect 46300 5480 46308 5772
rect 46342 5480 46346 5772
rect 46300 4678 46346 5480
rect 46952 6448 47102 6574
rect 46952 5252 46974 6448
rect 47068 5252 47102 6448
rect 46952 4928 47102 5252
rect 47592 5810 47638 6580
rect 47592 5794 47640 5810
rect 47592 5502 47606 5794
rect 47592 5486 47640 5502
rect 48660 5794 48706 6596
rect 48660 5502 48664 5794
rect 48698 5502 48706 5794
rect 46300 4386 46308 4678
rect 46342 4386 46346 4678
rect 46300 3584 46346 4386
rect 46300 3526 46308 3584
rect 45250 3276 45284 3292
rect 46284 3292 46308 3386
rect 46342 3526 46346 3584
rect 47592 4716 47638 5486
rect 47592 4700 47640 4716
rect 47592 4408 47606 4700
rect 47592 4392 47640 4408
rect 48660 4700 48706 5502
rect 48660 4408 48664 4700
rect 48698 4408 48706 4700
rect 47592 3622 47638 4392
rect 47592 3606 47640 3622
rect 47592 3548 47606 3606
rect 46342 3292 46366 3386
rect 48660 3606 48706 4408
rect 48660 3526 48664 3606
rect 47606 3298 47640 3314
rect 48644 3314 48664 3414
rect 48698 3526 48706 3606
rect 49712 7690 49722 7894
rect 49756 7946 49764 7982
rect 50780 7982 50814 7998
rect 49756 7894 49770 7946
rect 49756 7690 49758 7894
rect 49712 6888 49758 7690
rect 49712 6596 49722 6888
rect 49756 6596 49758 6888
rect 49712 5794 49758 6596
rect 49712 5502 49722 5794
rect 49756 5502 49758 5794
rect 49712 4700 49758 5502
rect 49712 4408 49722 4700
rect 49756 4408 49758 4700
rect 49712 3606 49758 4408
rect 49712 3548 49722 3606
rect 48698 3314 48726 3414
rect 46284 3248 46366 3292
rect 48644 3248 48726 3314
rect 49756 3548 49758 3606
rect 51812 7982 51896 8170
rect 50814 7690 50826 7894
rect 51812 7890 51838 7982
rect 50780 6888 50826 7690
rect 50814 6596 50826 6888
rect 50780 5794 50826 6596
rect 50814 5502 50826 5794
rect 50780 4700 50826 5502
rect 50814 4408 50826 4700
rect 50780 3606 50826 4408
rect 49722 3298 49756 3314
rect 50770 3314 50780 3386
rect 50814 3532 50826 3606
rect 51832 7690 51838 7890
rect 51872 7890 51896 7982
rect 52872 7982 52998 9016
rect 54052 8274 54178 9236
rect 55140 9236 55160 9336
rect 55194 9448 55202 9528
rect 56208 13612 56218 13816
rect 56252 13868 56260 13904
rect 57276 13904 57310 13920
rect 56252 13816 56266 13868
rect 56252 13612 56254 13816
rect 56208 12810 56254 13612
rect 56208 12518 56218 12810
rect 56252 12518 56254 12810
rect 56208 11716 56254 12518
rect 56208 11424 56218 11716
rect 56252 11424 56254 11716
rect 56208 10622 56254 11424
rect 56208 10330 56218 10622
rect 56252 10330 56254 10622
rect 56208 9528 56254 10330
rect 56208 9470 56218 9528
rect 55194 9236 55222 9336
rect 55140 9126 55222 9236
rect 56252 9470 56254 9528
rect 58308 13904 58392 14092
rect 57310 13612 57322 13816
rect 58308 13812 58334 13904
rect 57276 12810 57322 13612
rect 57310 12518 57322 12810
rect 57276 11716 57322 12518
rect 57310 11424 57322 11716
rect 57276 10622 57322 11424
rect 57310 10330 57322 10622
rect 57276 9528 57322 10330
rect 56218 9220 56252 9236
rect 57266 9236 57276 9308
rect 57310 9454 57322 9528
rect 58328 13612 58334 13812
rect 58368 13812 58392 13904
rect 59382 13904 59508 14886
rect 63156 14862 67606 14952
rect 69620 14874 74070 14964
rect 69632 14868 74070 14874
rect 76312 14924 76394 15034
rect 77424 15268 77426 15326
rect 79480 19702 79564 19890
rect 78482 19410 78494 19614
rect 79480 19610 79506 19702
rect 78448 18608 78494 19410
rect 78482 18316 78494 18608
rect 78448 17514 78494 18316
rect 78482 17222 78494 17514
rect 78448 16420 78494 17222
rect 78482 16128 78494 16420
rect 78448 15326 78494 16128
rect 77390 15018 77424 15034
rect 78438 15034 78448 15106
rect 78482 15252 78494 15326
rect 79500 19410 79506 19610
rect 79540 19610 79564 19702
rect 80564 19702 80598 19718
rect 79540 19410 79546 19610
rect 79500 18608 79546 19410
rect 79500 18316 79506 18608
rect 79540 18316 79546 18608
rect 79500 17514 79546 18316
rect 79500 17222 79506 17514
rect 79540 17222 79546 17514
rect 79500 16420 79546 17222
rect 79500 16128 79506 16420
rect 79540 16128 79546 16420
rect 79500 15326 79546 16128
rect 79500 15296 79506 15326
rect 78482 15034 78520 15106
rect 78438 14924 78520 15034
rect 79540 15296 79546 15326
rect 80556 19410 80564 19630
rect 81724 19714 81792 19892
rect 80598 19410 80602 19630
rect 80556 18608 80602 19410
rect 80556 18316 80564 18608
rect 80598 18316 80602 18608
rect 80556 17514 80602 18316
rect 81724 19422 81738 19714
rect 81772 19612 81792 19714
rect 82796 19714 82830 19730
rect 81724 19406 81772 19422
rect 82792 19422 82796 19620
rect 83828 19714 83896 19892
rect 83828 19626 83854 19714
rect 82830 19422 82838 19620
rect 81724 18636 81770 19406
rect 81724 18620 81772 18636
rect 81724 18328 81738 18620
rect 81724 18312 81772 18328
rect 82792 18620 82838 19422
rect 82792 18328 82796 18620
rect 82830 18328 82838 18620
rect 80556 17222 80564 17514
rect 80598 17222 80602 17514
rect 80556 16420 80602 17222
rect 81084 18180 81234 18306
rect 81084 16984 81106 18180
rect 81200 16984 81234 18180
rect 81084 16660 81234 16984
rect 81724 17542 81770 18312
rect 81724 17526 81772 17542
rect 81724 17234 81738 17526
rect 81724 17218 81772 17234
rect 82792 17526 82838 18328
rect 82792 17234 82796 17526
rect 82830 17234 82838 17526
rect 80556 16128 80564 16420
rect 80598 16128 80602 16420
rect 80556 15326 80602 16128
rect 80556 15268 80564 15326
rect 79506 15018 79540 15034
rect 80540 15034 80564 15128
rect 80598 15268 80602 15326
rect 81724 16448 81770 17218
rect 81724 16432 81772 16448
rect 81724 16140 81738 16432
rect 81724 16124 81772 16140
rect 82792 16432 82838 17234
rect 82792 16140 82796 16432
rect 82830 16140 82838 16432
rect 81724 15354 81770 16124
rect 81724 15338 81772 15354
rect 81724 15280 81738 15338
rect 80598 15034 80622 15128
rect 80540 14924 80622 15034
rect 82792 15338 82838 16140
rect 82792 15258 82796 15338
rect 81738 15030 81772 15046
rect 82776 15046 82796 15146
rect 82830 15258 82838 15338
rect 83844 19422 83854 19626
rect 83888 19678 83896 19714
rect 84912 19714 84946 19730
rect 83888 19626 83902 19678
rect 83888 19422 83890 19626
rect 83844 18620 83890 19422
rect 83844 18328 83854 18620
rect 83888 18328 83890 18620
rect 83844 17526 83890 18328
rect 83844 17234 83854 17526
rect 83888 17234 83890 17526
rect 83844 16432 83890 17234
rect 83844 16140 83854 16432
rect 83888 16140 83890 16432
rect 83844 15338 83890 16140
rect 83844 15280 83854 15338
rect 82830 15046 82858 15146
rect 82776 14936 82858 15046
rect 83888 15280 83890 15338
rect 85944 19714 86028 19902
rect 88356 19918 92790 19962
rect 94820 19930 99254 19974
rect 88356 19882 92798 19918
rect 94820 19894 99262 19930
rect 94820 19884 99110 19894
rect 88356 19872 92646 19882
rect 84946 19422 84958 19626
rect 85944 19622 85970 19714
rect 84912 18620 84958 19422
rect 84946 18328 84958 18620
rect 84912 17526 84958 18328
rect 84946 17234 84958 17526
rect 84912 16432 84958 17234
rect 84946 16140 84958 16432
rect 84912 15338 84958 16140
rect 83854 15030 83888 15046
rect 84902 15046 84912 15118
rect 84946 15264 84958 15338
rect 85964 19422 85970 19622
rect 86004 19622 86028 19714
rect 87028 19714 87062 19730
rect 86004 19422 86010 19622
rect 85964 18620 86010 19422
rect 85964 18328 85970 18620
rect 86004 18328 86010 18620
rect 85964 17526 86010 18328
rect 85964 17234 85970 17526
rect 86004 17234 86010 17526
rect 85964 16432 86010 17234
rect 85964 16140 85970 16432
rect 86004 16140 86010 16432
rect 85964 15338 86010 16140
rect 85964 15308 85970 15338
rect 84946 15046 84984 15118
rect 84902 14936 84984 15046
rect 86004 15308 86010 15338
rect 87020 19422 87028 19642
rect 88494 19694 88562 19872
rect 87062 19422 87066 19642
rect 87020 18620 87066 19422
rect 87020 18328 87028 18620
rect 87062 18328 87066 18620
rect 87020 17526 87066 18328
rect 88494 19402 88508 19694
rect 88542 19592 88562 19694
rect 89566 19694 89600 19710
rect 88494 19386 88542 19402
rect 89562 19402 89566 19600
rect 90598 19694 90666 19872
rect 90598 19606 90624 19694
rect 89600 19402 89608 19600
rect 88494 18616 88540 19386
rect 88494 18600 88542 18616
rect 88494 18308 88508 18600
rect 88494 18292 88542 18308
rect 89562 18600 89608 19402
rect 89562 18308 89566 18600
rect 89600 18308 89608 18600
rect 87020 17234 87028 17526
rect 87062 17234 87066 17526
rect 87020 16432 87066 17234
rect 87854 18160 88004 18286
rect 87854 16964 87876 18160
rect 87970 16964 88004 18160
rect 87854 16640 88004 16964
rect 88494 17522 88540 18292
rect 88494 17506 88542 17522
rect 88494 17214 88508 17506
rect 88494 17198 88542 17214
rect 89562 17506 89608 18308
rect 89562 17214 89566 17506
rect 89600 17214 89608 17506
rect 87020 16140 87028 16432
rect 87062 16140 87066 16432
rect 87020 15338 87066 16140
rect 87020 15280 87028 15338
rect 85970 15030 86004 15046
rect 87004 15046 87028 15140
rect 87062 15280 87066 15338
rect 88494 16428 88540 17198
rect 88494 16412 88542 16428
rect 88494 16120 88508 16412
rect 88494 16104 88542 16120
rect 89562 16412 89608 17214
rect 89562 16120 89566 16412
rect 89600 16120 89608 16412
rect 88494 15334 88540 16104
rect 88494 15318 88542 15334
rect 88494 15260 88508 15318
rect 87062 15046 87086 15140
rect 87004 14936 87086 15046
rect 89562 15318 89608 16120
rect 89562 15238 89566 15318
rect 88508 15010 88542 15026
rect 89546 15026 89566 15126
rect 89600 15238 89608 15318
rect 90614 19402 90624 19606
rect 90658 19658 90666 19694
rect 91682 19694 91716 19710
rect 90658 19606 90672 19658
rect 90658 19402 90660 19606
rect 90614 18600 90660 19402
rect 90614 18308 90624 18600
rect 90658 18308 90660 18600
rect 90614 17506 90660 18308
rect 90614 17214 90624 17506
rect 90658 17214 90660 17506
rect 90614 16412 90660 17214
rect 90614 16120 90624 16412
rect 90658 16120 90660 16412
rect 90614 15318 90660 16120
rect 90614 15260 90624 15318
rect 89600 15026 89628 15126
rect 63168 14856 67606 14862
rect 65282 14834 65364 14856
rect 71746 14846 71828 14868
rect 76312 14834 80762 14924
rect 82776 14846 87226 14936
rect 82788 14840 87226 14846
rect 89546 14916 89628 15026
rect 90658 15260 90660 15318
rect 92714 19694 92798 19882
rect 91716 19402 91728 19606
rect 92714 19602 92740 19694
rect 91682 18600 91728 19402
rect 91716 18308 91728 18600
rect 91682 17506 91728 18308
rect 91716 17214 91728 17506
rect 91682 16412 91728 17214
rect 91716 16120 91728 16412
rect 91682 15318 91728 16120
rect 90624 15010 90658 15026
rect 91672 15026 91682 15098
rect 91716 15244 91728 15318
rect 92734 19402 92740 19602
rect 92774 19602 92798 19694
rect 93798 19694 93832 19710
rect 92774 19402 92780 19602
rect 92734 18600 92780 19402
rect 92734 18308 92740 18600
rect 92774 18308 92780 18600
rect 92734 17506 92780 18308
rect 92734 17214 92740 17506
rect 92774 17214 92780 17506
rect 92734 16412 92780 17214
rect 92734 16120 92740 16412
rect 92774 16120 92780 16412
rect 92734 15318 92780 16120
rect 92734 15288 92740 15318
rect 91716 15026 91754 15098
rect 91672 14916 91754 15026
rect 92774 15288 92780 15318
rect 93790 19402 93798 19622
rect 94958 19706 95026 19884
rect 93832 19402 93836 19622
rect 93790 18600 93836 19402
rect 93790 18308 93798 18600
rect 93832 18308 93836 18600
rect 93790 17506 93836 18308
rect 94958 19414 94972 19706
rect 95006 19604 95026 19706
rect 96030 19706 96064 19722
rect 94958 19398 95006 19414
rect 96026 19414 96030 19612
rect 97062 19706 97130 19884
rect 97062 19618 97088 19706
rect 96064 19414 96072 19612
rect 94958 18628 95004 19398
rect 94958 18612 95006 18628
rect 94958 18320 94972 18612
rect 94958 18304 95006 18320
rect 96026 18612 96072 19414
rect 96026 18320 96030 18612
rect 96064 18320 96072 18612
rect 93790 17214 93798 17506
rect 93832 17214 93836 17506
rect 93790 16412 93836 17214
rect 94318 18172 94468 18298
rect 94318 16976 94340 18172
rect 94434 16976 94468 18172
rect 94318 16652 94468 16976
rect 94958 17534 95004 18304
rect 94958 17518 95006 17534
rect 94958 17226 94972 17518
rect 94958 17210 95006 17226
rect 96026 17518 96072 18320
rect 96026 17226 96030 17518
rect 96064 17226 96072 17518
rect 93790 16120 93798 16412
rect 93832 16120 93836 16412
rect 93790 15318 93836 16120
rect 93790 15260 93798 15318
rect 92740 15010 92774 15026
rect 93774 15026 93798 15120
rect 93832 15260 93836 15318
rect 94958 16440 95004 17210
rect 94958 16424 95006 16440
rect 94958 16132 94972 16424
rect 94958 16116 95006 16132
rect 96026 16424 96072 17226
rect 96026 16132 96030 16424
rect 96064 16132 96072 16424
rect 94958 15346 95004 16116
rect 94958 15330 95006 15346
rect 94958 15272 94972 15330
rect 93832 15026 93856 15120
rect 93774 14916 93856 15026
rect 96026 15330 96072 16132
rect 96026 15250 96030 15330
rect 94972 15022 95006 15038
rect 96010 15038 96030 15138
rect 96064 15250 96072 15330
rect 97078 19414 97088 19618
rect 97122 19670 97130 19706
rect 98146 19706 98180 19722
rect 97122 19618 97136 19670
rect 97122 19414 97124 19618
rect 97078 18612 97124 19414
rect 97078 18320 97088 18612
rect 97122 18320 97124 18612
rect 97078 17518 97124 18320
rect 97078 17226 97088 17518
rect 97122 17226 97124 17518
rect 97078 16424 97124 17226
rect 97078 16132 97088 16424
rect 97122 16132 97124 16424
rect 97078 15330 97124 16132
rect 97078 15272 97088 15330
rect 96064 15038 96092 15138
rect 96010 14928 96092 15038
rect 97122 15272 97124 15330
rect 99178 19706 99262 19894
rect 98180 19414 98192 19618
rect 99178 19614 99204 19706
rect 98146 18612 98192 19414
rect 98180 18320 98192 18612
rect 98146 17518 98192 18320
rect 98180 17226 98192 17518
rect 98146 16424 98192 17226
rect 98180 16132 98192 16424
rect 98146 15330 98192 16132
rect 97088 15022 97122 15038
rect 98136 15038 98146 15110
rect 98180 15256 98192 15330
rect 99198 19414 99204 19614
rect 99238 19614 99262 19706
rect 100262 19706 100296 19722
rect 99238 19414 99244 19614
rect 99198 18612 99244 19414
rect 99198 18320 99204 18612
rect 99238 18320 99244 18612
rect 99198 17518 99244 18320
rect 99198 17226 99204 17518
rect 99238 17226 99244 17518
rect 99198 16424 99244 17226
rect 99198 16132 99204 16424
rect 99238 16132 99244 16424
rect 99198 15330 99244 16132
rect 99198 15300 99204 15330
rect 98180 15038 98218 15110
rect 98136 14928 98218 15038
rect 99238 15300 99244 15330
rect 100254 19414 100262 19634
rect 100296 19414 100300 19634
rect 100254 18612 100300 19414
rect 100254 18320 100262 18612
rect 100296 18320 100300 18612
rect 100254 17518 100300 18320
rect 100254 17226 100262 17518
rect 100296 17226 100300 17518
rect 100254 16424 100300 17226
rect 100254 16132 100262 16424
rect 100296 16132 100300 16424
rect 100254 15330 100300 16132
rect 100254 15272 100262 15330
rect 99204 15022 99238 15038
rect 100238 15038 100262 15132
rect 100296 15272 100300 15330
rect 100630 19110 101276 19266
rect 100296 15038 100320 15132
rect 100238 14928 100320 15038
rect 100630 14992 100698 19110
rect 101188 14992 101276 19110
rect 76324 14828 80762 14834
rect 78438 14806 78520 14828
rect 84902 14818 84984 14840
rect 89546 14826 93996 14916
rect 96010 14838 100460 14928
rect 100630 14880 101276 14992
rect 96022 14832 100460 14838
rect 89558 14820 93996 14826
rect 91672 14798 91754 14820
rect 98136 14810 98218 14832
rect 62104 14150 62172 14160
rect 64208 14150 64276 14166
rect 66332 14150 66400 14182
rect 62104 14140 66400 14150
rect 61966 14096 66400 14140
rect 68572 14148 68640 14158
rect 70676 14148 70744 14164
rect 72800 14148 72868 14180
rect 68572 14138 72868 14148
rect 61966 14060 66408 14096
rect 61966 14050 66256 14060
rect 58368 13612 58374 13812
rect 59382 13808 59392 13904
rect 58328 12810 58374 13612
rect 58328 12518 58334 12810
rect 58368 12518 58374 12810
rect 58328 11716 58374 12518
rect 58328 11424 58334 11716
rect 58368 11424 58374 11716
rect 58328 10622 58374 11424
rect 58328 10330 58334 10622
rect 58368 10330 58374 10622
rect 58328 9528 58374 10330
rect 58328 9498 58334 9528
rect 57310 9236 57348 9308
rect 57266 9126 57348 9236
rect 58368 9498 58374 9528
rect 59384 13612 59392 13808
rect 59426 13808 59508 13904
rect 62104 13872 62172 14050
rect 59426 13612 59430 13808
rect 59384 12810 59430 13612
rect 59384 12518 59392 12810
rect 59426 12518 59430 12810
rect 62104 13580 62118 13872
rect 62152 13770 62172 13872
rect 63176 13872 63210 13888
rect 62104 13564 62152 13580
rect 63172 13580 63176 13778
rect 64208 13872 64276 14050
rect 64208 13784 64234 13872
rect 63210 13580 63218 13778
rect 62104 12794 62150 13564
rect 62104 12778 62152 12794
rect 59384 11716 59430 12518
rect 59384 11424 59392 11716
rect 59426 11424 59430 11716
rect 59384 10622 59430 11424
rect 59642 12542 60002 12694
rect 59642 11168 59698 12542
rect 59934 11168 60002 12542
rect 62104 12486 62118 12778
rect 62104 12470 62152 12486
rect 63172 12778 63218 13580
rect 63172 12486 63176 12778
rect 63210 12486 63218 12778
rect 59642 11002 60002 11168
rect 61464 12338 61614 12464
rect 61464 11142 61486 12338
rect 61580 11142 61614 12338
rect 61464 10818 61614 11142
rect 62104 11700 62150 12470
rect 62104 11684 62152 11700
rect 62104 11392 62118 11684
rect 62104 11376 62152 11392
rect 63172 11684 63218 12486
rect 63172 11392 63176 11684
rect 63210 11392 63218 11684
rect 59384 10330 59392 10622
rect 59426 10330 59430 10622
rect 59384 9528 59430 10330
rect 59384 9470 59392 9528
rect 58334 9220 58368 9236
rect 59368 9236 59392 9330
rect 59426 9470 59430 9528
rect 62104 10606 62150 11376
rect 62104 10590 62152 10606
rect 62104 10298 62118 10590
rect 62104 10282 62152 10298
rect 63172 10590 63218 11392
rect 63172 10298 63176 10590
rect 63210 10298 63218 10590
rect 62104 9512 62150 10282
rect 62104 9496 62152 9512
rect 62104 9438 62118 9496
rect 59426 9236 59450 9330
rect 59368 9216 59450 9236
rect 59368 9126 59494 9216
rect 63172 9496 63218 10298
rect 63172 9416 63176 9496
rect 62118 9188 62152 9204
rect 63156 9204 63176 9304
rect 63210 9416 63218 9496
rect 64224 13580 64234 13784
rect 64268 13836 64276 13872
rect 65292 13872 65326 13888
rect 64268 13784 64282 13836
rect 64268 13580 64270 13784
rect 64224 12778 64270 13580
rect 64224 12486 64234 12778
rect 64268 12486 64270 12778
rect 64224 11684 64270 12486
rect 64224 11392 64234 11684
rect 64268 11392 64270 11684
rect 64224 10590 64270 11392
rect 64224 10298 64234 10590
rect 64268 10298 64270 10590
rect 64224 9496 64270 10298
rect 64224 9438 64234 9496
rect 63210 9204 63238 9304
rect 55140 9036 59590 9126
rect 55152 9030 59590 9036
rect 63156 9094 63238 9204
rect 64268 9438 64270 9496
rect 66324 13872 66408 14060
rect 68434 14094 72868 14138
rect 75260 14122 75328 14132
rect 77364 14122 77432 14138
rect 79488 14122 79556 14154
rect 75260 14112 79556 14122
rect 68434 14058 72876 14094
rect 68434 14048 72724 14058
rect 65326 13580 65338 13784
rect 66324 13780 66350 13872
rect 65292 12778 65338 13580
rect 65326 12486 65338 12778
rect 65292 11684 65338 12486
rect 65326 11392 65338 11684
rect 65292 10590 65338 11392
rect 65326 10298 65338 10590
rect 65292 9496 65338 10298
rect 64234 9188 64268 9204
rect 65282 9204 65292 9276
rect 65326 9422 65338 9496
rect 66344 13580 66350 13780
rect 66384 13780 66408 13872
rect 67408 13872 67442 13888
rect 66384 13580 66390 13780
rect 66344 12778 66390 13580
rect 66344 12486 66350 12778
rect 66384 12486 66390 12778
rect 66344 11684 66390 12486
rect 66344 11392 66350 11684
rect 66384 11392 66390 11684
rect 66344 10590 66390 11392
rect 66344 10298 66350 10590
rect 66384 10298 66390 10590
rect 66344 9496 66390 10298
rect 66344 9466 66350 9496
rect 65326 9204 65364 9276
rect 65282 9094 65364 9204
rect 66384 9466 66390 9496
rect 67400 13580 67408 13800
rect 68572 13870 68640 14048
rect 67442 13580 67446 13800
rect 67400 12778 67446 13580
rect 67400 12486 67408 12778
rect 67442 12486 67446 12778
rect 67400 11684 67446 12486
rect 68572 13578 68586 13870
rect 68620 13768 68640 13870
rect 69644 13870 69678 13886
rect 68572 13562 68620 13578
rect 69640 13578 69644 13776
rect 70676 13870 70744 14048
rect 70676 13782 70702 13870
rect 69678 13578 69686 13776
rect 68572 12792 68618 13562
rect 68572 12776 68620 12792
rect 68572 12484 68586 12776
rect 68572 12468 68620 12484
rect 69640 12776 69686 13578
rect 69640 12484 69644 12776
rect 69678 12484 69686 12776
rect 67400 11392 67408 11684
rect 67442 11392 67446 11684
rect 67400 10590 67446 11392
rect 67932 12336 68082 12462
rect 67932 11140 67954 12336
rect 68048 11140 68082 12336
rect 67932 10816 68082 11140
rect 68572 11698 68618 12468
rect 68572 11682 68620 11698
rect 68572 11390 68586 11682
rect 68572 11374 68620 11390
rect 69640 11682 69686 12484
rect 69640 11390 69644 11682
rect 69678 11390 69686 11682
rect 67400 10298 67408 10590
rect 67442 10298 67446 10590
rect 67400 9496 67446 10298
rect 67400 9438 67408 9496
rect 66350 9188 66384 9204
rect 67384 9204 67408 9298
rect 67442 9438 67446 9496
rect 68572 10604 68618 11374
rect 68572 10588 68620 10604
rect 68572 10296 68586 10588
rect 68572 10280 68620 10296
rect 69640 10588 69686 11390
rect 69640 10296 69644 10588
rect 69678 10296 69686 10588
rect 68572 9510 68618 10280
rect 68572 9494 68620 9510
rect 68572 9436 68586 9494
rect 67442 9204 67466 9298
rect 67384 9094 67466 9204
rect 69640 9494 69686 10296
rect 69640 9414 69644 9494
rect 68586 9186 68620 9202
rect 69624 9202 69644 9302
rect 69678 9414 69686 9494
rect 70692 13578 70702 13782
rect 70736 13834 70744 13870
rect 71760 13870 71794 13886
rect 70736 13782 70750 13834
rect 70736 13578 70738 13782
rect 70692 12776 70738 13578
rect 70692 12484 70702 12776
rect 70736 12484 70738 12776
rect 70692 11682 70738 12484
rect 70692 11390 70702 11682
rect 70736 11390 70738 11682
rect 70692 10588 70738 11390
rect 70692 10296 70702 10588
rect 70736 10296 70738 10588
rect 70692 9494 70738 10296
rect 70692 9436 70702 9494
rect 69678 9202 69706 9302
rect 57266 9008 57348 9030
rect 56210 8274 56278 8290
rect 58334 8274 58402 8306
rect 54052 8264 58402 8274
rect 53968 8220 58402 8264
rect 53968 8184 58410 8220
rect 53968 8174 58258 8184
rect 54052 8070 54178 8174
rect 51872 7690 51878 7890
rect 52872 7790 52896 7982
rect 51832 6888 51878 7690
rect 51832 6596 51838 6888
rect 51872 6596 51878 6888
rect 51832 5794 51878 6596
rect 51832 5502 51838 5794
rect 51872 5502 51878 5794
rect 51832 4700 51878 5502
rect 51832 4408 51838 4700
rect 51872 4408 51878 4700
rect 51832 3606 51878 4408
rect 51832 3576 51838 3606
rect 50814 3314 50852 3386
rect 50770 3248 50852 3314
rect 51872 3576 51878 3606
rect 52888 7690 52896 7790
rect 52930 7790 52998 7982
rect 54106 7996 54174 8070
rect 52930 7690 52934 7790
rect 52888 6888 52934 7690
rect 52888 6596 52896 6888
rect 52930 6596 52934 6888
rect 52888 5794 52934 6596
rect 54106 7704 54120 7996
rect 54154 7894 54174 7996
rect 55178 7996 55212 8012
rect 54106 7688 54154 7704
rect 55174 7704 55178 7902
rect 56210 7996 56278 8174
rect 56210 7908 56236 7996
rect 55212 7704 55220 7902
rect 54106 6918 54152 7688
rect 54106 6902 54154 6918
rect 54106 6610 54120 6902
rect 54106 6594 54154 6610
rect 55174 6902 55220 7704
rect 55174 6610 55178 6902
rect 55212 6610 55220 6902
rect 52888 5502 52896 5794
rect 52930 5502 52934 5794
rect 52888 4700 52934 5502
rect 53466 6462 53616 6588
rect 53466 5266 53488 6462
rect 53582 5266 53616 6462
rect 53466 4942 53616 5266
rect 54106 5824 54152 6594
rect 54106 5808 54154 5824
rect 54106 5516 54120 5808
rect 54106 5500 54154 5516
rect 55174 5808 55220 6610
rect 55174 5516 55178 5808
rect 55212 5516 55220 5808
rect 52888 4408 52896 4700
rect 52930 4408 52934 4700
rect 52888 3606 52934 4408
rect 52888 3548 52896 3606
rect 51838 3298 51872 3314
rect 52872 3314 52896 3408
rect 52930 3548 52934 3606
rect 54106 4730 54152 5500
rect 54106 4714 54154 4730
rect 54106 4422 54120 4714
rect 54106 4406 54154 4422
rect 55174 4714 55220 5516
rect 55174 4422 55178 4714
rect 55212 4422 55220 4714
rect 54106 3636 54152 4406
rect 54106 3620 54154 3636
rect 54106 3562 54120 3620
rect 52930 3314 52954 3408
rect 52872 3248 52954 3314
rect 55174 3620 55220 4422
rect 55174 3540 55178 3620
rect 54120 3312 54154 3328
rect 55158 3328 55178 3428
rect 55212 3540 55220 3620
rect 56226 7704 56236 7908
rect 56270 7960 56278 7996
rect 57294 7996 57328 8012
rect 56270 7908 56284 7960
rect 56270 7704 56272 7908
rect 56226 6902 56272 7704
rect 56226 6610 56236 6902
rect 56270 6610 56272 6902
rect 56226 5808 56272 6610
rect 56226 5516 56236 5808
rect 56270 5516 56272 5808
rect 56226 4714 56272 5516
rect 56226 4422 56236 4714
rect 56270 4422 56272 4714
rect 56226 3620 56272 4422
rect 56226 3562 56236 3620
rect 55212 3328 55240 3428
rect 55158 3248 55240 3328
rect 56270 3562 56272 3620
rect 58326 7996 58410 8184
rect 57328 7704 57340 7908
rect 58326 7904 58352 7996
rect 57294 6902 57340 7704
rect 57328 6610 57340 6902
rect 57294 5808 57340 6610
rect 57328 5516 57340 5808
rect 57294 4714 57340 5516
rect 57328 4422 57340 4714
rect 57294 3620 57340 4422
rect 56236 3312 56270 3328
rect 57284 3328 57294 3400
rect 57328 3546 57340 3620
rect 58346 7704 58352 7904
rect 58386 7904 58410 7996
rect 59368 7996 59494 9030
rect 63156 9004 67606 9094
rect 63168 8998 67606 9004
rect 69624 9092 69706 9202
rect 70736 9436 70738 9494
rect 72792 13870 72876 14058
rect 75122 14068 79556 14112
rect 81728 14120 81796 14130
rect 83832 14120 83900 14136
rect 85956 14120 86024 14152
rect 81728 14110 86024 14120
rect 75122 14032 79564 14068
rect 75122 14022 79412 14032
rect 71794 13578 71806 13782
rect 72792 13778 72818 13870
rect 71760 12776 71806 13578
rect 71794 12484 71806 12776
rect 71760 11682 71806 12484
rect 71794 11390 71806 11682
rect 71760 10588 71806 11390
rect 71794 10296 71806 10588
rect 71760 9494 71806 10296
rect 70702 9186 70736 9202
rect 71750 9202 71760 9274
rect 71794 9420 71806 9494
rect 72812 13578 72818 13778
rect 72852 13778 72876 13870
rect 73876 13870 73910 13886
rect 72852 13578 72858 13778
rect 72812 12776 72858 13578
rect 72812 12484 72818 12776
rect 72852 12484 72858 12776
rect 72812 11682 72858 12484
rect 72812 11390 72818 11682
rect 72852 11390 72858 11682
rect 72812 10588 72858 11390
rect 72812 10296 72818 10588
rect 72852 10296 72858 10588
rect 72812 9494 72858 10296
rect 72812 9464 72818 9494
rect 71794 9202 71832 9274
rect 71750 9092 71832 9202
rect 72852 9464 72858 9494
rect 73868 13578 73876 13798
rect 75260 13844 75328 14022
rect 73910 13578 73914 13798
rect 73868 12776 73914 13578
rect 73868 12484 73876 12776
rect 73910 12484 73914 12776
rect 73868 11682 73914 12484
rect 75260 13552 75274 13844
rect 75308 13742 75328 13844
rect 76332 13844 76366 13860
rect 75260 13536 75308 13552
rect 76328 13552 76332 13750
rect 77364 13844 77432 14022
rect 77364 13756 77390 13844
rect 76366 13552 76374 13750
rect 75260 12766 75306 13536
rect 75260 12750 75308 12766
rect 75260 12458 75274 12750
rect 75260 12442 75308 12458
rect 76328 12750 76374 13552
rect 76328 12458 76332 12750
rect 76366 12458 76374 12750
rect 73868 11390 73876 11682
rect 73910 11390 73914 11682
rect 73868 10588 73914 11390
rect 74620 12310 74770 12436
rect 74620 11114 74642 12310
rect 74736 11114 74770 12310
rect 74620 10790 74770 11114
rect 75260 11672 75306 12442
rect 75260 11656 75308 11672
rect 75260 11364 75274 11656
rect 75260 11348 75308 11364
rect 76328 11656 76374 12458
rect 76328 11364 76332 11656
rect 76366 11364 76374 11656
rect 73868 10296 73876 10588
rect 73910 10296 73914 10588
rect 73868 9494 73914 10296
rect 73868 9436 73876 9494
rect 72818 9186 72852 9202
rect 73852 9202 73876 9296
rect 73910 9436 73914 9494
rect 75260 10578 75306 11348
rect 75260 10562 75308 10578
rect 75260 10270 75274 10562
rect 75260 10254 75308 10270
rect 76328 10562 76374 11364
rect 76328 10270 76332 10562
rect 76366 10270 76374 10562
rect 75260 9484 75306 10254
rect 75260 9468 75308 9484
rect 75260 9410 75274 9468
rect 73910 9202 73934 9296
rect 73852 9092 73934 9202
rect 76328 9468 76374 10270
rect 76328 9388 76332 9468
rect 75274 9160 75308 9176
rect 76312 9176 76332 9276
rect 76366 9388 76374 9468
rect 77380 13552 77390 13756
rect 77424 13808 77432 13844
rect 78448 13844 78482 13860
rect 77424 13756 77438 13808
rect 77424 13552 77426 13756
rect 77380 12750 77426 13552
rect 77380 12458 77390 12750
rect 77424 12458 77426 12750
rect 77380 11656 77426 12458
rect 77380 11364 77390 11656
rect 77424 11364 77426 11656
rect 77380 10562 77426 11364
rect 77380 10270 77390 10562
rect 77424 10270 77426 10562
rect 77380 9468 77426 10270
rect 77380 9410 77390 9468
rect 76366 9176 76394 9276
rect 69624 9002 74074 9092
rect 65282 8976 65364 8998
rect 69636 8996 74074 9002
rect 76312 9066 76394 9176
rect 77424 9410 77426 9468
rect 79480 13844 79564 14032
rect 81590 14066 86024 14110
rect 88494 14114 88562 14124
rect 90598 14114 90666 14130
rect 92722 14114 92790 14146
rect 88494 14104 92790 14114
rect 81590 14030 86032 14066
rect 81590 14020 85880 14030
rect 78482 13552 78494 13756
rect 79480 13752 79506 13844
rect 78448 12750 78494 13552
rect 78482 12458 78494 12750
rect 78448 11656 78494 12458
rect 78482 11364 78494 11656
rect 78448 10562 78494 11364
rect 78482 10270 78494 10562
rect 78448 9468 78494 10270
rect 77390 9160 77424 9176
rect 78438 9176 78448 9248
rect 78482 9394 78494 9468
rect 79500 13552 79506 13752
rect 79540 13752 79564 13844
rect 80564 13844 80598 13860
rect 79540 13552 79546 13752
rect 79500 12750 79546 13552
rect 79500 12458 79506 12750
rect 79540 12458 79546 12750
rect 79500 11656 79546 12458
rect 79500 11364 79506 11656
rect 79540 11364 79546 11656
rect 79500 10562 79546 11364
rect 79500 10270 79506 10562
rect 79540 10270 79546 10562
rect 79500 9468 79546 10270
rect 79500 9438 79506 9468
rect 78482 9176 78520 9248
rect 78438 9066 78520 9176
rect 79540 9438 79546 9468
rect 80556 13552 80564 13772
rect 81728 13842 81796 14020
rect 80598 13552 80602 13772
rect 80556 12750 80602 13552
rect 80556 12458 80564 12750
rect 80598 12458 80602 12750
rect 80556 11656 80602 12458
rect 81728 13550 81742 13842
rect 81776 13740 81796 13842
rect 82800 13842 82834 13858
rect 81728 13534 81776 13550
rect 82796 13550 82800 13748
rect 83832 13842 83900 14020
rect 83832 13754 83858 13842
rect 82834 13550 82842 13748
rect 81728 12764 81774 13534
rect 81728 12748 81776 12764
rect 81728 12456 81742 12748
rect 81728 12440 81776 12456
rect 82796 12748 82842 13550
rect 82796 12456 82800 12748
rect 82834 12456 82842 12748
rect 80556 11364 80564 11656
rect 80598 11364 80602 11656
rect 80556 10562 80602 11364
rect 81088 12308 81238 12434
rect 81088 11112 81110 12308
rect 81204 11112 81238 12308
rect 81088 10788 81238 11112
rect 81728 11670 81774 12440
rect 81728 11654 81776 11670
rect 81728 11362 81742 11654
rect 81728 11346 81776 11362
rect 82796 11654 82842 12456
rect 82796 11362 82800 11654
rect 82834 11362 82842 11654
rect 80556 10270 80564 10562
rect 80598 10270 80602 10562
rect 80556 9468 80602 10270
rect 80556 9410 80564 9468
rect 79506 9160 79540 9176
rect 80540 9176 80564 9270
rect 80598 9410 80602 9468
rect 81728 10576 81774 11346
rect 81728 10560 81776 10576
rect 81728 10268 81742 10560
rect 81728 10252 81776 10268
rect 82796 10560 82842 11362
rect 82796 10268 82800 10560
rect 82834 10268 82842 10560
rect 81728 9482 81774 10252
rect 81728 9466 81776 9482
rect 81728 9408 81742 9466
rect 80598 9176 80622 9270
rect 80540 9066 80622 9176
rect 82796 9466 82842 10268
rect 82796 9386 82800 9466
rect 81742 9158 81776 9174
rect 82780 9174 82800 9274
rect 82834 9386 82842 9466
rect 83848 13550 83858 13754
rect 83892 13806 83900 13842
rect 84916 13842 84950 13858
rect 83892 13754 83906 13806
rect 83892 13550 83894 13754
rect 83848 12748 83894 13550
rect 83848 12456 83858 12748
rect 83892 12456 83894 12748
rect 83848 11654 83894 12456
rect 83848 11362 83858 11654
rect 83892 11362 83894 11654
rect 83848 10560 83894 11362
rect 83848 10268 83858 10560
rect 83892 10268 83894 10560
rect 83848 9466 83894 10268
rect 83848 9408 83858 9466
rect 82834 9174 82862 9274
rect 71750 8974 71832 8996
rect 76312 8976 80762 9066
rect 76324 8970 80762 8976
rect 82780 9064 82862 9174
rect 83892 9408 83894 9466
rect 85948 13842 86032 14030
rect 88356 14060 92790 14104
rect 94962 14112 95030 14122
rect 97066 14112 97134 14128
rect 99190 14112 99258 14144
rect 94962 14102 99258 14112
rect 88356 14024 92798 14060
rect 88356 14014 92646 14024
rect 84950 13550 84962 13754
rect 85948 13750 85974 13842
rect 84916 12748 84962 13550
rect 84950 12456 84962 12748
rect 84916 11654 84962 12456
rect 84950 11362 84962 11654
rect 84916 10560 84962 11362
rect 84950 10268 84962 10560
rect 84916 9466 84962 10268
rect 83858 9158 83892 9174
rect 84906 9174 84916 9246
rect 84950 9392 84962 9466
rect 85968 13550 85974 13750
rect 86008 13750 86032 13842
rect 87032 13842 87066 13858
rect 86008 13550 86014 13750
rect 85968 12748 86014 13550
rect 85968 12456 85974 12748
rect 86008 12456 86014 12748
rect 85968 11654 86014 12456
rect 85968 11362 85974 11654
rect 86008 11362 86014 11654
rect 85968 10560 86014 11362
rect 85968 10268 85974 10560
rect 86008 10268 86014 10560
rect 85968 9466 86014 10268
rect 85968 9436 85974 9466
rect 84950 9174 84988 9246
rect 84906 9064 84988 9174
rect 86008 9436 86014 9466
rect 87024 13550 87032 13770
rect 88494 13836 88562 14014
rect 87066 13550 87070 13770
rect 87024 12748 87070 13550
rect 87024 12456 87032 12748
rect 87066 12456 87070 12748
rect 87024 11654 87070 12456
rect 88494 13544 88508 13836
rect 88542 13734 88562 13836
rect 89566 13836 89600 13852
rect 88494 13528 88542 13544
rect 89562 13544 89566 13742
rect 90598 13836 90666 14014
rect 90598 13748 90624 13836
rect 89600 13544 89608 13742
rect 88494 12758 88540 13528
rect 88494 12742 88542 12758
rect 88494 12450 88508 12742
rect 88494 12434 88542 12450
rect 89562 12742 89608 13544
rect 89562 12450 89566 12742
rect 89600 12450 89608 12742
rect 87024 11362 87032 11654
rect 87066 11362 87070 11654
rect 87024 10560 87070 11362
rect 87854 12302 88004 12428
rect 87854 11106 87876 12302
rect 87970 11106 88004 12302
rect 87854 10782 88004 11106
rect 88494 11664 88540 12434
rect 88494 11648 88542 11664
rect 88494 11356 88508 11648
rect 88494 11340 88542 11356
rect 89562 11648 89608 12450
rect 89562 11356 89566 11648
rect 89600 11356 89608 11648
rect 87024 10268 87032 10560
rect 87066 10268 87070 10560
rect 87024 9466 87070 10268
rect 87024 9408 87032 9466
rect 85974 9158 86008 9174
rect 87008 9174 87032 9268
rect 87066 9408 87070 9466
rect 88494 10570 88540 11340
rect 88494 10554 88542 10570
rect 88494 10262 88508 10554
rect 88494 10246 88542 10262
rect 89562 10554 89608 11356
rect 89562 10262 89566 10554
rect 89600 10262 89608 10554
rect 88494 9476 88540 10246
rect 88494 9460 88542 9476
rect 88494 9402 88508 9460
rect 87066 9174 87090 9268
rect 87008 9064 87090 9174
rect 89562 9460 89608 10262
rect 89562 9380 89566 9460
rect 88508 9152 88542 9168
rect 89546 9168 89566 9268
rect 89600 9380 89608 9460
rect 90614 13544 90624 13748
rect 90658 13800 90666 13836
rect 91682 13836 91716 13852
rect 90658 13748 90672 13800
rect 90658 13544 90660 13748
rect 90614 12742 90660 13544
rect 90614 12450 90624 12742
rect 90658 12450 90660 12742
rect 90614 11648 90660 12450
rect 90614 11356 90624 11648
rect 90658 11356 90660 11648
rect 90614 10554 90660 11356
rect 90614 10262 90624 10554
rect 90658 10262 90660 10554
rect 90614 9460 90660 10262
rect 90614 9402 90624 9460
rect 89600 9168 89628 9268
rect 82780 8974 87230 9064
rect 78438 8948 78520 8970
rect 82792 8968 87230 8974
rect 89546 9058 89628 9168
rect 90658 9402 90660 9460
rect 92714 13836 92798 14024
rect 94824 14058 99258 14102
rect 94824 14022 99266 14058
rect 94824 14012 99114 14022
rect 91716 13544 91728 13748
rect 92714 13744 92740 13836
rect 91682 12742 91728 13544
rect 91716 12450 91728 12742
rect 91682 11648 91728 12450
rect 91716 11356 91728 11648
rect 91682 10554 91728 11356
rect 91716 10262 91728 10554
rect 91682 9460 91728 10262
rect 90624 9152 90658 9168
rect 91672 9168 91682 9240
rect 91716 9386 91728 9460
rect 92734 13544 92740 13744
rect 92774 13744 92798 13836
rect 93798 13836 93832 13852
rect 92774 13544 92780 13744
rect 92734 12742 92780 13544
rect 92734 12450 92740 12742
rect 92774 12450 92780 12742
rect 92734 11648 92780 12450
rect 92734 11356 92740 11648
rect 92774 11356 92780 11648
rect 92734 10554 92780 11356
rect 92734 10262 92740 10554
rect 92774 10262 92780 10554
rect 92734 9460 92780 10262
rect 92734 9430 92740 9460
rect 91716 9168 91754 9240
rect 91672 9058 91754 9168
rect 92774 9430 92780 9460
rect 93790 13544 93798 13764
rect 94962 13834 95030 14012
rect 93832 13544 93836 13764
rect 93790 12742 93836 13544
rect 93790 12450 93798 12742
rect 93832 12450 93836 12742
rect 93790 11648 93836 12450
rect 94962 13542 94976 13834
rect 95010 13732 95030 13834
rect 96034 13834 96068 13850
rect 94962 13526 95010 13542
rect 96030 13542 96034 13740
rect 97066 13834 97134 14012
rect 97066 13746 97092 13834
rect 96068 13542 96076 13740
rect 94962 12756 95008 13526
rect 94962 12740 95010 12756
rect 94962 12448 94976 12740
rect 94962 12432 95010 12448
rect 96030 12740 96076 13542
rect 96030 12448 96034 12740
rect 96068 12448 96076 12740
rect 93790 11356 93798 11648
rect 93832 11356 93836 11648
rect 93790 10554 93836 11356
rect 94322 12300 94472 12426
rect 94322 11104 94344 12300
rect 94438 11104 94472 12300
rect 94322 10780 94472 11104
rect 94962 11662 95008 12432
rect 94962 11646 95010 11662
rect 94962 11354 94976 11646
rect 94962 11338 95010 11354
rect 96030 11646 96076 12448
rect 96030 11354 96034 11646
rect 96068 11354 96076 11646
rect 93790 10262 93798 10554
rect 93832 10262 93836 10554
rect 93790 9460 93836 10262
rect 93790 9402 93798 9460
rect 92740 9152 92774 9168
rect 93774 9168 93798 9262
rect 93832 9402 93836 9460
rect 94962 10568 95008 11338
rect 94962 10552 95010 10568
rect 94962 10260 94976 10552
rect 94962 10244 95010 10260
rect 96030 10552 96076 11354
rect 96030 10260 96034 10552
rect 96068 10260 96076 10552
rect 94962 9474 95008 10244
rect 94962 9458 95010 9474
rect 94962 9400 94976 9458
rect 93832 9168 93856 9262
rect 93774 9058 93856 9168
rect 96030 9458 96076 10260
rect 96030 9378 96034 9458
rect 94976 9150 95010 9166
rect 96014 9166 96034 9266
rect 96068 9378 96076 9458
rect 97082 13542 97092 13746
rect 97126 13798 97134 13834
rect 98150 13834 98184 13850
rect 97126 13746 97140 13798
rect 97126 13542 97128 13746
rect 97082 12740 97128 13542
rect 97082 12448 97092 12740
rect 97126 12448 97128 12740
rect 97082 11646 97128 12448
rect 97082 11354 97092 11646
rect 97126 11354 97128 11646
rect 97082 10552 97128 11354
rect 97082 10260 97092 10552
rect 97126 10260 97128 10552
rect 97082 9458 97128 10260
rect 97082 9400 97092 9458
rect 96068 9166 96096 9266
rect 89546 8968 93996 9058
rect 84906 8946 84988 8968
rect 89558 8962 93996 8968
rect 96014 9056 96096 9166
rect 97126 9400 97128 9458
rect 99182 13834 99266 14022
rect 98184 13542 98196 13746
rect 99182 13742 99208 13834
rect 98150 12740 98196 13542
rect 98184 12448 98196 12740
rect 98150 11646 98196 12448
rect 98184 11354 98196 11646
rect 98150 10552 98196 11354
rect 98184 10260 98196 10552
rect 98150 9458 98196 10260
rect 97092 9150 97126 9166
rect 98140 9166 98150 9238
rect 98184 9384 98196 9458
rect 99202 13542 99208 13742
rect 99242 13742 99266 13834
rect 100266 13834 100300 13850
rect 99242 13542 99248 13742
rect 99202 12740 99248 13542
rect 99202 12448 99208 12740
rect 99242 12448 99248 12740
rect 99202 11646 99248 12448
rect 99202 11354 99208 11646
rect 99242 11354 99248 11646
rect 99202 10552 99248 11354
rect 99202 10260 99208 10552
rect 99242 10260 99248 10552
rect 99202 9458 99248 10260
rect 99202 9428 99208 9458
rect 98184 9166 98222 9238
rect 98140 9056 98222 9166
rect 99242 9428 99248 9458
rect 100258 13542 100266 13762
rect 100300 13542 100304 13762
rect 100258 12740 100304 13542
rect 100258 12448 100266 12740
rect 100300 12448 100304 12740
rect 100258 11646 100304 12448
rect 100258 11354 100266 11646
rect 100300 11354 100304 11646
rect 100258 10552 100304 11354
rect 100258 10260 100266 10552
rect 100300 10260 100304 10552
rect 100258 9458 100304 10260
rect 100258 9400 100266 9458
rect 99208 9150 99242 9166
rect 100242 9166 100266 9260
rect 100300 9400 100304 9458
rect 100630 13700 101298 13902
rect 100630 9516 100742 13700
rect 101232 9516 101298 13700
rect 100630 9294 101298 9516
rect 100300 9166 100324 9260
rect 100242 9056 100324 9166
rect 96014 8966 100464 9056
rect 91672 8940 91754 8962
rect 96026 8960 100464 8966
rect 98140 8938 98222 8960
rect 62104 8292 62172 8302
rect 64208 8292 64276 8308
rect 66332 8292 66400 8324
rect 62104 8282 66400 8292
rect 61966 8238 66400 8282
rect 68576 8290 68644 8300
rect 70680 8290 70748 8306
rect 72804 8290 72872 8322
rect 68576 8280 72872 8290
rect 61966 8202 66408 8238
rect 61966 8192 66256 8202
rect 58386 7704 58392 7904
rect 59368 7832 59410 7996
rect 58346 6902 58392 7704
rect 58346 6610 58352 6902
rect 58386 6610 58392 6902
rect 58346 5808 58392 6610
rect 58346 5516 58352 5808
rect 58386 5516 58392 5808
rect 58346 4714 58392 5516
rect 58346 4422 58352 4714
rect 58386 4422 58392 4714
rect 58346 3620 58392 4422
rect 58346 3590 58352 3620
rect 57328 3328 57366 3400
rect 46284 3218 56720 3248
rect 57284 3218 57366 3328
rect 58386 3590 58392 3620
rect 59402 7704 59410 7832
rect 59444 7832 59494 7996
rect 62104 8014 62172 8192
rect 59444 7704 59448 7832
rect 59402 6902 59448 7704
rect 59402 6610 59410 6902
rect 59444 6610 59448 6902
rect 62104 7722 62118 8014
rect 62152 7912 62172 8014
rect 63176 8014 63210 8030
rect 62104 7706 62152 7722
rect 63172 7722 63176 7920
rect 64208 8014 64276 8192
rect 64208 7926 64234 8014
rect 63210 7722 63218 7920
rect 62104 6936 62150 7706
rect 62104 6920 62152 6936
rect 59402 5808 59448 6610
rect 59402 5516 59410 5808
rect 59444 5516 59448 5808
rect 59402 4714 59448 5516
rect 59600 6714 59948 6812
rect 59600 5340 59684 6714
rect 59850 5936 59948 6714
rect 62104 6628 62118 6920
rect 62104 6612 62152 6628
rect 63172 6920 63218 7722
rect 63172 6628 63176 6920
rect 63210 6628 63218 6920
rect 61464 6480 61614 6606
rect 59850 5340 60160 5936
rect 59600 5174 60160 5340
rect 59402 4422 59410 4714
rect 59444 4422 59448 4714
rect 59402 3620 59448 4422
rect 59402 3562 59410 3620
rect 58352 3312 58386 3328
rect 59386 3328 59410 3422
rect 59444 3562 59448 3620
rect 59444 3328 59468 3422
rect 59386 3218 59468 3328
rect 46284 3182 59608 3218
rect 42056 3122 59608 3182
rect 42056 3092 56720 3122
rect 57284 3100 57366 3122
rect 42068 3086 56720 3092
rect 44182 3064 44264 3086
rect 46354 3042 56720 3086
rect 59718 -184 60160 5174
rect 61464 5284 61486 6480
rect 61580 5284 61614 6480
rect 61464 4960 61614 5284
rect 62104 5842 62150 6612
rect 62104 5826 62152 5842
rect 62104 5534 62118 5826
rect 62104 5518 62152 5534
rect 63172 5826 63218 6628
rect 63172 5534 63176 5826
rect 63210 5534 63218 5826
rect 62104 4748 62150 5518
rect 62104 4732 62152 4748
rect 62104 4440 62118 4732
rect 62104 4424 62152 4440
rect 63172 4732 63218 5534
rect 63172 4440 63176 4732
rect 63210 4440 63218 4732
rect 62104 3654 62150 4424
rect 62104 3638 62152 3654
rect 62104 3580 62118 3638
rect 63172 3638 63218 4440
rect 63172 3558 63176 3638
rect 62118 3330 62152 3346
rect 63156 3346 63176 3446
rect 63210 3558 63218 3638
rect 64224 7722 64234 7926
rect 64268 7978 64276 8014
rect 65292 8014 65326 8030
rect 64268 7926 64282 7978
rect 64268 7722 64270 7926
rect 64224 6920 64270 7722
rect 64224 6628 64234 6920
rect 64268 6628 64270 6920
rect 64224 5826 64270 6628
rect 64224 5534 64234 5826
rect 64268 5534 64270 5826
rect 64224 4732 64270 5534
rect 64224 4440 64234 4732
rect 64268 4440 64270 4732
rect 64224 3638 64270 4440
rect 64224 3580 64234 3638
rect 63210 3346 63238 3446
rect 63156 3236 63238 3346
rect 64268 3580 64270 3638
rect 66324 8014 66408 8202
rect 68438 8236 72872 8280
rect 75260 8264 75328 8274
rect 77364 8264 77432 8280
rect 79488 8264 79556 8296
rect 75260 8254 79556 8264
rect 68438 8200 72880 8236
rect 68438 8190 72728 8200
rect 65326 7722 65338 7926
rect 66324 7922 66350 8014
rect 65292 6920 65338 7722
rect 65326 6628 65338 6920
rect 65292 5826 65338 6628
rect 65326 5534 65338 5826
rect 65292 4732 65338 5534
rect 65326 4440 65338 4732
rect 65292 3638 65338 4440
rect 64234 3330 64268 3346
rect 65282 3346 65292 3418
rect 65326 3564 65338 3638
rect 66344 7722 66350 7922
rect 66384 7922 66408 8014
rect 67408 8014 67442 8030
rect 66384 7722 66390 7922
rect 66344 6920 66390 7722
rect 66344 6628 66350 6920
rect 66384 6628 66390 6920
rect 66344 5826 66390 6628
rect 66344 5534 66350 5826
rect 66384 5534 66390 5826
rect 66344 4732 66390 5534
rect 66344 4440 66350 4732
rect 66384 4440 66390 4732
rect 66344 3638 66390 4440
rect 66344 3608 66350 3638
rect 65326 3346 65364 3418
rect 65282 3236 65364 3346
rect 66384 3608 66390 3638
rect 67400 7722 67408 7942
rect 68576 8012 68644 8190
rect 67442 7722 67446 7942
rect 67400 6920 67446 7722
rect 67400 6628 67408 6920
rect 67442 6628 67446 6920
rect 67400 5826 67446 6628
rect 68576 7720 68590 8012
rect 68624 7910 68644 8012
rect 69648 8012 69682 8028
rect 68576 7704 68624 7720
rect 69644 7720 69648 7918
rect 70680 8012 70748 8190
rect 70680 7924 70706 8012
rect 69682 7720 69690 7918
rect 68576 6934 68622 7704
rect 68576 6918 68624 6934
rect 68576 6626 68590 6918
rect 68576 6610 68624 6626
rect 69644 6918 69690 7720
rect 69644 6626 69648 6918
rect 69682 6626 69690 6918
rect 67400 5534 67408 5826
rect 67442 5534 67446 5826
rect 67936 6478 68086 6604
rect 67936 5814 67958 6478
rect 67400 4732 67446 5534
rect 67400 4440 67408 4732
rect 67442 4440 67446 4732
rect 67400 3638 67446 4440
rect 67400 3580 67408 3638
rect 66350 3330 66384 3346
rect 67384 3346 67408 3440
rect 67442 3580 67446 3638
rect 67706 5282 67958 5814
rect 68052 5814 68086 6478
rect 68576 5840 68622 6610
rect 68576 5824 68624 5840
rect 68052 5282 68258 5814
rect 67442 3346 67466 3440
rect 67384 3242 67466 3346
rect 67706 3242 68258 5282
rect 68576 5532 68590 5824
rect 68576 5516 68624 5532
rect 69644 5824 69690 6626
rect 69644 5532 69648 5824
rect 69682 5532 69690 5824
rect 68576 4746 68622 5516
rect 68576 4730 68624 4746
rect 68576 4438 68590 4730
rect 68576 4422 68624 4438
rect 69644 4730 69690 5532
rect 69644 4438 69648 4730
rect 69682 4438 69690 4730
rect 68576 3652 68622 4422
rect 68576 3636 68624 3652
rect 68576 3578 68590 3636
rect 69644 3636 69690 4438
rect 69644 3556 69648 3636
rect 68590 3328 68624 3344
rect 69628 3344 69648 3444
rect 69682 3556 69690 3636
rect 70696 7720 70706 7924
rect 70740 7976 70748 8012
rect 71764 8012 71798 8028
rect 70740 7924 70754 7976
rect 70740 7720 70742 7924
rect 70696 6918 70742 7720
rect 70696 6626 70706 6918
rect 70740 6626 70742 6918
rect 70696 5824 70742 6626
rect 70696 5532 70706 5824
rect 70740 5532 70742 5824
rect 70696 4730 70742 5532
rect 70696 4438 70706 4730
rect 70740 4438 70742 4730
rect 70696 3636 70742 4438
rect 70696 3578 70706 3636
rect 69682 3344 69710 3444
rect 69628 3242 69710 3344
rect 70740 3578 70742 3636
rect 72796 8012 72880 8200
rect 75122 8210 79556 8254
rect 81732 8262 81800 8272
rect 83836 8262 83904 8278
rect 85960 8262 86028 8294
rect 81732 8252 86028 8262
rect 75122 8174 79564 8210
rect 75122 8164 79412 8174
rect 71798 7720 71810 7924
rect 72796 7920 72822 8012
rect 71764 6918 71810 7720
rect 71798 6626 71810 6918
rect 71764 5824 71810 6626
rect 71798 5532 71810 5824
rect 71764 4730 71810 5532
rect 71798 4438 71810 4730
rect 71764 3636 71810 4438
rect 70706 3328 70740 3344
rect 71754 3344 71764 3416
rect 71798 3562 71810 3636
rect 72816 7720 72822 7920
rect 72856 7920 72880 8012
rect 73880 8012 73914 8028
rect 72856 7720 72862 7920
rect 72816 6918 72862 7720
rect 72816 6626 72822 6918
rect 72856 6626 72862 6918
rect 72816 5824 72862 6626
rect 72816 5532 72822 5824
rect 72856 5532 72862 5824
rect 72816 4730 72862 5532
rect 72816 4438 72822 4730
rect 72856 4438 72862 4730
rect 72816 3636 72862 4438
rect 72816 3606 72822 3636
rect 71798 3344 71836 3416
rect 67384 3236 69740 3242
rect 63156 3234 69740 3236
rect 71754 3234 71836 3344
rect 72856 3606 72862 3636
rect 73872 7720 73880 7940
rect 75260 7986 75328 8164
rect 73914 7720 73918 7940
rect 73872 6918 73918 7720
rect 73872 6626 73880 6918
rect 73914 6626 73918 6918
rect 73872 5824 73918 6626
rect 75260 7694 75274 7986
rect 75308 7884 75328 7986
rect 76332 7986 76366 8002
rect 75260 7678 75308 7694
rect 76328 7694 76332 7892
rect 77364 7986 77432 8164
rect 77364 7898 77390 7986
rect 76366 7694 76374 7892
rect 75260 6908 75306 7678
rect 75260 6892 75308 6908
rect 75260 6600 75274 6892
rect 75260 6584 75308 6600
rect 76328 6892 76374 7694
rect 76328 6600 76332 6892
rect 76366 6600 76374 6892
rect 74620 6452 74770 6578
rect 74620 5924 74642 6452
rect 73872 5532 73880 5824
rect 73914 5532 73918 5824
rect 73872 4730 73918 5532
rect 73872 4438 73880 4730
rect 73914 4438 73918 4730
rect 73872 3636 73918 4438
rect 73872 3578 73880 3636
rect 72822 3328 72856 3344
rect 73856 3344 73880 3438
rect 73914 3578 73918 3636
rect 74412 5256 74642 5924
rect 74736 5924 74770 6452
rect 74736 5256 74964 5924
rect 73914 3344 73938 3438
rect 73856 3234 73938 3344
rect 63156 3146 74078 3234
rect 63168 3140 74078 3146
rect 65282 3118 65364 3140
rect 67418 3138 74078 3140
rect 67418 3132 69740 3138
rect 67706 840 68258 3132
rect 71754 3116 71836 3138
rect 74412 804 74964 5256
rect 75260 5814 75306 6584
rect 75260 5798 75308 5814
rect 75260 5506 75274 5798
rect 75260 5490 75308 5506
rect 76328 5798 76374 6600
rect 76328 5506 76332 5798
rect 76366 5506 76374 5798
rect 75260 4720 75306 5490
rect 75260 4704 75308 4720
rect 75260 4412 75274 4704
rect 75260 4396 75308 4412
rect 76328 4704 76374 5506
rect 76328 4412 76332 4704
rect 76366 4412 76374 4704
rect 75260 3626 75306 4396
rect 75260 3610 75308 3626
rect 75260 3552 75274 3610
rect 76328 3610 76374 4412
rect 76328 3530 76332 3610
rect 75274 3302 75308 3318
rect 76312 3318 76332 3418
rect 76366 3530 76374 3610
rect 77380 7694 77390 7898
rect 77424 7950 77432 7986
rect 78448 7986 78482 8002
rect 77424 7898 77438 7950
rect 77424 7694 77426 7898
rect 77380 6892 77426 7694
rect 77380 6600 77390 6892
rect 77424 6600 77426 6892
rect 77380 5798 77426 6600
rect 77380 5506 77390 5798
rect 77424 5506 77426 5798
rect 77380 4704 77426 5506
rect 77380 4412 77390 4704
rect 77424 4412 77426 4704
rect 77380 3610 77426 4412
rect 77380 3552 77390 3610
rect 76366 3318 76394 3418
rect 76312 3208 76394 3318
rect 77424 3552 77426 3610
rect 79480 7986 79564 8174
rect 81594 8208 86028 8252
rect 88494 8256 88562 8266
rect 90598 8256 90666 8272
rect 92722 8256 92790 8288
rect 88494 8246 92790 8256
rect 81594 8172 86036 8208
rect 81594 8162 85884 8172
rect 78482 7694 78494 7898
rect 79480 7894 79506 7986
rect 78448 6892 78494 7694
rect 78482 6600 78494 6892
rect 78448 5798 78494 6600
rect 78482 5506 78494 5798
rect 78448 4704 78494 5506
rect 78482 4412 78494 4704
rect 78448 3610 78494 4412
rect 77390 3302 77424 3318
rect 78438 3318 78448 3390
rect 78482 3536 78494 3610
rect 79500 7694 79506 7894
rect 79540 7894 79564 7986
rect 80564 7986 80598 8002
rect 79540 7694 79546 7894
rect 79500 6892 79546 7694
rect 79500 6600 79506 6892
rect 79540 6600 79546 6892
rect 79500 5798 79546 6600
rect 79500 5506 79506 5798
rect 79540 5506 79546 5798
rect 79500 4704 79546 5506
rect 79500 4412 79506 4704
rect 79540 4412 79546 4704
rect 79500 3610 79546 4412
rect 79500 3580 79506 3610
rect 78482 3318 78520 3390
rect 78438 3208 78520 3318
rect 79540 3580 79546 3610
rect 80556 7694 80564 7914
rect 81732 7984 81800 8162
rect 80598 7694 80602 7914
rect 80556 6892 80602 7694
rect 80556 6600 80564 6892
rect 80598 6600 80602 6892
rect 80556 5798 80602 6600
rect 81732 7692 81746 7984
rect 81780 7882 81800 7984
rect 82804 7984 82838 8000
rect 81732 7676 81780 7692
rect 82800 7692 82804 7890
rect 83836 7984 83904 8162
rect 83836 7896 83862 7984
rect 82838 7692 82846 7890
rect 81732 6906 81778 7676
rect 81732 6890 81780 6906
rect 81732 6598 81746 6890
rect 81732 6582 81780 6598
rect 82800 6890 82846 7692
rect 82800 6598 82804 6890
rect 82838 6598 82846 6890
rect 80556 5506 80564 5798
rect 80598 5506 80602 5798
rect 80556 4704 80602 5506
rect 81092 6450 81242 6576
rect 81092 5254 81114 6450
rect 81208 5254 81242 6450
rect 81092 4930 81242 5254
rect 81732 5812 81778 6582
rect 81732 5796 81780 5812
rect 81732 5504 81746 5796
rect 81732 5488 81780 5504
rect 82800 5796 82846 6598
rect 82800 5504 82804 5796
rect 82838 5504 82846 5796
rect 80556 4412 80564 4704
rect 80598 4412 80602 4704
rect 80556 3610 80602 4412
rect 80556 3552 80564 3610
rect 79506 3302 79540 3318
rect 80540 3318 80564 3412
rect 80598 3552 80602 3610
rect 81732 4718 81778 5488
rect 81732 4702 81780 4718
rect 81732 4410 81746 4702
rect 81732 4394 81780 4410
rect 82800 4702 82846 5504
rect 82800 4410 82804 4702
rect 82838 4410 82846 4702
rect 81732 3624 81778 4394
rect 81732 3608 81780 3624
rect 81732 3550 81746 3608
rect 80598 3318 80622 3412
rect 80540 3214 80622 3318
rect 82800 3608 82846 4410
rect 82800 3528 82804 3608
rect 81746 3300 81780 3316
rect 82784 3316 82804 3416
rect 82838 3528 82846 3608
rect 83852 7692 83862 7896
rect 83896 7948 83904 7984
rect 84920 7984 84954 8000
rect 83896 7896 83910 7948
rect 83896 7692 83898 7896
rect 83852 6890 83898 7692
rect 83852 6598 83862 6890
rect 83896 6598 83898 6890
rect 83852 5796 83898 6598
rect 83852 5504 83862 5796
rect 83896 5504 83898 5796
rect 83852 4702 83898 5504
rect 83852 4410 83862 4702
rect 83896 4410 83898 4702
rect 83852 3608 83898 4410
rect 83852 3550 83862 3608
rect 82838 3316 82866 3416
rect 82784 3214 82866 3316
rect 83896 3550 83898 3608
rect 85952 7984 86036 8172
rect 88356 8202 92790 8246
rect 94966 8254 95034 8264
rect 97070 8254 97138 8270
rect 99194 8254 99262 8286
rect 94966 8244 99262 8254
rect 88356 8166 92798 8202
rect 88356 8156 92646 8166
rect 84954 7692 84966 7896
rect 85952 7892 85978 7984
rect 84920 6890 84966 7692
rect 84954 6598 84966 6890
rect 84920 5796 84966 6598
rect 84954 5504 84966 5796
rect 84920 4702 84966 5504
rect 84954 4410 84966 4702
rect 84920 3608 84966 4410
rect 83862 3300 83896 3316
rect 84910 3316 84920 3388
rect 84954 3534 84966 3608
rect 85972 7692 85978 7892
rect 86012 7892 86036 7984
rect 87036 7984 87070 8000
rect 86012 7692 86018 7892
rect 85972 6890 86018 7692
rect 85972 6598 85978 6890
rect 86012 6598 86018 6890
rect 85972 5796 86018 6598
rect 85972 5504 85978 5796
rect 86012 5504 86018 5796
rect 85972 4702 86018 5504
rect 85972 4410 85978 4702
rect 86012 4410 86018 4702
rect 85972 3608 86018 4410
rect 85972 3578 85978 3608
rect 84954 3316 84992 3388
rect 80540 3208 82896 3214
rect 76312 3206 82896 3208
rect 84910 3206 84992 3316
rect 86012 3578 86018 3608
rect 87028 7692 87036 7912
rect 88494 7978 88562 8156
rect 87070 7692 87074 7912
rect 87028 6890 87074 7692
rect 87028 6598 87036 6890
rect 87070 6598 87074 6890
rect 87028 5796 87074 6598
rect 88494 7686 88508 7978
rect 88542 7876 88562 7978
rect 89566 7978 89600 7994
rect 88494 7670 88542 7686
rect 89562 7686 89566 7884
rect 90598 7978 90666 8156
rect 90598 7890 90624 7978
rect 89600 7686 89608 7884
rect 88494 6900 88540 7670
rect 88494 6884 88542 6900
rect 88494 6592 88508 6884
rect 88494 6576 88542 6592
rect 89562 6884 89608 7686
rect 89562 6592 89566 6884
rect 89600 6592 89608 6884
rect 87028 5504 87036 5796
rect 87070 5504 87074 5796
rect 87028 4702 87074 5504
rect 87854 6444 88004 6570
rect 87854 5248 87876 6444
rect 87970 5248 88004 6444
rect 87854 4924 88004 5248
rect 88494 5806 88540 6576
rect 88494 5790 88542 5806
rect 88494 5498 88508 5790
rect 88494 5482 88542 5498
rect 89562 5790 89608 6592
rect 89562 5498 89566 5790
rect 89600 5498 89608 5790
rect 87028 4410 87036 4702
rect 87070 4410 87074 4702
rect 87028 3608 87074 4410
rect 87028 3550 87036 3608
rect 85978 3300 86012 3316
rect 87012 3316 87036 3410
rect 87070 3550 87074 3608
rect 88494 4712 88540 5482
rect 88494 4696 88542 4712
rect 88494 4404 88508 4696
rect 88494 4388 88542 4404
rect 89562 4696 89608 5498
rect 89562 4404 89566 4696
rect 89600 4404 89608 4696
rect 88494 3618 88540 4388
rect 88494 3602 88542 3618
rect 88494 3544 88508 3602
rect 87070 3316 87094 3410
rect 87012 3206 87094 3316
rect 89562 3602 89608 4404
rect 89562 3522 89566 3602
rect 88508 3294 88542 3310
rect 89546 3310 89566 3410
rect 89600 3522 89608 3602
rect 90614 7686 90624 7890
rect 90658 7942 90666 7978
rect 91682 7978 91716 7994
rect 90658 7890 90672 7942
rect 90658 7686 90660 7890
rect 90614 6884 90660 7686
rect 90614 6592 90624 6884
rect 90658 6592 90660 6884
rect 90614 5790 90660 6592
rect 90614 5498 90624 5790
rect 90658 5498 90660 5790
rect 90614 4696 90660 5498
rect 90614 4404 90624 4696
rect 90658 4404 90660 4696
rect 90614 3602 90660 4404
rect 90614 3544 90624 3602
rect 89600 3310 89628 3410
rect 76312 3118 87234 3206
rect 76324 3112 87234 3118
rect 78438 3090 78520 3112
rect 80574 3110 87234 3112
rect 89546 3200 89628 3310
rect 90658 3544 90660 3602
rect 92714 7978 92798 8166
rect 94828 8200 99262 8244
rect 94828 8164 99270 8200
rect 94828 8154 99118 8164
rect 91716 7686 91728 7890
rect 92714 7886 92740 7978
rect 91682 6884 91728 7686
rect 91716 6592 91728 6884
rect 91682 5790 91728 6592
rect 91716 5498 91728 5790
rect 91682 4696 91728 5498
rect 91716 4404 91728 4696
rect 91682 3602 91728 4404
rect 90624 3294 90658 3310
rect 91672 3310 91682 3382
rect 91716 3528 91728 3602
rect 92734 7686 92740 7886
rect 92774 7886 92798 7978
rect 93798 7978 93832 7994
rect 92774 7686 92780 7886
rect 92734 6884 92780 7686
rect 92734 6592 92740 6884
rect 92774 6592 92780 6884
rect 92734 5790 92780 6592
rect 92734 5498 92740 5790
rect 92774 5498 92780 5790
rect 92734 4696 92780 5498
rect 92734 4404 92740 4696
rect 92774 4404 92780 4696
rect 92734 3602 92780 4404
rect 92734 3572 92740 3602
rect 91716 3310 91754 3382
rect 91672 3200 91754 3310
rect 92774 3572 92780 3602
rect 93790 7686 93798 7906
rect 94966 7976 95034 8154
rect 93832 7686 93836 7906
rect 93790 6884 93836 7686
rect 93790 6592 93798 6884
rect 93832 6592 93836 6884
rect 93790 5790 93836 6592
rect 94966 7684 94980 7976
rect 95014 7874 95034 7976
rect 96038 7976 96072 7992
rect 94966 7668 95014 7684
rect 96034 7684 96038 7882
rect 97070 7976 97138 8154
rect 97070 7888 97096 7976
rect 96072 7684 96080 7882
rect 94966 6898 95012 7668
rect 94966 6882 95014 6898
rect 94966 6590 94980 6882
rect 94966 6574 95014 6590
rect 96034 6882 96080 7684
rect 96034 6590 96038 6882
rect 96072 6590 96080 6882
rect 93790 5498 93798 5790
rect 93832 5498 93836 5790
rect 93790 4696 93836 5498
rect 94326 6442 94476 6568
rect 94326 5246 94348 6442
rect 94442 5246 94476 6442
rect 94326 4922 94476 5246
rect 94966 5804 95012 6574
rect 94966 5788 95014 5804
rect 94966 5496 94980 5788
rect 94966 5480 95014 5496
rect 96034 5788 96080 6590
rect 96034 5496 96038 5788
rect 96072 5496 96080 5788
rect 93790 4404 93798 4696
rect 93832 4404 93836 4696
rect 93790 3602 93836 4404
rect 93790 3544 93798 3602
rect 92740 3294 92774 3310
rect 93774 3310 93798 3404
rect 93832 3544 93836 3602
rect 94966 4710 95012 5480
rect 94966 4694 95014 4710
rect 94966 4402 94980 4694
rect 94966 4386 95014 4402
rect 96034 4694 96080 5496
rect 96034 4402 96038 4694
rect 96072 4402 96080 4694
rect 94966 3616 95012 4386
rect 94966 3600 95014 3616
rect 94966 3542 94980 3600
rect 93832 3310 93856 3404
rect 93774 3206 93856 3310
rect 96034 3600 96080 4402
rect 96034 3520 96038 3600
rect 94980 3292 95014 3308
rect 96018 3308 96038 3408
rect 96072 3520 96080 3600
rect 97086 7684 97096 7888
rect 97130 7940 97138 7976
rect 98154 7976 98188 7992
rect 97130 7888 97144 7940
rect 97130 7684 97132 7888
rect 97086 6882 97132 7684
rect 97086 6590 97096 6882
rect 97130 6590 97132 6882
rect 97086 5788 97132 6590
rect 97086 5496 97096 5788
rect 97130 5496 97132 5788
rect 97086 4694 97132 5496
rect 97086 4402 97096 4694
rect 97130 4402 97132 4694
rect 97086 3600 97132 4402
rect 97086 3542 97096 3600
rect 96072 3308 96100 3408
rect 96018 3206 96100 3308
rect 97130 3542 97132 3600
rect 99186 7976 99270 8164
rect 98188 7684 98200 7888
rect 99186 7884 99212 7976
rect 98154 6882 98200 7684
rect 98188 6590 98200 6882
rect 98154 5788 98200 6590
rect 98188 5496 98200 5788
rect 98154 4694 98200 5496
rect 98188 4402 98200 4694
rect 98154 3600 98200 4402
rect 97096 3292 97130 3308
rect 98144 3308 98154 3380
rect 98188 3526 98200 3600
rect 99206 7684 99212 7884
rect 99246 7884 99270 7976
rect 100270 7976 100304 7992
rect 99246 7684 99252 7884
rect 99206 6882 99252 7684
rect 99206 6590 99212 6882
rect 99246 6590 99252 6882
rect 99206 5788 99252 6590
rect 99206 5496 99212 5788
rect 99246 5496 99252 5788
rect 99206 4694 99252 5496
rect 99206 4402 99212 4694
rect 99246 4402 99252 4694
rect 99206 3600 99252 4402
rect 99206 3570 99212 3600
rect 98188 3308 98226 3380
rect 93774 3200 96130 3206
rect 89546 3198 96130 3200
rect 98144 3198 98226 3308
rect 99246 3570 99252 3600
rect 100262 7684 100270 7904
rect 100304 7684 100308 7904
rect 100262 6882 100308 7684
rect 100262 6590 100270 6882
rect 100304 6590 100308 6882
rect 100262 5788 100308 6590
rect 100262 5496 100270 5788
rect 100304 5496 100308 5788
rect 100262 4694 100308 5496
rect 100262 4402 100270 4694
rect 100304 4402 100308 4694
rect 100262 3600 100308 4402
rect 100262 3542 100270 3600
rect 99212 3292 99246 3308
rect 100246 3308 100270 3402
rect 100304 3542 100308 3600
rect 100608 7468 101298 7712
rect 100304 3308 100328 3402
rect 100246 3198 100328 3308
rect 100608 3350 100786 7468
rect 101166 3350 101298 7468
rect 89546 3110 100468 3198
rect 100608 3172 101298 3350
rect 80574 3104 82896 3110
rect 84910 3088 84992 3110
rect 89558 3104 100468 3110
rect 91672 3082 91754 3104
rect 93808 3102 100468 3104
rect 93808 3096 96130 3102
rect 98144 3080 98226 3102
<< viali >>
rect 72632 74380 72838 74482
rect 80464 74422 80754 74572
rect 71338 73868 71372 74040
rect 43052 73478 45226 73680
rect 47060 73476 49234 73678
rect 51072 73476 53246 73678
rect 55082 73476 57256 73678
rect 71996 73868 72030 74040
rect 72654 73868 72688 74040
rect 73312 73868 73346 74040
rect 73970 73868 74004 74040
rect 75202 73848 75236 74020
rect 75860 73848 75894 74020
rect 76518 73848 76552 74020
rect 77176 73848 77210 74020
rect 77834 73848 77868 74020
rect 79052 73862 79086 74034
rect 79710 73862 79744 74034
rect 80368 73862 80402 74034
rect 81026 73862 81060 74034
rect 81684 73862 81718 74034
rect 42410 73194 42582 73228
rect 43104 73194 43276 73228
rect 43798 73194 43970 73228
rect 44492 73194 44664 73228
rect 45186 73194 45358 73228
rect 46418 73192 46590 73226
rect 47112 73192 47284 73226
rect 47806 73192 47978 73226
rect 48500 73192 48672 73226
rect 49194 73192 49366 73226
rect 50430 73192 50602 73226
rect 51124 73192 51296 73226
rect 51818 73192 51990 73226
rect 52512 73192 52684 73226
rect 53206 73192 53378 73226
rect 54440 73192 54612 73226
rect 55134 73192 55306 73226
rect 55828 73192 56000 73226
rect 56522 73192 56694 73226
rect 57216 73192 57388 73226
rect 42410 72536 42582 72570
rect 43104 72536 43276 72570
rect 43798 72536 43970 72570
rect 44492 72536 44664 72570
rect 45186 72536 45358 72570
rect 46418 72534 46590 72568
rect 47112 72534 47284 72568
rect 47806 72534 47978 72568
rect 48500 72534 48672 72568
rect 49194 72534 49366 72568
rect 42410 71878 42582 71912
rect 43104 71878 43276 71912
rect 43798 71878 43970 71912
rect 44492 71878 44664 71912
rect 45186 71878 45358 71912
rect 42410 71220 42582 71254
rect 43104 71220 43276 71254
rect 43798 71220 43970 71254
rect 44492 71220 44664 71254
rect 45186 71220 45358 71254
rect 50430 72534 50602 72568
rect 51124 72534 51296 72568
rect 51818 72534 51990 72568
rect 52512 72534 52684 72568
rect 53206 72534 53378 72568
rect 46418 71876 46590 71910
rect 47112 71876 47284 71910
rect 47806 71876 47978 71910
rect 48500 71876 48672 71910
rect 49194 71876 49366 71910
rect 46418 71218 46590 71252
rect 47112 71218 47284 71252
rect 47806 71218 47978 71252
rect 48500 71218 48672 71252
rect 49194 71218 49366 71252
rect 42410 70562 42582 70596
rect 43104 70562 43276 70596
rect 43798 70562 43970 70596
rect 44492 70562 44664 70596
rect 45186 70562 45358 70596
rect 54440 72534 54612 72568
rect 55134 72534 55306 72568
rect 55828 72534 56000 72568
rect 56522 72534 56694 72568
rect 57216 72534 57388 72568
rect 50430 71876 50602 71910
rect 51124 71876 51296 71910
rect 51818 71876 51990 71910
rect 52512 71876 52684 71910
rect 53206 71876 53378 71910
rect 50430 71218 50602 71252
rect 51124 71218 51296 71252
rect 51818 71218 51990 71252
rect 52512 71218 52684 71252
rect 53206 71218 53378 71252
rect 46418 70560 46590 70594
rect 47112 70560 47284 70594
rect 47806 70560 47978 70594
rect 48500 70560 48672 70594
rect 49194 70560 49366 70594
rect 54440 71876 54612 71910
rect 55134 71876 55306 71910
rect 55828 71876 56000 71910
rect 56522 71876 56694 71910
rect 57216 71876 57388 71910
rect 54440 71218 54612 71252
rect 55134 71218 55306 71252
rect 55828 71218 56000 71252
rect 56522 71218 56694 71252
rect 57216 71218 57388 71252
rect 50430 70560 50602 70594
rect 51124 70560 51296 70594
rect 51818 70560 51990 70594
rect 52512 70560 52684 70594
rect 53206 70560 53378 70594
rect 54440 70560 54612 70594
rect 55134 70560 55306 70594
rect 55828 70560 56000 70594
rect 56522 70560 56694 70594
rect 57216 70560 57388 70594
rect 42410 69904 42582 69938
rect 43104 69904 43276 69938
rect 43798 69904 43970 69938
rect 44492 69904 44664 69938
rect 45186 69904 45358 69938
rect 46418 69902 46590 69936
rect 47112 69902 47284 69936
rect 47806 69902 47978 69936
rect 48500 69902 48672 69936
rect 49194 69902 49366 69936
rect 50430 69902 50602 69936
rect 51124 69902 51296 69936
rect 51818 69902 51990 69936
rect 52512 69902 52684 69936
rect 53206 69902 53378 69936
rect 54440 69902 54612 69936
rect 55134 69902 55306 69936
rect 55828 69902 56000 69936
rect 56522 69902 56694 69936
rect 57216 69902 57388 69936
rect 71066 70412 71150 72980
rect 71310 72954 71344 73126
rect 71310 72260 71344 72432
rect 71310 71566 71344 71738
rect 71310 70872 71344 71044
rect 71310 70178 71344 70350
rect 71968 72954 72002 73126
rect 71968 72260 72002 72432
rect 71968 71566 72002 71738
rect 71968 70872 72002 71044
rect 43044 69280 45218 69482
rect 47038 69280 49212 69482
rect 51060 69280 53234 69482
rect 55082 69280 57256 69482
rect 57740 69482 57844 69662
rect 71968 70178 72002 70350
rect 72626 72954 72660 73126
rect 72626 72260 72660 72432
rect 72626 71566 72660 71738
rect 72626 70872 72660 71044
rect 72626 70178 72660 70350
rect 73284 72954 73318 73126
rect 73284 72260 73318 72432
rect 73284 71566 73318 71738
rect 73284 70872 73318 71044
rect 73284 70178 73318 70350
rect 73942 72954 73976 73126
rect 73942 72260 73976 72432
rect 73942 71566 73976 71738
rect 73942 70872 73976 71044
rect 73942 70178 73976 70350
rect 74930 70392 75014 72960
rect 75174 72934 75208 73106
rect 75174 72240 75208 72412
rect 75174 71546 75208 71718
rect 75174 70852 75208 71024
rect 75174 70158 75208 70330
rect 75832 72934 75866 73106
rect 75832 72240 75866 72412
rect 75832 71546 75866 71718
rect 75832 70852 75866 71024
rect 42402 68996 42574 69030
rect 43096 68996 43268 69030
rect 43790 68996 43962 69030
rect 44484 68996 44656 69030
rect 45178 68996 45350 69030
rect 46396 68996 46568 69030
rect 47090 68996 47262 69030
rect 47784 68996 47956 69030
rect 48478 68996 48650 69030
rect 49172 68996 49344 69030
rect 50418 68996 50590 69030
rect 51112 68996 51284 69030
rect 51806 68996 51978 69030
rect 52500 68996 52672 69030
rect 53194 68996 53366 69030
rect 54440 68996 54612 69030
rect 55134 68996 55306 69030
rect 55828 68996 56000 69030
rect 56522 68996 56694 69030
rect 57216 68996 57388 69030
rect 42402 68338 42574 68372
rect 43096 68338 43268 68372
rect 43790 68338 43962 68372
rect 44484 68338 44656 68372
rect 45178 68338 45350 68372
rect 46396 68338 46568 68372
rect 47090 68338 47262 68372
rect 47784 68338 47956 68372
rect 48478 68338 48650 68372
rect 49172 68338 49344 68372
rect 42402 67680 42574 67714
rect 43096 67680 43268 67714
rect 43790 67680 43962 67714
rect 44484 67680 44656 67714
rect 45178 67680 45350 67714
rect 42402 67022 42574 67056
rect 43096 67022 43268 67056
rect 43790 67022 43962 67056
rect 44484 67022 44656 67056
rect 45178 67022 45350 67056
rect 1086 65834 2490 65904
rect 3754 65830 5158 65900
rect 6428 65836 7832 65906
rect 9074 65836 10478 65906
rect 11728 65830 13132 65900
rect 14382 65836 15786 65906
rect 17008 65840 18412 65910
rect 19562 65816 20520 65924
rect 50418 68338 50590 68372
rect 51112 68338 51284 68372
rect 51806 68338 51978 68372
rect 52500 68338 52672 68372
rect 53194 68338 53366 68372
rect 46396 67680 46568 67714
rect 47090 67680 47262 67714
rect 47784 67680 47956 67714
rect 48478 67680 48650 67714
rect 49172 67680 49344 67714
rect 46396 67022 46568 67056
rect 47090 67022 47262 67056
rect 47784 67022 47956 67056
rect 48478 67022 48650 67056
rect 49172 67022 49344 67056
rect 42402 66364 42574 66398
rect 43096 66364 43268 66398
rect 43790 66364 43962 66398
rect 44484 66364 44656 66398
rect 45178 66364 45350 66398
rect 54440 68338 54612 68372
rect 55134 68338 55306 68372
rect 55828 68338 56000 68372
rect 56522 68338 56694 68372
rect 57216 68338 57388 68372
rect 50418 67680 50590 67714
rect 51112 67680 51284 67714
rect 51806 67680 51978 67714
rect 52500 67680 52672 67714
rect 53194 67680 53366 67714
rect 50418 67022 50590 67056
rect 51112 67022 51284 67056
rect 51806 67022 51978 67056
rect 52500 67022 52672 67056
rect 53194 67022 53366 67056
rect 46396 66364 46568 66398
rect 47090 66364 47262 66398
rect 47784 66364 47956 66398
rect 48478 66364 48650 66398
rect 49172 66364 49344 66398
rect 54440 67680 54612 67714
rect 55134 67680 55306 67714
rect 55828 67680 56000 67714
rect 56522 67680 56694 67714
rect 57216 67680 57388 67714
rect 54440 67022 54612 67056
rect 55134 67022 55306 67056
rect 55828 67022 56000 67056
rect 56522 67022 56694 67056
rect 57216 67022 57388 67056
rect 50418 66364 50590 66398
rect 51112 66364 51284 66398
rect 51806 66364 51978 66398
rect 52500 66364 52672 66398
rect 53194 66364 53366 66398
rect 71062 66636 71146 69204
rect 71306 69178 71340 69350
rect 71306 68484 71340 68656
rect 71306 67790 71340 67962
rect 71306 67096 71340 67268
rect 54440 66364 54612 66398
rect 55134 66364 55306 66398
rect 55828 66364 56000 66398
rect 56522 66364 56694 66398
rect 57216 66364 57388 66398
rect 71306 66402 71340 66574
rect 71964 69178 71998 69350
rect 75832 70158 75866 70330
rect 76490 72934 76524 73106
rect 76490 72240 76524 72412
rect 76490 71546 76524 71718
rect 76490 70852 76524 71024
rect 76490 70158 76524 70330
rect 77148 72934 77182 73106
rect 77148 72240 77182 72412
rect 77148 71546 77182 71718
rect 77148 70852 77182 71024
rect 77148 70158 77182 70330
rect 77806 72934 77840 73106
rect 77806 72240 77840 72412
rect 77806 71546 77840 71718
rect 77806 70852 77840 71024
rect 77806 70158 77840 70330
rect 78780 70406 78864 72974
rect 79024 72948 79058 73120
rect 79024 72254 79058 72426
rect 79024 71560 79058 71732
rect 79024 70866 79058 71038
rect 79024 70172 79058 70344
rect 79682 72948 79716 73120
rect 79682 72254 79716 72426
rect 79682 71560 79716 71732
rect 79682 70866 79716 71038
rect 71964 68484 71998 68656
rect 71964 67790 71998 67962
rect 71964 67096 71998 67268
rect 42402 65706 42574 65740
rect 43096 65706 43268 65740
rect 43790 65706 43962 65740
rect 44484 65706 44656 65740
rect 45178 65706 45350 65740
rect 46396 65706 46568 65740
rect 47090 65706 47262 65740
rect 47784 65706 47956 65740
rect 48478 65706 48650 65740
rect 49172 65706 49344 65740
rect 50418 65706 50590 65740
rect 51112 65706 51284 65740
rect 51806 65706 51978 65740
rect 52500 65706 52672 65740
rect 53194 65706 53366 65740
rect 54440 65706 54612 65740
rect 55134 65706 55306 65740
rect 55828 65706 56000 65740
rect 56522 65706 56694 65740
rect 57216 65706 57388 65740
rect 71964 66402 71998 66574
rect 72622 69178 72656 69350
rect 72622 68484 72656 68656
rect 72622 67790 72656 67962
rect 72622 67096 72656 67268
rect 72622 66402 72656 66574
rect 73280 69178 73314 69350
rect 73280 68484 73314 68656
rect 73280 67790 73314 67962
rect 73280 67096 73314 67268
rect 73280 66402 73314 66574
rect 73938 69178 73972 69350
rect 73938 68484 73972 68656
rect 73938 67790 73972 67962
rect 73938 67096 73972 67268
rect 73938 66402 73972 66574
rect 74926 66616 75010 69184
rect 75170 69158 75204 69330
rect 75170 68464 75204 68636
rect 75170 67770 75204 67942
rect 75170 67076 75204 67248
rect 75170 66382 75204 66554
rect 75828 69158 75862 69330
rect 79682 70172 79716 70344
rect 80340 72948 80374 73120
rect 80340 72254 80374 72426
rect 80340 71560 80374 71732
rect 80340 70866 80374 71038
rect 80340 70172 80374 70344
rect 80998 72948 81032 73120
rect 80998 72254 81032 72426
rect 80998 71560 81032 71732
rect 80998 70866 81032 71038
rect 80998 70172 81032 70344
rect 81656 72948 81690 73120
rect 81656 72254 81690 72426
rect 81656 71560 81690 71732
rect 81656 70866 81690 71038
rect 81656 70172 81690 70344
rect 75828 68464 75862 68636
rect 75828 67770 75862 67942
rect 75828 67076 75862 67248
rect 19572 65586 19744 65620
rect 20266 65586 20438 65620
rect 966 65536 1138 65570
rect 1660 65536 1832 65570
rect 2354 65536 2526 65570
rect 3634 65532 3806 65566
rect 4328 65532 4500 65566
rect 5022 65532 5194 65566
rect 6308 65538 6480 65572
rect 7002 65538 7174 65572
rect 7696 65538 7868 65572
rect 8954 65538 9126 65572
rect 9648 65538 9820 65572
rect 10342 65538 10514 65572
rect 11608 65532 11780 65566
rect 12302 65532 12474 65566
rect 12996 65532 13168 65566
rect 14262 65538 14434 65572
rect 14956 65538 15128 65572
rect 15650 65538 15822 65572
rect 16888 65542 17060 65576
rect 17582 65542 17754 65576
rect 18276 65542 18448 65576
rect 966 64878 1138 64912
rect 1660 64878 1832 64912
rect 2354 64878 2526 64912
rect 966 64220 1138 64254
rect 1660 64220 1832 64254
rect 2354 64220 2526 64254
rect 966 63562 1138 63596
rect 1660 63562 1832 63596
rect 2354 63562 2526 63596
rect 966 62904 1138 62938
rect 1660 62904 1832 62938
rect 2354 62904 2526 62938
rect 966 62246 1138 62280
rect 1660 62246 1832 62280
rect 2354 62246 2526 62280
rect 3634 64874 3806 64908
rect 4328 64874 4500 64908
rect 5022 64874 5194 64908
rect 3634 64216 3806 64250
rect 4328 64216 4500 64250
rect 5022 64216 5194 64250
rect 3634 63558 3806 63592
rect 4328 63558 4500 63592
rect 5022 63558 5194 63592
rect 3634 62900 3806 62934
rect 4328 62900 4500 62934
rect 5022 62900 5194 62934
rect 3634 62242 3806 62276
rect 4328 62242 4500 62276
rect 5022 62242 5194 62276
rect 966 61588 1138 61622
rect 1660 61588 1832 61622
rect 2354 61588 2526 61622
rect 966 60930 1138 60964
rect 1660 60930 1832 60964
rect 2354 60930 2526 60964
rect 3086 60716 3304 61070
rect 6308 64880 6480 64914
rect 7002 64880 7174 64914
rect 7696 64880 7868 64914
rect 6308 64222 6480 64256
rect 7002 64222 7174 64256
rect 7696 64222 7868 64256
rect 6308 63564 6480 63598
rect 7002 63564 7174 63598
rect 7696 63564 7868 63598
rect 6308 62906 6480 62940
rect 7002 62906 7174 62940
rect 7696 62906 7868 62940
rect 6308 62248 6480 62282
rect 7002 62248 7174 62282
rect 7696 62248 7868 62282
rect 3634 61584 3806 61618
rect 4328 61584 4500 61618
rect 5022 61584 5194 61618
rect 3634 60926 3806 60960
rect 4328 60926 4500 60960
rect 5022 60926 5194 60960
rect 5720 60742 5956 61104
rect 8954 64880 9126 64914
rect 9648 64880 9820 64914
rect 10342 64880 10514 64914
rect 8954 64222 9126 64256
rect 9648 64222 9820 64256
rect 10342 64222 10514 64256
rect 8954 63564 9126 63598
rect 9648 63564 9820 63598
rect 10342 63564 10514 63598
rect 8954 62906 9126 62940
rect 9648 62906 9820 62940
rect 10342 62906 10514 62940
rect 8954 62248 9126 62282
rect 9648 62248 9820 62282
rect 10342 62248 10514 62282
rect 6308 61590 6480 61624
rect 7002 61590 7174 61624
rect 7696 61590 7868 61624
rect 6308 60932 6480 60966
rect 7002 60932 7174 60966
rect 7696 60932 7868 60966
rect 8380 60692 8582 61180
rect 11608 64874 11780 64908
rect 12302 64874 12474 64908
rect 12996 64874 13168 64908
rect 11608 64216 11780 64250
rect 12302 64216 12474 64250
rect 12996 64216 13168 64250
rect 11608 63558 11780 63592
rect 12302 63558 12474 63592
rect 12996 63558 13168 63592
rect 11608 62900 11780 62934
rect 12302 62900 12474 62934
rect 12996 62900 13168 62934
rect 11608 62242 11780 62276
rect 12302 62242 12474 62276
rect 12996 62242 13168 62276
rect 8954 61590 9126 61624
rect 9648 61590 9820 61624
rect 10342 61590 10514 61624
rect 8954 60932 9126 60966
rect 9648 60932 9820 60966
rect 10342 60932 10514 60966
rect 11056 60658 11274 61096
rect 14262 64880 14434 64914
rect 14956 64880 15128 64914
rect 15650 64880 15822 64914
rect 14262 64222 14434 64256
rect 14956 64222 15128 64256
rect 15650 64222 15822 64256
rect 14262 63564 14434 63598
rect 14956 63564 15128 63598
rect 15650 63564 15822 63598
rect 14262 62906 14434 62940
rect 14956 62906 15128 62940
rect 15650 62906 15822 62940
rect 14262 62248 14434 62282
rect 14956 62248 15128 62282
rect 15650 62248 15822 62282
rect 11608 61584 11780 61618
rect 12302 61584 12474 61618
rect 12996 61584 13168 61618
rect 11608 60926 11780 60960
rect 12302 60926 12474 60960
rect 12996 60926 13168 60960
rect 13706 60700 13874 61128
rect 16888 64884 17060 64918
rect 17582 64884 17754 64918
rect 18276 64884 18448 64918
rect 19572 64928 19744 64962
rect 20266 64928 20438 64962
rect 16888 64226 17060 64260
rect 17582 64226 17754 64260
rect 18276 64226 18448 64260
rect 16888 63568 17060 63602
rect 17582 63568 17754 63602
rect 18276 63568 18448 63602
rect 16888 62910 17060 62944
rect 17582 62910 17754 62944
rect 18276 62910 18448 62944
rect 16888 62252 17060 62286
rect 17582 62252 17754 62286
rect 18276 62252 18448 62286
rect 14262 61590 14434 61624
rect 14956 61590 15128 61624
rect 15650 61590 15822 61624
rect 14262 60932 14434 60966
rect 14956 60932 15128 60966
rect 15650 60932 15822 60966
rect 16322 60800 16576 61070
rect 43032 64806 45206 65008
rect 47040 64804 49214 65006
rect 51052 64804 53226 65006
rect 55062 64804 57236 65006
rect 42390 64522 42562 64556
rect 43084 64522 43256 64556
rect 43778 64522 43950 64556
rect 44472 64522 44644 64556
rect 45166 64522 45338 64556
rect 46398 64520 46570 64554
rect 47092 64520 47264 64554
rect 47786 64520 47958 64554
rect 48480 64520 48652 64554
rect 49174 64520 49346 64554
rect 50410 64520 50582 64554
rect 51104 64520 51276 64554
rect 51798 64520 51970 64554
rect 52492 64520 52664 64554
rect 53186 64520 53358 64554
rect 54420 64520 54592 64554
rect 55114 64520 55286 64554
rect 55808 64520 55980 64554
rect 56502 64520 56674 64554
rect 57196 64520 57368 64554
rect 19572 64270 19744 64304
rect 20266 64270 20438 64304
rect 20732 64074 20782 64112
rect 19572 63612 19744 63646
rect 20266 63612 20438 63646
rect 41840 64136 42022 64304
rect 42390 63864 42562 63898
rect 43084 63864 43256 63898
rect 43778 63864 43950 63898
rect 44472 63864 44644 63898
rect 45166 63864 45338 63898
rect 19572 62954 19744 62988
rect 20266 62954 20438 62988
rect 19572 62296 19744 62330
rect 20266 62296 20438 62330
rect 16888 61594 17060 61628
rect 17582 61594 17754 61628
rect 18276 61594 18448 61628
rect 16888 60936 17060 60970
rect 17582 60936 17754 60970
rect 18276 60936 18448 60970
rect 18872 60816 19082 61162
rect 46398 63862 46570 63896
rect 47092 63862 47264 63896
rect 47786 63862 47958 63896
rect 48480 63862 48652 63896
rect 49174 63862 49346 63896
rect 42390 63206 42562 63240
rect 43084 63206 43256 63240
rect 43778 63206 43950 63240
rect 44472 63206 44644 63240
rect 45166 63206 45338 63240
rect 42390 62548 42562 62582
rect 43084 62548 43256 62582
rect 43778 62548 43950 62582
rect 44472 62548 44644 62582
rect 45166 62548 45338 62582
rect 19572 61638 19744 61672
rect 20266 61638 20438 61672
rect 19572 60980 19744 61014
rect 20266 60980 20438 61014
rect 50410 63862 50582 63896
rect 51104 63862 51276 63896
rect 51798 63862 51970 63896
rect 52492 63862 52664 63896
rect 53186 63862 53358 63896
rect 46398 63204 46570 63238
rect 47092 63204 47264 63238
rect 47786 63204 47958 63238
rect 48480 63204 48652 63238
rect 49174 63204 49346 63238
rect 46398 62546 46570 62580
rect 47092 62546 47264 62580
rect 47786 62546 47958 62580
rect 48480 62546 48652 62580
rect 49174 62546 49346 62580
rect 42390 61890 42562 61924
rect 43084 61890 43256 61924
rect 43778 61890 43950 61924
rect 44472 61890 44644 61924
rect 45166 61890 45338 61924
rect 19572 60322 19744 60356
rect 20266 60322 20438 60356
rect 966 60272 1138 60306
rect 1660 60272 1832 60306
rect 2354 60272 2526 60306
rect 3634 60268 3806 60302
rect 4328 60268 4500 60302
rect 5022 60268 5194 60302
rect 6308 60274 6480 60308
rect 7002 60274 7174 60308
rect 7696 60274 7868 60308
rect 8954 60274 9126 60308
rect 9648 60274 9820 60308
rect 10342 60274 10514 60308
rect 11608 60268 11780 60302
rect 12302 60268 12474 60302
rect 12996 60268 13168 60302
rect 14262 60274 14434 60308
rect 14956 60274 15128 60308
rect 15650 60274 15822 60308
rect 16888 60278 17060 60312
rect 17582 60278 17754 60312
rect 18276 60278 18448 60312
rect 54420 63862 54592 63896
rect 55114 63862 55286 63896
rect 55808 63862 55980 63896
rect 56502 63862 56674 63896
rect 57196 63862 57368 63896
rect 50410 63204 50582 63238
rect 51104 63204 51276 63238
rect 51798 63204 51970 63238
rect 52492 63204 52664 63238
rect 53186 63204 53358 63238
rect 50410 62546 50582 62580
rect 51104 62546 51276 62580
rect 51798 62546 51970 62580
rect 52492 62546 52664 62580
rect 53186 62546 53358 62580
rect 46398 61888 46570 61922
rect 47092 61888 47264 61922
rect 47786 61888 47958 61922
rect 48480 61888 48652 61922
rect 49174 61888 49346 61922
rect 54420 63204 54592 63238
rect 55114 63204 55286 63238
rect 55808 63204 55980 63238
rect 56502 63204 56674 63238
rect 57196 63204 57368 63238
rect 54420 62546 54592 62580
rect 55114 62546 55286 62580
rect 55808 62546 55980 62580
rect 56502 62546 56674 62580
rect 57196 62546 57368 62580
rect 50410 61888 50582 61922
rect 51104 61888 51276 61922
rect 51798 61888 51970 61922
rect 52492 61888 52664 61922
rect 53186 61888 53358 61922
rect 71062 62866 71146 65434
rect 71306 65408 71340 65580
rect 71306 64714 71340 64886
rect 71306 64020 71340 64192
rect 71306 63326 71340 63498
rect 71306 62632 71340 62804
rect 71964 65408 71998 65580
rect 75828 66382 75862 66554
rect 76486 69158 76520 69330
rect 76486 68464 76520 68636
rect 76486 67770 76520 67942
rect 76486 67076 76520 67248
rect 76486 66382 76520 66554
rect 77144 69158 77178 69330
rect 77144 68464 77178 68636
rect 77144 67770 77178 67942
rect 77144 67076 77178 67248
rect 77144 66382 77178 66554
rect 77802 69158 77836 69330
rect 77802 68464 77836 68636
rect 77802 67770 77836 67942
rect 77802 67076 77836 67248
rect 77802 66382 77836 66554
rect 78776 66630 78860 69198
rect 79020 69172 79054 69344
rect 79020 68478 79054 68650
rect 79020 67784 79054 67956
rect 79020 67090 79054 67262
rect 79020 66396 79054 66568
rect 79678 69172 79712 69344
rect 79678 68478 79712 68650
rect 79678 67784 79712 67956
rect 79678 67090 79712 67262
rect 79678 66396 79712 66568
rect 80336 69172 80370 69344
rect 80336 68478 80370 68650
rect 80336 67784 80370 67956
rect 80336 67090 80370 67262
rect 80336 66396 80370 66568
rect 80994 69172 81028 69344
rect 80994 68478 81028 68650
rect 80994 67784 81028 67956
rect 80994 67090 81028 67262
rect 80994 66396 81028 66568
rect 81652 69172 81686 69344
rect 81652 68478 81686 68650
rect 81652 67784 81686 67956
rect 81652 67090 81686 67262
rect 81652 66396 81686 66568
rect 71964 64714 71998 64886
rect 71964 64020 71998 64192
rect 71964 63326 71998 63498
rect 71964 62632 71998 62804
rect 72622 65408 72656 65580
rect 72622 64714 72656 64886
rect 72622 64020 72656 64192
rect 72622 63326 72656 63498
rect 72622 62632 72656 62804
rect 73280 65408 73314 65580
rect 73280 64714 73314 64886
rect 73280 64020 73314 64192
rect 73280 63326 73314 63498
rect 73280 62632 73314 62804
rect 73938 65408 73972 65580
rect 73938 64714 73972 64886
rect 73938 64020 73972 64192
rect 73938 63326 73972 63498
rect 73938 62632 73972 62804
rect 74926 62846 75010 65414
rect 75170 65388 75204 65560
rect 75170 64694 75204 64866
rect 75170 64000 75204 64172
rect 75170 63306 75204 63478
rect 75170 62612 75204 62784
rect 75828 65388 75862 65560
rect 75828 64694 75862 64866
rect 75828 64000 75862 64172
rect 75828 63306 75862 63478
rect 54420 61888 54592 61922
rect 55114 61888 55286 61922
rect 55808 61888 55980 61922
rect 56502 61888 56674 61922
rect 57196 61888 57368 61922
rect 42390 61232 42562 61266
rect 43084 61232 43256 61266
rect 43778 61232 43950 61266
rect 44472 61232 44644 61266
rect 45166 61232 45338 61266
rect 46398 61230 46570 61264
rect 47092 61230 47264 61264
rect 47786 61230 47958 61264
rect 48480 61230 48652 61264
rect 49174 61230 49346 61264
rect 50410 61230 50582 61264
rect 51104 61230 51276 61264
rect 51798 61230 51970 61264
rect 52492 61230 52664 61264
rect 53186 61230 53358 61264
rect 54420 61230 54592 61264
rect 55114 61230 55286 61264
rect 55808 61230 55980 61264
rect 56502 61230 56674 61264
rect 57196 61230 57368 61264
rect 43024 60608 45198 60810
rect 47018 60608 49192 60810
rect 51040 60608 53214 60810
rect 55062 60608 57236 60810
rect 57798 60588 57940 61090
rect 42382 60324 42554 60358
rect 43076 60324 43248 60358
rect 43770 60324 43942 60358
rect 44464 60324 44636 60358
rect 45158 60324 45330 60358
rect 46376 60324 46548 60358
rect 47070 60324 47242 60358
rect 47764 60324 47936 60358
rect 48458 60324 48630 60358
rect 49152 60324 49324 60358
rect 50398 60324 50570 60358
rect 51092 60324 51264 60358
rect 51786 60324 51958 60358
rect 52480 60324 52652 60358
rect 53174 60324 53346 60358
rect 54420 60324 54592 60358
rect 55114 60324 55286 60358
rect 55808 60324 55980 60358
rect 56502 60324 56674 60358
rect 57196 60324 57368 60358
rect 1058 59566 2462 59636
rect 3726 59562 5130 59632
rect 6400 59568 7804 59638
rect 9046 59568 10450 59638
rect 11700 59562 13104 59632
rect 14354 59568 15758 59638
rect 16980 59572 18384 59642
rect 19534 59548 20492 59656
rect 42382 59666 42554 59700
rect 43076 59666 43248 59700
rect 43770 59666 43942 59700
rect 44464 59666 44636 59700
rect 45158 59666 45330 59700
rect 19544 59318 19716 59352
rect 20238 59318 20410 59352
rect 938 59268 1110 59302
rect 1632 59268 1804 59302
rect 2326 59268 2498 59302
rect 3606 59264 3778 59298
rect 4300 59264 4472 59298
rect 4994 59264 5166 59298
rect 6280 59270 6452 59304
rect 6974 59270 7146 59304
rect 7668 59270 7840 59304
rect 8926 59270 9098 59304
rect 9620 59270 9792 59304
rect 10314 59270 10486 59304
rect 11580 59264 11752 59298
rect 12274 59264 12446 59298
rect 12968 59264 13140 59298
rect 14234 59270 14406 59304
rect 14928 59270 15100 59304
rect 15622 59270 15794 59304
rect 16860 59274 17032 59308
rect 17554 59274 17726 59308
rect 18248 59274 18420 59308
rect 938 58610 1110 58644
rect 1632 58610 1804 58644
rect 2326 58610 2498 58644
rect 338 56766 438 57716
rect 938 57952 1110 57986
rect 1632 57952 1804 57986
rect 2326 57952 2498 57986
rect 938 57294 1110 57328
rect 1632 57294 1804 57328
rect 2326 57294 2498 57328
rect 938 56636 1110 56670
rect 1632 56636 1804 56670
rect 2326 56636 2498 56670
rect 938 55978 1110 56012
rect 1632 55978 1804 56012
rect 2326 55978 2498 56012
rect 3606 58606 3778 58640
rect 4300 58606 4472 58640
rect 4994 58606 5166 58640
rect 3606 57948 3778 57982
rect 4300 57948 4472 57982
rect 4994 57948 5166 57982
rect 3606 57290 3778 57324
rect 4300 57290 4472 57324
rect 4994 57290 5166 57324
rect 3606 56632 3778 56666
rect 4300 56632 4472 56666
rect 4994 56632 5166 56666
rect 3606 55974 3778 56008
rect 4300 55974 4472 56008
rect 4994 55974 5166 56008
rect 938 55320 1110 55354
rect 1632 55320 1804 55354
rect 2326 55320 2498 55354
rect 938 54662 1110 54696
rect 1632 54662 1804 54696
rect 2326 54662 2498 54696
rect 3058 54448 3276 54802
rect 6280 58612 6452 58646
rect 6974 58612 7146 58646
rect 7668 58612 7840 58646
rect 6280 57954 6452 57988
rect 6974 57954 7146 57988
rect 7668 57954 7840 57988
rect 6280 57296 6452 57330
rect 6974 57296 7146 57330
rect 7668 57296 7840 57330
rect 6280 56638 6452 56672
rect 6974 56638 7146 56672
rect 7668 56638 7840 56672
rect 6280 55980 6452 56014
rect 6974 55980 7146 56014
rect 7668 55980 7840 56014
rect 3606 55316 3778 55350
rect 4300 55316 4472 55350
rect 4994 55316 5166 55350
rect 3606 54658 3778 54692
rect 4300 54658 4472 54692
rect 4994 54658 5166 54692
rect 5692 54474 5928 54836
rect 8926 58612 9098 58646
rect 9620 58612 9792 58646
rect 10314 58612 10486 58646
rect 8926 57954 9098 57988
rect 9620 57954 9792 57988
rect 10314 57954 10486 57988
rect 8926 57296 9098 57330
rect 9620 57296 9792 57330
rect 10314 57296 10486 57330
rect 8926 56638 9098 56672
rect 9620 56638 9792 56672
rect 10314 56638 10486 56672
rect 8926 55980 9098 56014
rect 9620 55980 9792 56014
rect 10314 55980 10486 56014
rect 6280 55322 6452 55356
rect 6974 55322 7146 55356
rect 7668 55322 7840 55356
rect 6280 54664 6452 54698
rect 6974 54664 7146 54698
rect 7668 54664 7840 54698
rect 8352 54424 8554 54912
rect 11580 58606 11752 58640
rect 12274 58606 12446 58640
rect 12968 58606 13140 58640
rect 11580 57948 11752 57982
rect 12274 57948 12446 57982
rect 12968 57948 13140 57982
rect 11580 57290 11752 57324
rect 12274 57290 12446 57324
rect 12968 57290 13140 57324
rect 11580 56632 11752 56666
rect 12274 56632 12446 56666
rect 12968 56632 13140 56666
rect 11580 55974 11752 56008
rect 12274 55974 12446 56008
rect 12968 55974 13140 56008
rect 8926 55322 9098 55356
rect 9620 55322 9792 55356
rect 10314 55322 10486 55356
rect 8926 54664 9098 54698
rect 9620 54664 9792 54698
rect 10314 54664 10486 54698
rect 11028 54390 11246 54828
rect 14234 58612 14406 58646
rect 14928 58612 15100 58646
rect 15622 58612 15794 58646
rect 14234 57954 14406 57988
rect 14928 57954 15100 57988
rect 15622 57954 15794 57988
rect 14234 57296 14406 57330
rect 14928 57296 15100 57330
rect 15622 57296 15794 57330
rect 14234 56638 14406 56672
rect 14928 56638 15100 56672
rect 15622 56638 15794 56672
rect 14234 55980 14406 56014
rect 14928 55980 15100 56014
rect 15622 55980 15794 56014
rect 11580 55316 11752 55350
rect 12274 55316 12446 55350
rect 12968 55316 13140 55350
rect 11580 54658 11752 54692
rect 12274 54658 12446 54692
rect 12968 54658 13140 54692
rect 13678 54432 13846 54860
rect 16860 58616 17032 58650
rect 17554 58616 17726 58650
rect 18248 58616 18420 58650
rect 19544 58660 19716 58694
rect 20238 58660 20410 58694
rect 16860 57958 17032 57992
rect 17554 57958 17726 57992
rect 18248 57958 18420 57992
rect 16860 57300 17032 57334
rect 17554 57300 17726 57334
rect 18248 57300 18420 57334
rect 16860 56642 17032 56676
rect 17554 56642 17726 56676
rect 18248 56642 18420 56676
rect 16860 55984 17032 56018
rect 17554 55984 17726 56018
rect 18248 55984 18420 56018
rect 14234 55322 14406 55356
rect 14928 55322 15100 55356
rect 15622 55322 15794 55356
rect 14234 54664 14406 54698
rect 14928 54664 15100 54698
rect 15622 54664 15794 54698
rect 16294 54532 16548 54802
rect 46376 59666 46548 59700
rect 47070 59666 47242 59700
rect 47764 59666 47936 59700
rect 48458 59666 48630 59700
rect 49152 59666 49324 59700
rect 42382 59008 42554 59042
rect 43076 59008 43248 59042
rect 43770 59008 43942 59042
rect 44464 59008 44636 59042
rect 45158 59008 45330 59042
rect 42382 58350 42554 58384
rect 43076 58350 43248 58384
rect 43770 58350 43942 58384
rect 44464 58350 44636 58384
rect 45158 58350 45330 58384
rect 19544 58002 19716 58036
rect 20238 58002 20410 58036
rect 19544 57344 19716 57378
rect 20238 57344 20410 57378
rect 23634 57446 23806 57480
rect 24328 57446 24500 57480
rect 25022 57446 25194 57480
rect 25716 57446 25888 57480
rect 26410 57446 26582 57480
rect 27104 57446 27276 57480
rect 27798 57446 27970 57480
rect 28492 57446 28664 57480
rect 29186 57446 29358 57480
rect 29880 57446 30052 57480
rect 50398 59666 50570 59700
rect 51092 59666 51264 59700
rect 51786 59666 51958 59700
rect 52480 59666 52652 59700
rect 53174 59666 53346 59700
rect 46376 59008 46548 59042
rect 47070 59008 47242 59042
rect 47764 59008 47936 59042
rect 48458 59008 48630 59042
rect 49152 59008 49324 59042
rect 46376 58350 46548 58384
rect 47070 58350 47242 58384
rect 47764 58350 47936 58384
rect 48458 58350 48630 58384
rect 49152 58350 49324 58384
rect 42382 57692 42554 57726
rect 43076 57692 43248 57726
rect 43770 57692 43942 57726
rect 44464 57692 44636 57726
rect 45158 57692 45330 57726
rect 54420 59666 54592 59700
rect 55114 59666 55286 59700
rect 55808 59666 55980 59700
rect 56502 59666 56674 59700
rect 57196 59666 57368 59700
rect 50398 59008 50570 59042
rect 51092 59008 51264 59042
rect 51786 59008 51958 59042
rect 52480 59008 52652 59042
rect 53174 59008 53346 59042
rect 50398 58350 50570 58384
rect 51092 58350 51264 58384
rect 51786 58350 51958 58384
rect 52480 58350 52652 58384
rect 53174 58350 53346 58384
rect 46376 57692 46548 57726
rect 47070 57692 47242 57726
rect 47764 57692 47936 57726
rect 48458 57692 48630 57726
rect 49152 57692 49324 57726
rect 54420 59008 54592 59042
rect 55114 59008 55286 59042
rect 55808 59008 55980 59042
rect 56502 59008 56674 59042
rect 57196 59008 57368 59042
rect 71062 59102 71146 61670
rect 71306 61644 71340 61816
rect 71306 60950 71340 61122
rect 71306 60256 71340 60428
rect 71306 59562 71340 59734
rect 71964 61644 71998 61816
rect 75828 62612 75862 62784
rect 76486 65388 76520 65560
rect 76486 64694 76520 64866
rect 76486 64000 76520 64172
rect 76486 63306 76520 63478
rect 76486 62612 76520 62784
rect 77144 65388 77178 65560
rect 77144 64694 77178 64866
rect 77144 64000 77178 64172
rect 77144 63306 77178 63478
rect 77144 62612 77178 62784
rect 77802 65388 77836 65560
rect 77802 64694 77836 64866
rect 77802 64000 77836 64172
rect 77802 63306 77836 63478
rect 77802 62612 77836 62784
rect 78776 62860 78860 65428
rect 79020 65402 79054 65574
rect 79020 64708 79054 64880
rect 79020 64014 79054 64186
rect 79020 63320 79054 63492
rect 79020 62626 79054 62798
rect 79678 65402 79712 65574
rect 79678 64708 79712 64880
rect 79678 64014 79712 64186
rect 79678 63320 79712 63492
rect 71964 60950 71998 61122
rect 71964 60256 71998 60428
rect 71964 59562 71998 59734
rect 54420 58350 54592 58384
rect 55114 58350 55286 58384
rect 55808 58350 55980 58384
rect 56502 58350 56674 58384
rect 57196 58350 57368 58384
rect 50398 57692 50570 57726
rect 51092 57692 51264 57726
rect 51786 57692 51958 57726
rect 52480 57692 52652 57726
rect 53174 57692 53346 57726
rect 71306 58868 71340 59040
rect 71964 58868 71998 59040
rect 72622 61644 72656 61816
rect 72622 60950 72656 61122
rect 72622 60256 72656 60428
rect 72622 59562 72656 59734
rect 72622 58868 72656 59040
rect 73280 61644 73314 61816
rect 79678 62626 79712 62798
rect 80336 65402 80370 65574
rect 80336 64708 80370 64880
rect 80336 64014 80370 64186
rect 80336 63320 80370 63492
rect 80336 62626 80370 62798
rect 80994 65402 81028 65574
rect 80994 64708 81028 64880
rect 80994 64014 81028 64186
rect 80994 63320 81028 63492
rect 80994 62626 81028 62798
rect 81652 65402 81686 65574
rect 81652 64708 81686 64880
rect 81652 64014 81686 64186
rect 81652 63320 81686 63492
rect 81652 62626 81686 62798
rect 73280 60950 73314 61122
rect 73280 60256 73314 60428
rect 73280 59562 73314 59734
rect 73280 58868 73314 59040
rect 73938 61644 73972 61816
rect 73938 60950 73972 61122
rect 73938 60256 73972 60428
rect 73938 59562 73972 59734
rect 73938 58868 73972 59040
rect 74926 59082 75010 61650
rect 75170 61624 75204 61796
rect 75170 60930 75204 61102
rect 75170 60236 75204 60408
rect 75170 59542 75204 59714
rect 75828 61624 75862 61796
rect 75828 60930 75862 61102
rect 75828 60236 75862 60408
rect 75828 59542 75862 59714
rect 75170 58848 75204 59020
rect 54420 57692 54592 57726
rect 55114 57692 55286 57726
rect 55808 57692 55980 57726
rect 56502 57692 56674 57726
rect 57196 57692 57368 57726
rect 42382 57034 42554 57068
rect 43076 57034 43248 57068
rect 43770 57034 43942 57068
rect 44464 57034 44636 57068
rect 45158 57034 45330 57068
rect 46376 57034 46548 57068
rect 47070 57034 47242 57068
rect 47764 57034 47936 57068
rect 48458 57034 48630 57068
rect 49152 57034 49324 57068
rect 50398 57034 50570 57068
rect 51092 57034 51264 57068
rect 51786 57034 51958 57068
rect 52480 57034 52652 57068
rect 53174 57034 53346 57068
rect 54420 57034 54592 57068
rect 55114 57034 55286 57068
rect 55808 57034 55980 57068
rect 56502 57034 56674 57068
rect 57196 57034 57368 57068
rect 23634 56788 23806 56822
rect 24328 56788 24500 56822
rect 25022 56788 25194 56822
rect 25716 56788 25888 56822
rect 26410 56788 26582 56822
rect 27104 56788 27276 56822
rect 27798 56788 27970 56822
rect 28492 56788 28664 56822
rect 29186 56788 29358 56822
rect 29880 56788 30052 56822
rect 19544 56686 19716 56720
rect 20238 56686 20410 56720
rect 19544 56028 19716 56062
rect 20238 56028 20410 56062
rect 16860 55326 17032 55360
rect 17554 55326 17726 55360
rect 18248 55326 18420 55360
rect 16860 54668 17032 54702
rect 17554 54668 17726 54702
rect 18248 54668 18420 54702
rect 18844 54548 19054 54894
rect 30348 56782 30386 56840
rect 58868 56840 59184 57288
rect 23634 56130 23806 56164
rect 24328 56130 24500 56164
rect 25022 56130 25194 56164
rect 25716 56130 25888 56164
rect 26410 56130 26582 56164
rect 27104 56130 27276 56164
rect 27798 56130 27970 56164
rect 28492 56130 28664 56164
rect 29186 56130 29358 56164
rect 29880 56130 30052 56164
rect 42976 56218 45150 56420
rect 46984 56216 49158 56418
rect 50996 56216 53170 56418
rect 55006 56216 57180 56418
rect 24408 55788 25052 55844
rect 28824 55902 29468 55946
rect 42334 55934 42506 55968
rect 43028 55934 43200 55968
rect 43722 55934 43894 55968
rect 44416 55934 44588 55968
rect 45110 55934 45282 55968
rect 46342 55932 46514 55966
rect 47036 55932 47208 55966
rect 47730 55932 47902 55966
rect 48424 55932 48596 55966
rect 49118 55932 49290 55966
rect 50354 55932 50526 55966
rect 51048 55932 51220 55966
rect 51742 55932 51914 55966
rect 52436 55932 52608 55966
rect 53130 55932 53302 55966
rect 54364 55932 54536 55966
rect 55058 55932 55230 55966
rect 55752 55932 55924 55966
rect 56446 55932 56618 55966
rect 57140 55932 57312 55966
rect 23640 55556 23812 55590
rect 24334 55556 24506 55590
rect 25028 55556 25200 55590
rect 25722 55556 25894 55590
rect 26416 55556 26588 55590
rect 27110 55556 27282 55590
rect 27804 55556 27976 55590
rect 28498 55556 28670 55590
rect 29192 55556 29364 55590
rect 29886 55556 30058 55590
rect 19544 55370 19716 55404
rect 20238 55370 20410 55404
rect 19544 54712 19716 54746
rect 20238 54712 20410 54746
rect 23006 55000 23088 55346
rect 23640 54898 23812 54932
rect 24334 54898 24506 54932
rect 25028 54898 25200 54932
rect 25722 54898 25894 54932
rect 26416 54898 26588 54932
rect 27110 54898 27282 54932
rect 27804 54898 27976 54932
rect 28498 54898 28670 54932
rect 29192 54898 29364 54932
rect 29886 54898 30058 54932
rect 20690 54456 20770 54624
rect 23316 54452 23374 54720
rect 23640 54240 23812 54274
rect 24334 54240 24506 54274
rect 25028 54240 25200 54274
rect 25722 54240 25894 54274
rect 26416 54240 26588 54274
rect 27110 54240 27282 54274
rect 27804 54240 27976 54274
rect 28498 54240 28670 54274
rect 29192 54240 29364 54274
rect 29886 54240 30058 54274
rect 42334 55276 42506 55310
rect 43028 55276 43200 55310
rect 43722 55276 43894 55310
rect 44416 55276 44588 55310
rect 45110 55276 45282 55310
rect 19544 54054 19716 54088
rect 20238 54054 20410 54088
rect 938 54004 1110 54038
rect 1632 54004 1804 54038
rect 2326 54004 2498 54038
rect 3606 54000 3778 54034
rect 4300 54000 4472 54034
rect 4994 54000 5166 54034
rect 6280 54006 6452 54040
rect 6974 54006 7146 54040
rect 7668 54006 7840 54040
rect 8926 54006 9098 54040
rect 9620 54006 9792 54040
rect 10314 54006 10486 54040
rect 11580 54000 11752 54034
rect 12274 54000 12446 54034
rect 12968 54000 13140 54034
rect 14234 54006 14406 54040
rect 14928 54006 15100 54040
rect 15622 54006 15794 54040
rect 16860 54010 17032 54044
rect 17554 54010 17726 54044
rect 18248 54010 18420 54044
rect 24414 53898 25058 53954
rect 28830 54012 29474 54056
rect 46342 55274 46514 55308
rect 47036 55274 47208 55308
rect 47730 55274 47902 55308
rect 48424 55274 48596 55308
rect 49118 55274 49290 55308
rect 42334 54618 42506 54652
rect 43028 54618 43200 54652
rect 43722 54618 43894 54652
rect 44416 54618 44588 54652
rect 45110 54618 45282 54652
rect 42334 53960 42506 53994
rect 43028 53960 43200 53994
rect 43722 53960 43894 53994
rect 44416 53960 44588 53994
rect 45110 53960 45282 53994
rect 23656 53614 23828 53648
rect 24350 53614 24522 53648
rect 25044 53614 25216 53648
rect 25738 53614 25910 53648
rect 26432 53614 26604 53648
rect 27126 53614 27298 53648
rect 27820 53614 27992 53648
rect 28514 53614 28686 53648
rect 29208 53614 29380 53648
rect 29902 53614 30074 53648
rect 1058 53200 2462 53270
rect 3726 53196 5130 53266
rect 6400 53202 7804 53272
rect 9046 53202 10450 53272
rect 11700 53196 13104 53266
rect 14354 53202 15758 53272
rect 16980 53206 18384 53276
rect 19534 53182 20492 53290
rect 19544 52952 19716 52986
rect 20238 52952 20410 52986
rect 938 52902 1110 52936
rect 1632 52902 1804 52936
rect 2326 52902 2498 52936
rect 3606 52898 3778 52932
rect 4300 52898 4472 52932
rect 4994 52898 5166 52932
rect 6280 52904 6452 52938
rect 6974 52904 7146 52938
rect 7668 52904 7840 52938
rect 8926 52904 9098 52938
rect 9620 52904 9792 52938
rect 10314 52904 10486 52938
rect 11580 52898 11752 52932
rect 12274 52898 12446 52932
rect 12968 52898 13140 52932
rect 14234 52904 14406 52938
rect 14928 52904 15100 52938
rect 15622 52904 15794 52938
rect 16860 52908 17032 52942
rect 17554 52908 17726 52942
rect 18248 52908 18420 52942
rect 23656 52956 23828 52990
rect 24350 52956 24522 52990
rect 25044 52956 25216 52990
rect 25738 52956 25910 52990
rect 26432 52956 26604 52990
rect 27126 52956 27298 52990
rect 27820 52956 27992 52990
rect 28514 52956 28686 52990
rect 29208 52956 29380 52990
rect 29902 52956 30074 52990
rect 30390 52964 30444 53048
rect 938 52244 1110 52278
rect 1632 52244 1804 52278
rect 2326 52244 2498 52278
rect 938 51586 1110 51620
rect 1632 51586 1804 51620
rect 2326 51586 2498 51620
rect 938 50928 1110 50962
rect 1632 50928 1804 50962
rect 2326 50928 2498 50962
rect 938 50270 1110 50304
rect 1632 50270 1804 50304
rect 2326 50270 2498 50304
rect 938 49612 1110 49646
rect 1632 49612 1804 49646
rect 2326 49612 2498 49646
rect 3606 52240 3778 52274
rect 4300 52240 4472 52274
rect 4994 52240 5166 52274
rect 3606 51582 3778 51616
rect 4300 51582 4472 51616
rect 4994 51582 5166 51616
rect 3606 50924 3778 50958
rect 4300 50924 4472 50958
rect 4994 50924 5166 50958
rect 3606 50266 3778 50300
rect 4300 50266 4472 50300
rect 4994 50266 5166 50300
rect 3606 49608 3778 49642
rect 4300 49608 4472 49642
rect 4994 49608 5166 49642
rect 938 48954 1110 48988
rect 1632 48954 1804 48988
rect 2326 48954 2498 48988
rect 938 48296 1110 48330
rect 1632 48296 1804 48330
rect 2326 48296 2498 48330
rect 3058 48082 3276 48436
rect 6280 52246 6452 52280
rect 6974 52246 7146 52280
rect 7668 52246 7840 52280
rect 6280 51588 6452 51622
rect 6974 51588 7146 51622
rect 7668 51588 7840 51622
rect 6280 50930 6452 50964
rect 6974 50930 7146 50964
rect 7668 50930 7840 50964
rect 6280 50272 6452 50306
rect 6974 50272 7146 50306
rect 7668 50272 7840 50306
rect 6280 49614 6452 49648
rect 6974 49614 7146 49648
rect 7668 49614 7840 49648
rect 3606 48950 3778 48984
rect 4300 48950 4472 48984
rect 4994 48950 5166 48984
rect 3606 48292 3778 48326
rect 4300 48292 4472 48326
rect 4994 48292 5166 48326
rect 5692 48108 5928 48470
rect 8926 52246 9098 52280
rect 9620 52246 9792 52280
rect 10314 52246 10486 52280
rect 8926 51588 9098 51622
rect 9620 51588 9792 51622
rect 10314 51588 10486 51622
rect 8926 50930 9098 50964
rect 9620 50930 9792 50964
rect 10314 50930 10486 50964
rect 8926 50272 9098 50306
rect 9620 50272 9792 50306
rect 10314 50272 10486 50306
rect 8926 49614 9098 49648
rect 9620 49614 9792 49648
rect 10314 49614 10486 49648
rect 6280 48956 6452 48990
rect 6974 48956 7146 48990
rect 7668 48956 7840 48990
rect 6280 48298 6452 48332
rect 6974 48298 7146 48332
rect 7668 48298 7840 48332
rect 8352 48058 8554 48546
rect 11580 52240 11752 52274
rect 12274 52240 12446 52274
rect 12968 52240 13140 52274
rect 11580 51582 11752 51616
rect 12274 51582 12446 51616
rect 12968 51582 13140 51616
rect 11580 50924 11752 50958
rect 12274 50924 12446 50958
rect 12968 50924 13140 50958
rect 11580 50266 11752 50300
rect 12274 50266 12446 50300
rect 12968 50266 13140 50300
rect 11580 49608 11752 49642
rect 12274 49608 12446 49642
rect 12968 49608 13140 49642
rect 8926 48956 9098 48990
rect 9620 48956 9792 48990
rect 10314 48956 10486 48990
rect 8926 48298 9098 48332
rect 9620 48298 9792 48332
rect 10314 48298 10486 48332
rect 11028 48024 11246 48462
rect 14234 52246 14406 52280
rect 14928 52246 15100 52280
rect 15622 52246 15794 52280
rect 14234 51588 14406 51622
rect 14928 51588 15100 51622
rect 15622 51588 15794 51622
rect 14234 50930 14406 50964
rect 14928 50930 15100 50964
rect 15622 50930 15794 50964
rect 14234 50272 14406 50306
rect 14928 50272 15100 50306
rect 15622 50272 15794 50306
rect 14234 49614 14406 49648
rect 14928 49614 15100 49648
rect 15622 49614 15794 49648
rect 11580 48950 11752 48984
rect 12274 48950 12446 48984
rect 12968 48950 13140 48984
rect 11580 48292 11752 48326
rect 12274 48292 12446 48326
rect 12968 48292 13140 48326
rect 13678 48066 13846 48494
rect 16860 52250 17032 52284
rect 17554 52250 17726 52284
rect 18248 52250 18420 52284
rect 19544 52294 19716 52328
rect 20238 52294 20410 52328
rect 16860 51592 17032 51626
rect 17554 51592 17726 51626
rect 18248 51592 18420 51626
rect 16860 50934 17032 50968
rect 17554 50934 17726 50968
rect 18248 50934 18420 50968
rect 16860 50276 17032 50310
rect 17554 50276 17726 50310
rect 18248 50276 18420 50310
rect 16860 49618 17032 49652
rect 17554 49618 17726 49652
rect 18248 49618 18420 49652
rect 14234 48956 14406 48990
rect 14928 48956 15100 48990
rect 15622 48956 15794 48990
rect 14234 48298 14406 48332
rect 14928 48298 15100 48332
rect 15622 48298 15794 48332
rect 16294 48166 16548 48436
rect 50354 55274 50526 55308
rect 51048 55274 51220 55308
rect 51742 55274 51914 55308
rect 52436 55274 52608 55308
rect 53130 55274 53302 55308
rect 46342 54616 46514 54650
rect 47036 54616 47208 54650
rect 47730 54616 47902 54650
rect 48424 54616 48596 54650
rect 49118 54616 49290 54650
rect 46342 53958 46514 53992
rect 47036 53958 47208 53992
rect 47730 53958 47902 53992
rect 48424 53958 48596 53992
rect 49118 53958 49290 53992
rect 42334 53302 42506 53336
rect 43028 53302 43200 53336
rect 43722 53302 43894 53336
rect 44416 53302 44588 53336
rect 45110 53302 45282 53336
rect 23656 52298 23828 52332
rect 24350 52298 24522 52332
rect 25044 52298 25216 52332
rect 25738 52298 25910 52332
rect 26432 52298 26604 52332
rect 27126 52298 27298 52332
rect 27820 52298 27992 52332
rect 28514 52298 28686 52332
rect 29208 52298 29380 52332
rect 29902 52298 30074 52332
rect 54364 55274 54536 55308
rect 55058 55274 55230 55308
rect 55752 55274 55924 55308
rect 56446 55274 56618 55308
rect 57140 55274 57312 55308
rect 50354 54616 50526 54650
rect 51048 54616 51220 54650
rect 51742 54616 51914 54650
rect 52436 54616 52608 54650
rect 53130 54616 53302 54650
rect 50354 53958 50526 53992
rect 51048 53958 51220 53992
rect 51742 53958 51914 53992
rect 52436 53958 52608 53992
rect 53130 53958 53302 53992
rect 46342 53300 46514 53334
rect 47036 53300 47208 53334
rect 47730 53300 47902 53334
rect 48424 53300 48596 53334
rect 49118 53300 49290 53334
rect 54364 54616 54536 54650
rect 55058 54616 55230 54650
rect 55752 54616 55924 54650
rect 56446 54616 56618 54650
rect 57140 54616 57312 54650
rect 54364 53958 54536 53992
rect 55058 53958 55230 53992
rect 55752 53958 55924 53992
rect 56446 53958 56618 53992
rect 57140 53958 57312 53992
rect 50354 53300 50526 53334
rect 51048 53300 51220 53334
rect 51742 53300 51914 53334
rect 52436 53300 52608 53334
rect 53130 53300 53302 53334
rect 54364 53300 54536 53334
rect 55058 53300 55230 53334
rect 55752 53300 55924 53334
rect 56446 53300 56618 53334
rect 57140 53300 57312 53334
rect 42334 52644 42506 52678
rect 43028 52644 43200 52678
rect 43722 52644 43894 52678
rect 44416 52644 44588 52678
rect 45110 52644 45282 52678
rect 46342 52642 46514 52676
rect 47036 52642 47208 52676
rect 47730 52642 47902 52676
rect 48424 52642 48596 52676
rect 49118 52642 49290 52676
rect 50354 52642 50526 52676
rect 51048 52642 51220 52676
rect 51742 52642 51914 52676
rect 52436 52642 52608 52676
rect 53130 52642 53302 52676
rect 54364 52642 54536 52676
rect 55058 52642 55230 52676
rect 55752 52642 55924 52676
rect 56446 52642 56618 52676
rect 57140 52642 57312 52676
rect 24430 51956 25074 52012
rect 28846 52070 29490 52114
rect 19544 51636 19716 51670
rect 20238 51636 20410 51670
rect 19544 50978 19716 51012
rect 20238 50978 20410 51012
rect 19544 50320 19716 50354
rect 20238 50320 20410 50354
rect 19544 49662 19716 49696
rect 20238 49662 20410 49696
rect 16860 48960 17032 48994
rect 17554 48960 17726 48994
rect 18248 48960 18420 48994
rect 16860 48302 17032 48336
rect 17554 48302 17726 48336
rect 18248 48302 18420 48336
rect 18844 48182 19054 48528
rect 19544 49004 19716 49038
rect 20238 49004 20410 49038
rect 20690 48694 20742 48728
rect 19544 48346 19716 48380
rect 20238 48346 20410 48380
rect 19544 47688 19716 47722
rect 20238 47688 20410 47722
rect 938 47638 1110 47672
rect 1632 47638 1804 47672
rect 2326 47638 2498 47672
rect 3606 47634 3778 47668
rect 4300 47634 4472 47668
rect 4994 47634 5166 47668
rect 6280 47640 6452 47674
rect 6974 47640 7146 47674
rect 7668 47640 7840 47674
rect 8926 47640 9098 47674
rect 9620 47640 9792 47674
rect 10314 47640 10486 47674
rect 11580 47634 11752 47668
rect 12274 47634 12446 47668
rect 12968 47634 13140 47668
rect 14234 47640 14406 47674
rect 14928 47640 15100 47674
rect 15622 47640 15794 47674
rect 16860 47644 17032 47678
rect 17554 47644 17726 47678
rect 18248 47644 18420 47678
rect 2730 47258 4298 47334
rect 9218 47266 10514 47394
rect 14392 47244 15472 47360
rect 17118 47292 18328 47394
rect 19582 47256 20426 47364
rect 42968 52020 45142 52222
rect 46962 52020 49136 52222
rect 50984 52020 53158 52222
rect 55006 52020 57180 52222
rect 57636 52026 57760 52328
rect 42326 51736 42498 51770
rect 43020 51736 43192 51770
rect 43714 51736 43886 51770
rect 44408 51736 44580 51770
rect 45102 51736 45274 51770
rect 46320 51736 46492 51770
rect 47014 51736 47186 51770
rect 47708 51736 47880 51770
rect 48402 51736 48574 51770
rect 49096 51736 49268 51770
rect 50342 51736 50514 51770
rect 51036 51736 51208 51770
rect 51730 51736 51902 51770
rect 52424 51736 52596 51770
rect 53118 51736 53290 51770
rect 54364 51736 54536 51770
rect 55058 51736 55230 51770
rect 55752 51736 55924 51770
rect 56446 51736 56618 51770
rect 57140 51736 57312 51770
rect 42326 51078 42498 51112
rect 43020 51078 43192 51112
rect 43714 51078 43886 51112
rect 44408 51078 44580 51112
rect 45102 51078 45274 51112
rect 46320 51078 46492 51112
rect 47014 51078 47186 51112
rect 47708 51078 47880 51112
rect 48402 51078 48574 51112
rect 49096 51078 49268 51112
rect 42326 50420 42498 50454
rect 43020 50420 43192 50454
rect 43714 50420 43886 50454
rect 44408 50420 44580 50454
rect 45102 50420 45274 50454
rect 42326 49762 42498 49796
rect 43020 49762 43192 49796
rect 43714 49762 43886 49796
rect 44408 49762 44580 49796
rect 45102 49762 45274 49796
rect 50342 51078 50514 51112
rect 51036 51078 51208 51112
rect 51730 51078 51902 51112
rect 52424 51078 52596 51112
rect 53118 51078 53290 51112
rect 46320 50420 46492 50454
rect 47014 50420 47186 50454
rect 47708 50420 47880 50454
rect 48402 50420 48574 50454
rect 49096 50420 49268 50454
rect 46320 49762 46492 49796
rect 47014 49762 47186 49796
rect 47708 49762 47880 49796
rect 48402 49762 48574 49796
rect 49096 49762 49268 49796
rect 42326 49104 42498 49138
rect 43020 49104 43192 49138
rect 43714 49104 43886 49138
rect 44408 49104 44580 49138
rect 45102 49104 45274 49138
rect 54364 51078 54536 51112
rect 55058 51078 55230 51112
rect 55752 51078 55924 51112
rect 56446 51078 56618 51112
rect 57140 51078 57312 51112
rect 50342 50420 50514 50454
rect 51036 50420 51208 50454
rect 51730 50420 51902 50454
rect 52424 50420 52596 50454
rect 53118 50420 53290 50454
rect 50342 49762 50514 49796
rect 51036 49762 51208 49796
rect 51730 49762 51902 49796
rect 52424 49762 52596 49796
rect 53118 49762 53290 49796
rect 46320 49104 46492 49138
rect 47014 49104 47186 49138
rect 47708 49104 47880 49138
rect 48402 49104 48574 49138
rect 49096 49104 49268 49138
rect 54364 50420 54536 50454
rect 55058 50420 55230 50454
rect 55752 50420 55924 50454
rect 56446 50420 56618 50454
rect 57140 50420 57312 50454
rect 54364 49762 54536 49796
rect 55058 49762 55230 49796
rect 55752 49762 55924 49796
rect 56446 49762 56618 49796
rect 57140 49762 57312 49796
rect 50342 49104 50514 49138
rect 51036 49104 51208 49138
rect 51730 49104 51902 49138
rect 52424 49104 52596 49138
rect 53118 49104 53290 49138
rect 54364 49104 54536 49138
rect 55058 49104 55230 49138
rect 55752 49104 55924 49138
rect 56446 49104 56618 49138
rect 57140 49104 57312 49138
rect 42326 48446 42498 48480
rect 43020 48446 43192 48480
rect 43714 48446 43886 48480
rect 44408 48446 44580 48480
rect 45102 48446 45274 48480
rect 46320 48446 46492 48480
rect 47014 48446 47186 48480
rect 47708 48446 47880 48480
rect 48402 48446 48574 48480
rect 49096 48446 49268 48480
rect 50342 48446 50514 48480
rect 51036 48446 51208 48480
rect 51730 48446 51902 48480
rect 52424 48446 52596 48480
rect 53118 48446 53290 48480
rect 54364 48446 54536 48480
rect 55058 48446 55230 48480
rect 55752 48446 55924 48480
rect 56446 48446 56618 48480
rect 57140 48446 57312 48480
rect 42872 47994 44786 48112
rect 46870 47968 49234 48126
rect 50844 47954 53232 48086
rect 54540 47954 57088 48140
rect 71062 55326 71146 57894
rect 71306 57868 71340 58040
rect 71306 57174 71340 57346
rect 71306 56480 71340 56652
rect 71306 55786 71340 55958
rect 71964 57868 71998 58040
rect 75828 58848 75862 59020
rect 76486 61624 76520 61796
rect 76486 60930 76520 61102
rect 76486 60236 76520 60408
rect 76486 59542 76520 59714
rect 76486 58848 76520 59020
rect 77144 61624 77178 61796
rect 77144 60930 77178 61102
rect 77144 60236 77178 60408
rect 77144 59542 77178 59714
rect 77144 58848 77178 59020
rect 77802 61624 77836 61796
rect 77802 60930 77836 61102
rect 77802 60236 77836 60408
rect 77802 59542 77836 59714
rect 77802 58848 77836 59020
rect 78776 59096 78860 61664
rect 79020 61638 79054 61810
rect 79020 60944 79054 61116
rect 79020 60250 79054 60422
rect 79020 59556 79054 59728
rect 79678 61638 79712 61810
rect 79678 60944 79712 61116
rect 79678 60250 79712 60422
rect 79678 59556 79712 59728
rect 79020 58862 79054 59034
rect 71964 57174 71998 57346
rect 71964 56480 71998 56652
rect 71964 55786 71998 55958
rect 71306 55092 71340 55264
rect 71964 55092 71998 55264
rect 72622 57868 72656 58040
rect 72622 57174 72656 57346
rect 72622 56480 72656 56652
rect 72622 55786 72656 55958
rect 72622 55092 72656 55264
rect 73280 57868 73314 58040
rect 73280 57174 73314 57346
rect 73280 56480 73314 56652
rect 73280 55786 73314 55958
rect 73280 55092 73314 55264
rect 73938 57868 73972 58040
rect 73938 57174 73972 57346
rect 73938 56480 73972 56652
rect 73938 55786 73972 55958
rect 73938 55092 73972 55264
rect 74926 55306 75010 57874
rect 75170 57848 75204 58020
rect 75170 57154 75204 57326
rect 75170 56460 75204 56632
rect 75170 55766 75204 55938
rect 75828 57848 75862 58020
rect 79678 58862 79712 59034
rect 80336 61638 80370 61810
rect 80336 60944 80370 61116
rect 80336 60250 80370 60422
rect 80336 59556 80370 59728
rect 80336 58862 80370 59034
rect 80994 61638 81028 61810
rect 80994 60944 81028 61116
rect 80994 60250 81028 60422
rect 80994 59556 81028 59728
rect 80994 58862 81028 59034
rect 81652 61638 81686 61810
rect 81652 60944 81686 61116
rect 81652 60250 81686 60422
rect 81652 59556 81686 59728
rect 81652 58862 81686 59034
rect 75828 57154 75862 57326
rect 75828 56460 75862 56632
rect 75828 55766 75862 55938
rect 75170 55072 75204 55244
rect 75828 55072 75862 55244
rect 76486 57848 76520 58020
rect 76486 57154 76520 57326
rect 76486 56460 76520 56632
rect 76486 55766 76520 55938
rect 76486 55072 76520 55244
rect 77144 57848 77178 58020
rect 77144 57154 77178 57326
rect 77144 56460 77178 56632
rect 77144 55766 77178 55938
rect 77144 55072 77178 55244
rect 77802 57848 77836 58020
rect 77802 57154 77836 57326
rect 77802 56460 77836 56632
rect 77802 55766 77836 55938
rect 77802 55072 77836 55244
rect 78776 55320 78860 57888
rect 79020 57862 79054 58034
rect 79020 57168 79054 57340
rect 79020 56474 79054 56646
rect 79020 55780 79054 55952
rect 79678 57862 79712 58034
rect 79678 57168 79712 57340
rect 79678 56474 79712 56646
rect 79678 55780 79712 55952
rect 79020 55086 79054 55258
rect 79678 55086 79712 55258
rect 80336 57862 80370 58034
rect 80336 57168 80370 57340
rect 80336 56474 80370 56646
rect 80336 55780 80370 55952
rect 80336 55086 80370 55258
rect 80994 57862 81028 58034
rect 80994 57168 81028 57340
rect 80994 56474 81028 56646
rect 80994 55780 81028 55952
rect 80994 55086 81028 55258
rect 81652 57862 81686 58034
rect 81652 57168 81686 57340
rect 81652 56474 81686 56646
rect 81652 55780 81686 55952
rect 81652 55086 81686 55258
rect 71066 51554 71150 54122
rect 71310 54096 71344 54268
rect 71310 53402 71344 53574
rect 71310 52708 71344 52880
rect 71310 52014 71344 52186
rect 71310 51320 71344 51492
rect 71968 54096 72002 54268
rect 71968 53402 72002 53574
rect 71968 52708 72002 52880
rect 71968 52014 72002 52186
rect 71968 51320 72002 51492
rect 72626 54096 72660 54268
rect 72626 53402 72660 53574
rect 72626 52708 72660 52880
rect 72626 52014 72660 52186
rect 72626 51320 72660 51492
rect 73284 54096 73318 54268
rect 73284 53402 73318 53574
rect 73284 52708 73318 52880
rect 73284 52014 73318 52186
rect 73284 51320 73318 51492
rect 73942 54096 73976 54268
rect 73942 53402 73976 53574
rect 73942 52708 73976 52880
rect 73942 52014 73976 52186
rect 73942 51320 73976 51492
rect 74930 51534 75014 54102
rect 75174 54076 75208 54248
rect 75174 53382 75208 53554
rect 75174 52688 75208 52860
rect 75174 51994 75208 52166
rect 75174 51300 75208 51472
rect 75832 54076 75866 54248
rect 75832 53382 75866 53554
rect 75832 52688 75866 52860
rect 75832 51994 75866 52166
rect 75832 51300 75866 51472
rect 76490 54076 76524 54248
rect 76490 53382 76524 53554
rect 76490 52688 76524 52860
rect 76490 51994 76524 52166
rect 76490 51300 76524 51472
rect 77148 54076 77182 54248
rect 77148 53382 77182 53554
rect 77148 52688 77182 52860
rect 77148 51994 77182 52166
rect 77148 51300 77182 51472
rect 77806 54076 77840 54248
rect 77806 53382 77840 53554
rect 77806 52688 77840 52860
rect 77806 51994 77840 52166
rect 77806 51300 77840 51472
rect 78780 51548 78864 54116
rect 79024 54090 79058 54262
rect 79024 53396 79058 53568
rect 79024 52702 79058 52874
rect 79024 52008 79058 52180
rect 79024 51314 79058 51486
rect 79682 54090 79716 54262
rect 79682 53396 79716 53568
rect 79682 52702 79716 52874
rect 79682 52008 79716 52180
rect 79682 51314 79716 51486
rect 80340 54090 80374 54262
rect 80340 53396 80374 53568
rect 80340 52702 80374 52874
rect 80340 52008 80374 52180
rect 80340 51314 80374 51486
rect 80998 54090 81032 54262
rect 80998 53396 81032 53568
rect 80998 52702 81032 52874
rect 80998 52008 81032 52180
rect 80998 51314 81032 51486
rect 81656 54090 81690 54262
rect 81924 54218 82048 54890
rect 83303 54065 83337 54099
rect 83399 54065 83433 54099
rect 83495 54065 83529 54099
rect 83591 54065 83625 54099
rect 83687 54065 83721 54099
rect 83783 54065 83817 54099
rect 83879 54065 83913 54099
rect 83975 54065 84009 54099
rect 84071 54065 84105 54099
rect 84167 54065 84201 54099
rect 84263 54065 84297 54099
rect 84359 54065 84393 54099
rect 84455 54065 84489 54099
rect 84551 54065 84585 54099
rect 84647 54065 84681 54099
rect 84743 54065 84777 54099
rect 84839 54065 84873 54099
rect 84935 54065 84969 54099
rect 85031 54065 85065 54099
rect 85127 54065 85161 54099
rect 85223 54065 85257 54099
rect 85319 54065 85353 54099
rect 85415 54065 85449 54099
rect 85511 54065 85545 54099
rect 85607 54065 85641 54099
rect 85703 54065 85737 54099
rect 85799 54065 85833 54099
rect 85895 54065 85929 54099
rect 85991 54065 86025 54099
rect 86087 54065 86121 54099
rect 86183 54065 86217 54099
rect 86279 54065 86313 54099
rect 83404 53969 83438 54003
rect 83476 53969 83510 54003
rect 81656 53396 81690 53568
rect 83382 53640 83448 53700
rect 83882 53976 83916 54003
rect 83882 53969 83892 53976
rect 83892 53969 83916 53976
rect 83687 53658 83721 53692
rect 83390 53347 83424 53381
rect 83462 53347 83496 53381
rect 83534 53347 83568 53381
rect 83970 53605 84020 53606
rect 83970 53571 83971 53605
rect 83971 53571 84005 53605
rect 84005 53571 84020 53605
rect 83970 53550 84020 53571
rect 83870 53460 83920 53498
rect 83718 53347 83752 53381
rect 83790 53347 83824 53381
rect 84368 53969 84402 54003
rect 84440 53969 84474 54003
rect 84512 53969 84546 54003
rect 84836 53998 84870 54003
rect 84836 53969 84846 53998
rect 84846 53969 84870 53998
rect 84908 53969 84942 54003
rect 84980 53969 85014 54003
rect 84167 53658 84201 53692
rect 84710 53347 84744 53381
rect 84782 53347 84816 53381
rect 84854 53347 84888 53381
rect 85375 53969 85409 54003
rect 85447 53969 85481 54003
rect 85519 53969 85553 54003
rect 85726 53969 85760 54003
rect 85798 53969 85832 54003
rect 85870 53969 85904 54003
rect 86032 53969 86066 54003
rect 86104 53999 86138 54003
rect 86104 53969 86116 53999
rect 86116 53969 86138 53999
rect 86176 53969 86210 54003
rect 85223 53658 85257 53692
rect 86270 53586 86316 53630
rect 85504 53347 85538 53381
rect 85576 53347 85610 53381
rect 85648 53347 85682 53381
rect 86025 53347 86059 53381
rect 86097 53347 86131 53381
rect 86169 53347 86203 53381
rect 83303 53251 83337 53285
rect 83399 53251 83433 53285
rect 83495 53251 83529 53285
rect 83591 53251 83625 53285
rect 83687 53251 83721 53285
rect 83783 53251 83817 53285
rect 83879 53251 83913 53285
rect 83975 53251 84009 53285
rect 84071 53251 84105 53285
rect 84167 53251 84201 53285
rect 84263 53251 84297 53285
rect 84359 53251 84393 53285
rect 84455 53251 84489 53285
rect 84551 53251 84585 53285
rect 84647 53251 84681 53285
rect 84743 53251 84777 53285
rect 84839 53251 84873 53285
rect 84935 53251 84969 53285
rect 85031 53251 85065 53285
rect 85127 53251 85161 53285
rect 85223 53251 85257 53285
rect 85319 53251 85353 53285
rect 85415 53251 85449 53285
rect 85511 53251 85545 53285
rect 85607 53251 85641 53285
rect 85703 53251 85737 53285
rect 85799 53251 85833 53285
rect 85895 53251 85929 53285
rect 85991 53251 86025 53285
rect 86087 53251 86121 53285
rect 86183 53251 86217 53285
rect 86279 53251 86313 53285
rect 81656 52702 81690 52874
rect 81656 52008 81690 52180
rect 81656 51314 81690 51486
rect 77384 50850 77634 51008
rect 75734 48226 76396 48690
rect 66184 46248 66696 46524
rect 24382 44696 25184 44984
rect 39408 44424 41694 45004
rect 11074 43646 11216 43708
rect 1958 42760 1992 43052
rect 1958 41666 1992 41958
rect 1326 40322 1420 41518
rect 1958 40572 1992 40864
rect 1958 39478 1992 39770
rect 1958 38384 1992 38676
rect 3016 42760 3050 43052
rect 3016 41666 3050 41958
rect 3016 40572 3050 40864
rect 3016 39478 3050 39770
rect 3016 38384 3050 38676
rect 4074 42760 4108 43052
rect 4074 41666 4108 41958
rect 4074 40572 4108 40864
rect 4074 39478 4108 39770
rect 4074 38384 4108 38676
rect 5132 42760 5166 43052
rect 5132 41666 5166 41958
rect 5132 40572 5166 40864
rect 5132 39478 5166 39770
rect 5132 38384 5166 38676
rect 6190 42760 6224 43052
rect 6190 41666 6224 41958
rect 6190 40572 6224 40864
rect 6190 39478 6224 39770
rect 6190 38384 6224 38676
rect 7248 42760 7282 43052
rect 7248 41666 7282 41958
rect 8472 42768 8506 43060
rect 8472 41674 8506 41966
rect 7248 40572 7282 40864
rect 7840 40330 7934 41526
rect 8472 40580 8506 40872
rect 7248 39478 7282 39770
rect 7248 38384 7282 38676
rect 8472 39486 8506 39778
rect 8472 38392 8506 38684
rect 9530 42768 9564 43060
rect 9530 41674 9564 41966
rect 9530 40580 9564 40872
rect 9530 39486 9564 39778
rect 1958 36944 1992 37236
rect 1958 35850 1992 36142
rect 1326 34506 1420 35702
rect 1958 34756 1992 35048
rect 1958 33662 1992 33954
rect 1958 32568 1992 32860
rect 3016 36944 3050 37236
rect 3016 35850 3050 36142
rect 3016 34756 3050 35048
rect 3016 33662 3050 33954
rect 3016 32568 3050 32860
rect 4074 36944 4108 37236
rect 4074 35850 4108 36142
rect 4074 34756 4108 35048
rect 4074 33662 4108 33954
rect 4074 32568 4108 32860
rect 5132 36944 5166 37236
rect 5132 35850 5166 36142
rect 5132 34756 5166 35048
rect 5132 33662 5166 33954
rect 5132 32568 5166 32860
rect 6190 36944 6224 37236
rect 9530 38392 9564 38684
rect 10588 42768 10622 43060
rect 10588 41674 10622 41966
rect 10588 40580 10622 40872
rect 10588 39486 10622 39778
rect 10588 38392 10622 38684
rect 11646 42768 11680 43060
rect 11646 41674 11680 41966
rect 11646 40580 11680 40872
rect 11646 39486 11680 39778
rect 11646 38392 11680 38684
rect 12704 42768 12738 43060
rect 12704 41674 12738 41966
rect 12704 40580 12738 40872
rect 12704 39486 12738 39778
rect 12704 38392 12738 38684
rect 13762 42768 13796 43060
rect 13762 41674 13796 41966
rect 14978 42776 15012 43068
rect 14978 41682 15012 41974
rect 13762 40580 13796 40872
rect 14346 40338 14440 41534
rect 14978 40588 15012 40880
rect 13762 39486 13796 39778
rect 13762 38392 13796 38684
rect 14978 39494 15012 39786
rect 14978 38400 15012 38692
rect 16036 42776 16070 43068
rect 16036 41682 16070 41974
rect 16036 40588 16070 40880
rect 16036 39494 16070 39786
rect 6190 35850 6224 36142
rect 6190 34756 6224 35048
rect 6190 33662 6224 33954
rect 6190 32568 6224 32860
rect 7248 36944 7282 37236
rect 7248 35850 7282 36142
rect 8472 36952 8506 37244
rect 8472 35858 8506 36150
rect 7248 34756 7282 35048
rect 7840 34514 7934 35710
rect 8472 34764 8506 35056
rect 7248 33662 7282 33954
rect 7248 32568 7282 32860
rect 8472 33670 8506 33962
rect 8472 32576 8506 32868
rect 9530 36952 9564 37244
rect 9530 35858 9564 36150
rect 9530 34764 9564 35056
rect 9530 33670 9564 33962
rect 1958 31110 1992 31402
rect 1958 30016 1992 30308
rect 1326 28672 1420 29868
rect 1958 28922 1992 29214
rect 1958 27828 1992 28120
rect 1958 26734 1992 27026
rect 3016 31110 3050 31402
rect 3016 30016 3050 30308
rect 3016 28922 3050 29214
rect 3016 27828 3050 28120
rect 3016 26734 3050 27026
rect 4074 31110 4108 31402
rect 4074 30016 4108 30308
rect 4074 28922 4108 29214
rect 4074 27828 4108 28120
rect 4074 26734 4108 27026
rect 5132 31110 5166 31402
rect 5132 30016 5166 30308
rect 5132 28922 5166 29214
rect 5132 27828 5166 28120
rect 5132 26734 5166 27026
rect 6190 31110 6224 31402
rect 9530 32576 9564 32868
rect 10588 36952 10622 37244
rect 10588 35858 10622 36150
rect 10588 34764 10622 35056
rect 10588 33670 10622 33962
rect 10588 32576 10622 32868
rect 11646 36952 11680 37244
rect 16036 38400 16070 38692
rect 17094 42776 17128 43068
rect 17094 41682 17128 41974
rect 17094 40588 17128 40880
rect 17094 39494 17128 39786
rect 17094 38400 17128 38692
rect 18152 42776 18186 43068
rect 18152 41682 18186 41974
rect 18152 40588 18186 40880
rect 18152 39494 18186 39786
rect 18152 38400 18186 38692
rect 19210 42776 19244 43068
rect 19210 41682 19244 41974
rect 19210 40588 19244 40880
rect 19210 39494 19244 39786
rect 19210 38400 19244 38692
rect 20268 42776 20302 43068
rect 20268 41682 20302 41974
rect 21468 42760 21502 43052
rect 22526 42760 22560 43052
rect 21468 41666 21502 41958
rect 22526 41666 22560 41958
rect 20268 40588 20302 40880
rect 20836 40322 20930 41518
rect 21468 40572 21502 40864
rect 22526 40572 22560 40864
rect 20268 39494 20302 39786
rect 21468 39478 21502 39770
rect 22526 39478 22560 39770
rect 20268 38400 20302 38692
rect 21468 38384 21502 38676
rect 11646 35858 11680 36150
rect 11646 34764 11680 35056
rect 11646 33670 11680 33962
rect 11646 32576 11680 32868
rect 12704 36952 12738 37244
rect 12704 35858 12738 36150
rect 12704 34764 12738 35056
rect 12704 33670 12738 33962
rect 12704 32576 12738 32868
rect 13762 36952 13796 37244
rect 13762 35858 13796 36150
rect 14978 36960 15012 37252
rect 14978 35866 15012 36158
rect 13762 34764 13796 35056
rect 14346 34522 14440 35718
rect 14978 34772 15012 35064
rect 13762 33670 13796 33962
rect 13762 32576 13796 32868
rect 14978 33678 15012 33970
rect 14978 32584 15012 32876
rect 16036 36960 16070 37252
rect 16036 35866 16070 36158
rect 16036 34772 16070 35064
rect 16036 33678 16070 33970
rect 6190 30016 6224 30308
rect 6190 28922 6224 29214
rect 6190 27828 6224 28120
rect 6190 26734 6224 27026
rect 7248 31110 7282 31402
rect 7248 30016 7282 30308
rect 8472 31118 8506 31410
rect 8472 30024 8506 30316
rect 7248 28922 7282 29214
rect 7840 28680 7934 29876
rect 8472 28930 8506 29222
rect 7248 27828 7282 28120
rect 7248 26734 7282 27026
rect 8472 27836 8506 28128
rect 8472 26742 8506 27034
rect 9530 31118 9564 31410
rect 9530 30024 9564 30316
rect 9530 28930 9564 29222
rect 9530 27836 9564 28128
rect 1958 25274 1992 25566
rect 1958 24180 1992 24472
rect 1326 22836 1420 24032
rect 1958 23086 1992 23378
rect 1958 21992 1992 22284
rect 1958 20898 1992 21190
rect 3016 25274 3050 25566
rect 3016 24180 3050 24472
rect 3016 23086 3050 23378
rect 3016 21992 3050 22284
rect 3016 20898 3050 21190
rect 4074 25274 4108 25566
rect 4074 24180 4108 24472
rect 4074 23086 4108 23378
rect 4074 21992 4108 22284
rect 4074 20898 4108 21190
rect 5132 25274 5166 25566
rect 5132 24180 5166 24472
rect 5132 23086 5166 23378
rect 5132 21992 5166 22284
rect 5132 20898 5166 21190
rect 6190 25274 6224 25566
rect 9530 26742 9564 27034
rect 10588 31118 10622 31410
rect 10588 30024 10622 30316
rect 10588 28930 10622 29222
rect 10588 27836 10622 28128
rect 10588 26742 10622 27034
rect 11646 31118 11680 31410
rect 16036 32584 16070 32876
rect 17094 36960 17128 37252
rect 17094 35866 17128 36158
rect 17094 34772 17128 35064
rect 17094 33678 17128 33970
rect 17094 32584 17128 32876
rect 18152 36960 18186 37252
rect 18152 35866 18186 36158
rect 18152 34772 18186 35064
rect 18152 33678 18186 33970
rect 18152 32584 18186 32876
rect 19210 36960 19244 37252
rect 22526 38384 22560 38676
rect 23584 42760 23618 43052
rect 23584 41666 23618 41958
rect 23584 40572 23618 40864
rect 23584 39478 23618 39770
rect 23584 38384 23618 38676
rect 24642 42760 24676 43052
rect 24642 41666 24676 41958
rect 24642 40572 24676 40864
rect 24642 39478 24676 39770
rect 24642 38384 24676 38676
rect 25700 42760 25734 43052
rect 25700 41666 25734 41958
rect 25700 40572 25734 40864
rect 25700 39478 25734 39770
rect 25700 38384 25734 38676
rect 26758 42760 26792 43052
rect 26758 41666 26792 41958
rect 27990 42776 28024 43068
rect 29048 42776 29082 43068
rect 27990 41682 28024 41974
rect 29048 41682 29082 41974
rect 26758 40572 26792 40864
rect 27358 40338 27452 41534
rect 27990 40588 28024 40880
rect 29048 40588 29082 40880
rect 26758 39478 26792 39770
rect 27990 39494 28024 39786
rect 29048 39494 29082 39786
rect 26758 38384 26792 38676
rect 27990 38400 28024 38692
rect 19210 35866 19244 36158
rect 19210 34772 19244 35064
rect 19210 33678 19244 33970
rect 19210 32584 19244 32876
rect 20268 36960 20302 37252
rect 20268 35866 20302 36158
rect 21468 36944 21502 37236
rect 22526 36944 22560 37236
rect 21468 35850 21502 36142
rect 22526 35850 22560 36142
rect 20268 34772 20302 35064
rect 20836 34506 20930 35702
rect 21468 34756 21502 35048
rect 22526 34756 22560 35048
rect 20268 33678 20302 33970
rect 21468 33662 21502 33954
rect 22526 33662 22560 33954
rect 20268 32584 20302 32876
rect 21468 32568 21502 32860
rect 11646 30024 11680 30316
rect 11646 28930 11680 29222
rect 11646 27836 11680 28128
rect 11646 26742 11680 27034
rect 12704 31118 12738 31410
rect 12704 30024 12738 30316
rect 12704 28930 12738 29222
rect 12704 27836 12738 28128
rect 12704 26742 12738 27034
rect 13762 31118 13796 31410
rect 13762 30024 13796 30316
rect 14978 31126 15012 31418
rect 14978 30032 15012 30324
rect 13762 28930 13796 29222
rect 14346 28688 14440 29884
rect 14978 28938 15012 29230
rect 13762 27836 13796 28128
rect 13762 26742 13796 27034
rect 14978 27844 15012 28136
rect 14978 26750 15012 27042
rect 16036 31126 16070 31418
rect 16036 30032 16070 30324
rect 16036 28938 16070 29230
rect 16036 27844 16070 28136
rect 6190 24180 6224 24472
rect 6190 23086 6224 23378
rect 6190 21992 6224 22284
rect 6190 20898 6224 21190
rect 7248 25274 7282 25566
rect 7248 24180 7282 24472
rect 8472 25282 8506 25574
rect 8472 24188 8506 24480
rect 7248 23086 7282 23378
rect 7840 22844 7934 24040
rect 8472 23094 8506 23386
rect 7248 21992 7282 22284
rect 7248 20898 7282 21190
rect 8472 22000 8506 22292
rect 8472 20906 8506 21198
rect 9530 25282 9564 25574
rect 9530 24188 9564 24480
rect 9530 23094 9564 23386
rect 9530 22000 9564 22292
rect 1958 19410 1992 19702
rect 1958 18316 1992 18608
rect 1326 16972 1420 18168
rect 1958 17222 1992 17514
rect 1958 16128 1992 16420
rect 1958 15034 1992 15326
rect 3016 19410 3050 19702
rect 3016 18316 3050 18608
rect 3016 17222 3050 17514
rect 3016 16128 3050 16420
rect 3016 15034 3050 15326
rect 4074 19410 4108 19702
rect 4074 18316 4108 18608
rect 4074 17222 4108 17514
rect 4074 16128 4108 16420
rect 4074 15034 4108 15326
rect 5132 19410 5166 19702
rect 5132 18316 5166 18608
rect 5132 17222 5166 17514
rect 5132 16128 5166 16420
rect 5132 15034 5166 15326
rect 6190 19410 6224 19702
rect 9530 20906 9564 21198
rect 10588 25282 10622 25574
rect 10588 24188 10622 24480
rect 10588 23094 10622 23386
rect 10588 22000 10622 22292
rect 10588 20906 10622 21198
rect 11646 25282 11680 25574
rect 16036 26750 16070 27042
rect 17094 31126 17128 31418
rect 17094 30032 17128 30324
rect 17094 28938 17128 29230
rect 17094 27844 17128 28136
rect 17094 26750 17128 27042
rect 18152 31126 18186 31418
rect 18152 30032 18186 30324
rect 18152 28938 18186 29230
rect 18152 27844 18186 28136
rect 18152 26750 18186 27042
rect 19210 31126 19244 31418
rect 22526 32568 22560 32860
rect 23584 36944 23618 37236
rect 23584 35850 23618 36142
rect 23584 34756 23618 35048
rect 23584 33662 23618 33954
rect 23584 32568 23618 32860
rect 24642 36944 24676 37236
rect 24642 35850 24676 36142
rect 24642 34756 24676 35048
rect 24642 33662 24676 33954
rect 24642 32568 24676 32860
rect 25700 36944 25734 37236
rect 29048 38400 29082 38692
rect 30106 42776 30140 43068
rect 30106 41682 30140 41974
rect 30106 40588 30140 40880
rect 30106 39494 30140 39786
rect 30106 38400 30140 38692
rect 31164 42776 31198 43068
rect 31164 41682 31198 41974
rect 31164 40588 31198 40880
rect 31164 39494 31198 39786
rect 31164 38400 31198 38692
rect 32222 42776 32256 43068
rect 32222 41682 32256 41974
rect 32222 40588 32256 40880
rect 32222 39494 32256 39786
rect 32222 38400 32256 38692
rect 33280 42776 33314 43068
rect 33280 41682 33314 41974
rect 34500 42782 34534 43074
rect 35558 42782 35592 43074
rect 34500 41688 34534 41980
rect 35558 41688 35592 41980
rect 33280 40588 33314 40880
rect 33868 40344 33962 41540
rect 34500 40594 34534 40886
rect 35558 40594 35592 40886
rect 33280 39494 33314 39786
rect 34500 39500 34534 39792
rect 35558 39500 35592 39792
rect 33280 38400 33314 38692
rect 34500 38406 34534 38698
rect 25700 35850 25734 36142
rect 25700 34756 25734 35048
rect 25700 33662 25734 33954
rect 25700 32568 25734 32860
rect 26758 36944 26792 37236
rect 26758 35850 26792 36142
rect 27990 36960 28024 37252
rect 29048 36960 29082 37252
rect 27990 35866 28024 36158
rect 29048 35866 29082 36158
rect 26758 34756 26792 35048
rect 27358 34522 27452 35718
rect 27990 34772 28024 35064
rect 29048 34772 29082 35064
rect 26758 33662 26792 33954
rect 27990 33678 28024 33970
rect 29048 33678 29082 33970
rect 26758 32568 26792 32860
rect 27990 32584 28024 32876
rect 19210 30032 19244 30324
rect 19210 28938 19244 29230
rect 19210 27844 19244 28136
rect 19210 26750 19244 27042
rect 20268 31126 20302 31418
rect 20268 30032 20302 30324
rect 21468 31110 21502 31402
rect 22526 31110 22560 31402
rect 21468 30016 21502 30308
rect 22526 30016 22560 30308
rect 20268 28938 20302 29230
rect 20836 28672 20930 29868
rect 21468 28922 21502 29214
rect 22526 28922 22560 29214
rect 20268 27844 20302 28136
rect 21468 27828 21502 28120
rect 22526 27828 22560 28120
rect 20268 26750 20302 27042
rect 21468 26734 21502 27026
rect 11646 24188 11680 24480
rect 11646 23094 11680 23386
rect 11646 22000 11680 22292
rect 11646 20906 11680 21198
rect 12704 25282 12738 25574
rect 12704 24188 12738 24480
rect 12704 23094 12738 23386
rect 12704 22000 12738 22292
rect 12704 20906 12738 21198
rect 13762 25282 13796 25574
rect 13762 24188 13796 24480
rect 14978 25290 15012 25582
rect 14978 24196 15012 24488
rect 13762 23094 13796 23386
rect 14346 22852 14440 24048
rect 14978 23102 15012 23394
rect 13762 22000 13796 22292
rect 13762 20906 13796 21198
rect 14978 22008 15012 22300
rect 14978 20914 15012 21206
rect 16036 25290 16070 25582
rect 16036 24196 16070 24488
rect 16036 23102 16070 23394
rect 16036 22008 16070 22300
rect 6190 18316 6224 18608
rect 6190 17222 6224 17514
rect 6190 16128 6224 16420
rect 6190 15034 6224 15326
rect 7248 19410 7282 19702
rect 7248 18316 7282 18608
rect 8472 19418 8506 19710
rect 8472 18324 8506 18616
rect 7248 17222 7282 17514
rect 7840 16980 7934 18176
rect 8472 17230 8506 17522
rect 7248 16128 7282 16420
rect 7248 15034 7282 15326
rect 8472 16136 8506 16428
rect 8472 15042 8506 15334
rect 9530 19418 9564 19710
rect 9530 18324 9564 18616
rect 9530 17230 9564 17522
rect 9530 16136 9564 16428
rect 1968 13554 2002 13846
rect 1968 12460 2002 12752
rect 1336 11116 1430 12312
rect 1968 11366 2002 11658
rect 1968 10272 2002 10564
rect 1968 9178 2002 9470
rect 3026 13554 3060 13846
rect 3026 12460 3060 12752
rect 3026 11366 3060 11658
rect 3026 10272 3060 10564
rect 3026 9178 3060 9470
rect 4084 13554 4118 13846
rect 4084 12460 4118 12752
rect 4084 11366 4118 11658
rect 4084 10272 4118 10564
rect 4084 9178 4118 9470
rect 5142 13554 5176 13846
rect 5142 12460 5176 12752
rect 5142 11366 5176 11658
rect 5142 10272 5176 10564
rect 5142 9178 5176 9470
rect 6200 13554 6234 13846
rect 9530 15042 9564 15334
rect 10588 19418 10622 19710
rect 10588 18324 10622 18616
rect 10588 17230 10622 17522
rect 10588 16136 10622 16428
rect 10588 15042 10622 15334
rect 11646 19418 11680 19710
rect 16036 20914 16070 21206
rect 17094 25290 17128 25582
rect 17094 24196 17128 24488
rect 17094 23102 17128 23394
rect 17094 22008 17128 22300
rect 17094 20914 17128 21206
rect 18152 25290 18186 25582
rect 18152 24196 18186 24488
rect 18152 23102 18186 23394
rect 18152 22008 18186 22300
rect 18152 20914 18186 21206
rect 19210 25290 19244 25582
rect 22526 26734 22560 27026
rect 23584 31110 23618 31402
rect 23584 30016 23618 30308
rect 23584 28922 23618 29214
rect 23584 27828 23618 28120
rect 23584 26734 23618 27026
rect 24642 31110 24676 31402
rect 24642 30016 24676 30308
rect 24642 28922 24676 29214
rect 24642 27828 24676 28120
rect 24642 26734 24676 27026
rect 25700 31110 25734 31402
rect 29048 32584 29082 32876
rect 30106 36960 30140 37252
rect 30106 35866 30140 36158
rect 30106 34772 30140 35064
rect 30106 33678 30140 33970
rect 30106 32584 30140 32876
rect 31164 36960 31198 37252
rect 31164 35866 31198 36158
rect 31164 34772 31198 35064
rect 31164 33678 31198 33970
rect 31164 32584 31198 32876
rect 32222 36960 32256 37252
rect 35558 38406 35592 38698
rect 36616 42782 36650 43074
rect 36616 41688 36650 41980
rect 36616 40594 36650 40886
rect 36616 39500 36650 39792
rect 36616 38406 36650 38698
rect 37674 42782 37708 43074
rect 49622 43720 49866 43888
rect 63846 43492 64132 43614
rect 68426 43844 68848 43922
rect 37674 41688 37708 41980
rect 37674 40594 37708 40886
rect 37674 39500 37708 39792
rect 37674 38406 37708 38698
rect 38732 42782 38766 43074
rect 39790 42782 39824 43074
rect 40990 42782 41024 43074
rect 42048 42782 42082 43074
rect 38732 41688 38766 41980
rect 38732 40594 38766 40886
rect 38732 39500 38766 39792
rect 38732 38406 38766 38698
rect 39790 41688 39824 41980
rect 40990 41688 41024 41980
rect 42048 41688 42082 41980
rect 39790 40594 39824 40886
rect 40358 40344 40452 41540
rect 40990 40594 41024 40886
rect 42048 40594 42082 40886
rect 39790 39500 39824 39792
rect 39790 38406 39824 38698
rect 40990 39500 41024 39792
rect 42048 39500 42082 39792
rect 40990 38406 41024 38698
rect 32222 35866 32256 36158
rect 32222 34772 32256 35064
rect 32222 33678 32256 33970
rect 32222 32584 32256 32876
rect 33280 36960 33314 37252
rect 33280 35866 33314 36158
rect 34500 36966 34534 37258
rect 35558 36966 35592 37258
rect 34500 35872 34534 36164
rect 35558 35872 35592 36164
rect 33280 34772 33314 35064
rect 33868 34528 33962 35724
rect 34500 34778 34534 35070
rect 35558 34778 35592 35070
rect 33280 33678 33314 33970
rect 33280 32584 33314 32876
rect 34500 33684 34534 33976
rect 35558 33684 35592 33976
rect 34500 32590 34534 32882
rect 25700 30016 25734 30308
rect 25700 28922 25734 29214
rect 25700 27828 25734 28120
rect 25700 26734 25734 27026
rect 26758 31110 26792 31402
rect 26758 30016 26792 30308
rect 27990 31126 28024 31418
rect 29048 31126 29082 31418
rect 27990 30032 28024 30324
rect 29048 30032 29082 30324
rect 26758 28922 26792 29214
rect 27358 28688 27452 29884
rect 27990 28938 28024 29230
rect 29048 28938 29082 29230
rect 26758 27828 26792 28120
rect 27990 27844 28024 28136
rect 29048 27844 29082 28136
rect 26758 26734 26792 27026
rect 27990 26750 28024 27042
rect 19210 24196 19244 24488
rect 19210 23102 19244 23394
rect 19210 22008 19244 22300
rect 19210 20914 19244 21206
rect 20268 25290 20302 25582
rect 20268 24196 20302 24488
rect 21468 25274 21502 25566
rect 22526 25274 22560 25566
rect 21468 24180 21502 24472
rect 22526 24180 22560 24472
rect 20268 23102 20302 23394
rect 20836 22836 20930 24032
rect 21468 23086 21502 23378
rect 22526 23086 22560 23378
rect 20268 22008 20302 22300
rect 20268 20914 20302 21206
rect 21468 21992 21502 22284
rect 22526 21992 22560 22284
rect 21468 20898 21502 21190
rect 11646 18324 11680 18616
rect 11646 17230 11680 17522
rect 11646 16136 11680 16428
rect 11646 15042 11680 15334
rect 12704 19418 12738 19710
rect 12704 18324 12738 18616
rect 12704 17230 12738 17522
rect 12704 16136 12738 16428
rect 12704 15042 12738 15334
rect 13762 19418 13796 19710
rect 13762 18324 13796 18616
rect 14978 19426 15012 19718
rect 14978 18332 15012 18624
rect 13762 17230 13796 17522
rect 14346 16988 14440 18184
rect 14978 17238 15012 17530
rect 13762 16136 13796 16428
rect 13762 15042 13796 15334
rect 14978 16144 15012 16436
rect 14978 15050 15012 15342
rect 16036 19426 16070 19718
rect 16036 18332 16070 18624
rect 16036 17238 16070 17530
rect 16036 16144 16070 16436
rect 6200 12460 6234 12752
rect 6200 11366 6234 11658
rect 6200 10272 6234 10564
rect 6200 9178 6234 9470
rect 7258 13554 7292 13846
rect 7258 12460 7292 12752
rect 8482 13562 8516 13854
rect 8482 12468 8516 12760
rect 7258 11366 7292 11658
rect 7850 11124 7944 12320
rect 8482 11374 8516 11666
rect 7258 10272 7292 10564
rect 7258 9178 7292 9470
rect 8482 10280 8516 10572
rect 8482 9186 8516 9478
rect 9540 13562 9574 13854
rect 9540 12468 9574 12760
rect 9540 11374 9574 11666
rect 9540 10280 9574 10572
rect 1986 7646 2020 7938
rect 3044 7646 3078 7938
rect 1986 6552 2020 6844
rect 3044 6552 3078 6844
rect 1354 5208 1448 6404
rect 1986 5458 2020 5750
rect 3044 5458 3078 5750
rect 1986 4364 2020 4656
rect 3044 4364 3078 4656
rect 1986 3270 2020 3562
rect 3044 3270 3078 3562
rect 4102 7646 4136 7938
rect 4102 6552 4136 6844
rect 4102 5458 4136 5750
rect 4102 4364 4136 4656
rect 4102 3270 4136 3562
rect 5160 7646 5194 7938
rect 5160 6552 5194 6844
rect 5160 5458 5194 5750
rect 5160 4364 5194 4656
rect 5160 3270 5194 3562
rect 6218 7646 6252 7938
rect 9540 9186 9574 9478
rect 10598 13562 10632 13854
rect 10598 12468 10632 12760
rect 10598 11374 10632 11666
rect 10598 10280 10632 10572
rect 10598 9186 10632 9478
rect 11656 13562 11690 13854
rect 11656 12468 11690 12760
rect 11656 11374 11690 11666
rect 11656 10280 11690 10572
rect 11656 9186 11690 9478
rect 12714 13562 12748 13854
rect 16036 15050 16070 15342
rect 17094 19426 17128 19718
rect 17094 18332 17128 18624
rect 17094 17238 17128 17530
rect 17094 16144 17128 16436
rect 17094 15050 17128 15342
rect 18152 19426 18186 19718
rect 18152 18332 18186 18624
rect 18152 17238 18186 17530
rect 18152 16144 18186 16436
rect 18152 15050 18186 15342
rect 19210 19426 19244 19718
rect 22526 20898 22560 21190
rect 23584 25274 23618 25566
rect 23584 24180 23618 24472
rect 23584 23086 23618 23378
rect 23584 21992 23618 22284
rect 23584 20898 23618 21190
rect 24642 25274 24676 25566
rect 24642 24180 24676 24472
rect 24642 23086 24676 23378
rect 24642 21992 24676 22284
rect 24642 20898 24676 21190
rect 25700 25274 25734 25566
rect 29048 26750 29082 27042
rect 30106 31126 30140 31418
rect 30106 30032 30140 30324
rect 30106 28938 30140 29230
rect 30106 27844 30140 28136
rect 30106 26750 30140 27042
rect 31164 31126 31198 31418
rect 31164 30032 31198 30324
rect 31164 28938 31198 29230
rect 31164 27844 31198 28136
rect 31164 26750 31198 27042
rect 32222 31126 32256 31418
rect 35558 32590 35592 32882
rect 36616 36966 36650 37258
rect 36616 35872 36650 36164
rect 36616 34778 36650 35070
rect 36616 33684 36650 33976
rect 36616 32590 36650 32882
rect 37674 36966 37708 37258
rect 37674 35872 37708 36164
rect 37674 34778 37708 35070
rect 37674 33684 37708 33976
rect 37674 32590 37708 32882
rect 38732 36966 38766 37258
rect 42048 38406 42082 38698
rect 43106 42782 43140 43074
rect 43106 41688 43140 41980
rect 43106 40594 43140 40886
rect 43106 39500 43140 39792
rect 43106 38406 43140 38698
rect 44164 42782 44198 43074
rect 44164 41688 44198 41980
rect 44164 40594 44198 40886
rect 44164 39500 44198 39792
rect 44164 38406 44198 38698
rect 45222 42782 45256 43074
rect 46280 42782 46314 43074
rect 47578 42804 47612 43096
rect 48636 42804 48670 43096
rect 45222 41688 45256 41980
rect 45222 40594 45256 40886
rect 45222 39500 45256 39792
rect 45222 38406 45256 38698
rect 46280 41688 46314 41980
rect 47578 41710 47612 42002
rect 48636 41710 48670 42002
rect 46280 40594 46314 40886
rect 46946 40366 47040 41562
rect 47578 40616 47612 40908
rect 48636 40616 48670 40908
rect 46280 39500 46314 39792
rect 46280 38406 46314 38698
rect 47578 39522 47612 39814
rect 48636 39522 48670 39814
rect 47578 38428 47612 38720
rect 38732 35872 38766 36164
rect 38732 34778 38766 35070
rect 38732 33684 38766 33976
rect 38732 32590 38766 32882
rect 39790 36966 39824 37258
rect 39790 35872 39824 36164
rect 40990 36966 41024 37258
rect 42048 36966 42082 37258
rect 40990 35872 41024 36164
rect 42048 35872 42082 36164
rect 39790 34778 39824 35070
rect 40358 34528 40452 35724
rect 40990 34778 41024 35070
rect 42048 34778 42082 35070
rect 39790 33684 39824 33976
rect 39790 32590 39824 32882
rect 40990 33684 41024 33976
rect 42048 33684 42082 33976
rect 40990 32590 41024 32882
rect 32222 30032 32256 30324
rect 32222 28938 32256 29230
rect 32222 27844 32256 28136
rect 32222 26750 32256 27042
rect 33280 31126 33314 31418
rect 33280 30032 33314 30324
rect 34500 31132 34534 31424
rect 35558 31132 35592 31424
rect 34500 30038 34534 30330
rect 35558 30038 35592 30330
rect 33280 28938 33314 29230
rect 33868 28694 33962 29890
rect 34500 28944 34534 29236
rect 35558 28944 35592 29236
rect 33280 27844 33314 28136
rect 33280 26750 33314 27042
rect 34500 27850 34534 28142
rect 35558 27850 35592 28142
rect 34500 26756 34534 27048
rect 25700 24180 25734 24472
rect 25700 23086 25734 23378
rect 25700 21992 25734 22284
rect 25700 20898 25734 21190
rect 26758 25274 26792 25566
rect 26758 24180 26792 24472
rect 27990 25290 28024 25582
rect 29048 25290 29082 25582
rect 27990 24196 28024 24488
rect 29048 24196 29082 24488
rect 26758 23086 26792 23378
rect 27358 22852 27452 24048
rect 27990 23102 28024 23394
rect 29048 23102 29082 23394
rect 26758 21992 26792 22284
rect 27990 22008 28024 22300
rect 29048 22008 29082 22300
rect 26758 20898 26792 21190
rect 27990 20914 28024 21206
rect 19210 18332 19244 18624
rect 19210 17238 19244 17530
rect 19210 16144 19244 16436
rect 19210 15050 19244 15342
rect 20268 19426 20302 19718
rect 20268 18332 20302 18624
rect 21468 19410 21502 19702
rect 22526 19410 22560 19702
rect 21468 18316 21502 18608
rect 22526 18316 22560 18608
rect 20268 17238 20302 17530
rect 20836 16972 20930 18168
rect 21468 17222 21502 17514
rect 22526 17222 22560 17514
rect 20268 16144 20302 16436
rect 20268 15050 20302 15342
rect 21468 16128 21502 16420
rect 22526 16128 22560 16420
rect 21468 15034 21502 15326
rect 12714 12468 12748 12760
rect 12714 11374 12748 11666
rect 12714 10280 12748 10572
rect 12714 9186 12748 9478
rect 13772 13562 13806 13854
rect 13772 12468 13806 12760
rect 14988 13570 15022 13862
rect 14988 12476 15022 12768
rect 13772 11374 13806 11666
rect 14356 11132 14450 12328
rect 14988 11382 15022 11674
rect 13772 10280 13806 10572
rect 13772 9186 13806 9478
rect 14988 10288 15022 10580
rect 14988 9194 15022 9486
rect 16046 13570 16080 13862
rect 16046 12476 16080 12768
rect 16046 11382 16080 11674
rect 16046 10288 16080 10580
rect 6218 6552 6252 6844
rect 6218 5458 6252 5750
rect 6218 4364 6252 4656
rect 6218 3270 6252 3562
rect 7276 7646 7310 7938
rect 7276 6552 7310 6844
rect 8500 7654 8534 7946
rect 9558 7654 9592 7946
rect 8500 6560 8534 6852
rect 9558 6560 9592 6852
rect 7276 5458 7310 5750
rect 7868 5216 7962 6412
rect 8500 5466 8534 5758
rect 9558 5466 9592 5758
rect 7276 4364 7310 4656
rect 7276 3270 7310 3562
rect 8500 4372 8534 4664
rect 9558 4372 9592 4664
rect 8500 3278 8534 3570
rect 9558 3278 9592 3570
rect 10616 7654 10650 7946
rect 10616 6560 10650 6852
rect 10616 5466 10650 5758
rect 10616 4372 10650 4664
rect 10616 3278 10650 3570
rect 11674 7654 11708 7946
rect 11674 6560 11708 6852
rect 11674 5466 11708 5758
rect 11674 4372 11708 4664
rect 11674 3278 11708 3570
rect 12732 7654 12766 7946
rect 16046 9194 16080 9486
rect 17104 13570 17138 13862
rect 17104 12476 17138 12768
rect 17104 11382 17138 11674
rect 17104 10288 17138 10580
rect 17104 9194 17138 9486
rect 18162 13570 18196 13862
rect 18162 12476 18196 12768
rect 18162 11382 18196 11674
rect 18162 10288 18196 10580
rect 18162 9194 18196 9486
rect 19220 13570 19254 13862
rect 22526 15034 22560 15326
rect 23584 19410 23618 19702
rect 23584 18316 23618 18608
rect 23584 17222 23618 17514
rect 23584 16128 23618 16420
rect 23584 15034 23618 15326
rect 24642 19410 24676 19702
rect 24642 18316 24676 18608
rect 24642 17222 24676 17514
rect 24642 16128 24676 16420
rect 24642 15034 24676 15326
rect 25700 19410 25734 19702
rect 29048 20914 29082 21206
rect 30106 25290 30140 25582
rect 30106 24196 30140 24488
rect 30106 23102 30140 23394
rect 30106 22008 30140 22300
rect 30106 20914 30140 21206
rect 31164 25290 31198 25582
rect 31164 24196 31198 24488
rect 31164 23102 31198 23394
rect 31164 22008 31198 22300
rect 31164 20914 31198 21206
rect 32222 25290 32256 25582
rect 35558 26756 35592 27048
rect 36616 31132 36650 31424
rect 36616 30038 36650 30330
rect 36616 28944 36650 29236
rect 36616 27850 36650 28142
rect 36616 26756 36650 27048
rect 37674 31132 37708 31424
rect 37674 30038 37708 30330
rect 37674 28944 37708 29236
rect 37674 27850 37708 28142
rect 37674 26756 37708 27048
rect 38732 31132 38766 31424
rect 42048 32590 42082 32882
rect 43106 36966 43140 37258
rect 43106 35872 43140 36164
rect 43106 34778 43140 35070
rect 43106 33684 43140 33976
rect 43106 32590 43140 32882
rect 44164 36966 44198 37258
rect 44164 35872 44198 36164
rect 44164 34778 44198 35070
rect 44164 33684 44198 33976
rect 44164 32590 44198 32882
rect 45222 36966 45256 37258
rect 48636 38428 48670 38720
rect 49694 42804 49728 43096
rect 49694 41710 49728 42002
rect 49694 40616 49728 40908
rect 49694 39522 49728 39814
rect 49694 38428 49728 38720
rect 50752 42804 50786 43096
rect 50752 41710 50786 42002
rect 50752 40616 50786 40908
rect 50752 39522 50786 39814
rect 50752 38428 50786 38720
rect 51810 42804 51844 43096
rect 52868 42804 52902 43096
rect 54092 42818 54126 43110
rect 55150 42818 55184 43110
rect 51810 41710 51844 42002
rect 51810 40616 51844 40908
rect 51810 39522 51844 39814
rect 51810 38428 51844 38720
rect 52868 41710 52902 42002
rect 54092 41724 54126 42016
rect 55150 41724 55184 42016
rect 52868 40616 52902 40908
rect 53460 40380 53554 41576
rect 54092 40630 54126 40922
rect 55150 40630 55184 40922
rect 52868 39522 52902 39814
rect 52868 38428 52902 38720
rect 54092 39536 54126 39828
rect 55150 39536 55184 39828
rect 54092 38442 54126 38734
rect 45222 35872 45256 36164
rect 45222 34778 45256 35070
rect 45222 33684 45256 33976
rect 45222 32590 45256 32882
rect 46280 36966 46314 37258
rect 46280 35872 46314 36164
rect 47578 36988 47612 37280
rect 48636 36988 48670 37280
rect 47578 35894 47612 36186
rect 48636 35894 48670 36186
rect 46280 34778 46314 35070
rect 46946 34550 47040 35746
rect 47578 34800 47612 35092
rect 48636 34800 48670 35092
rect 46280 33684 46314 33976
rect 46280 32590 46314 32882
rect 47578 33706 47612 33998
rect 48636 33706 48670 33998
rect 47578 32612 47612 32904
rect 38732 30038 38766 30330
rect 38732 28944 38766 29236
rect 38732 27850 38766 28142
rect 38732 26756 38766 27048
rect 39790 31132 39824 31424
rect 39790 30038 39824 30330
rect 40990 31132 41024 31424
rect 42048 31132 42082 31424
rect 40990 30038 41024 30330
rect 42048 30038 42082 30330
rect 39790 28944 39824 29236
rect 40358 28694 40452 29890
rect 40990 28944 41024 29236
rect 42048 28944 42082 29236
rect 39790 27850 39824 28142
rect 39790 26756 39824 27048
rect 40990 27850 41024 28142
rect 42048 27850 42082 28142
rect 40990 26756 41024 27048
rect 32222 24196 32256 24488
rect 32222 23102 32256 23394
rect 32222 22008 32256 22300
rect 32222 20914 32256 21206
rect 33280 25290 33314 25582
rect 33280 24196 33314 24488
rect 34500 25296 34534 25588
rect 35558 25296 35592 25588
rect 34500 24202 34534 24494
rect 35558 24202 35592 24494
rect 33280 23102 33314 23394
rect 33868 22858 33962 24054
rect 34500 23108 34534 23400
rect 35558 23108 35592 23400
rect 33280 22008 33314 22300
rect 33280 20914 33314 21206
rect 34500 22014 34534 22306
rect 35558 22014 35592 22306
rect 34500 20920 34534 21212
rect 25700 18316 25734 18608
rect 25700 17222 25734 17514
rect 25700 16128 25734 16420
rect 25700 15034 25734 15326
rect 26758 19410 26792 19702
rect 26758 18316 26792 18608
rect 27990 19426 28024 19718
rect 29048 19426 29082 19718
rect 27990 18332 28024 18624
rect 29048 18332 29082 18624
rect 26758 17222 26792 17514
rect 27358 16988 27452 18184
rect 27990 17238 28024 17530
rect 29048 17238 29082 17530
rect 26758 16128 26792 16420
rect 27990 16144 28024 16436
rect 29048 16144 29082 16436
rect 26758 15034 26792 15326
rect 27990 15050 28024 15342
rect 19220 12476 19254 12768
rect 19220 11382 19254 11674
rect 19220 10288 19254 10580
rect 19220 9194 19254 9486
rect 20278 13570 20312 13862
rect 20278 12476 20312 12768
rect 21478 13554 21512 13846
rect 22536 13554 22570 13846
rect 21478 12460 21512 12752
rect 22536 12460 22570 12752
rect 20278 11382 20312 11674
rect 20846 11116 20940 12312
rect 21478 11366 21512 11658
rect 22536 11366 22570 11658
rect 20278 10288 20312 10580
rect 20278 9194 20312 9486
rect 21478 10272 21512 10564
rect 22536 10272 22570 10564
rect 21478 9178 21512 9470
rect 12732 6560 12766 6852
rect 12732 5466 12766 5758
rect 12732 4372 12766 4664
rect 12732 3278 12766 3570
rect 13790 7654 13824 7946
rect 13790 6560 13824 6852
rect 15006 7662 15040 7954
rect 16064 7662 16098 7954
rect 15006 6568 15040 6860
rect 16064 6568 16098 6860
rect 13790 5466 13824 5758
rect 14374 5224 14468 6420
rect 15006 5474 15040 5766
rect 16064 5474 16098 5766
rect 13790 4372 13824 4664
rect 13790 3278 13824 3570
rect 15006 4380 15040 4672
rect 16064 4380 16098 4672
rect 15006 3286 15040 3578
rect 16064 3286 16098 3578
rect 17122 7662 17156 7954
rect 17122 6568 17156 6860
rect 17122 5474 17156 5766
rect 17122 4380 17156 4672
rect 17122 3286 17156 3578
rect 18180 7662 18214 7954
rect 18180 6568 18214 6860
rect 18180 5474 18214 5766
rect 18180 4380 18214 4672
rect 18180 3286 18214 3578
rect 19238 7662 19272 7954
rect 22536 9178 22570 9470
rect 23594 13554 23628 13846
rect 23594 12460 23628 12752
rect 23594 11366 23628 11658
rect 23594 10272 23628 10564
rect 23594 9178 23628 9470
rect 24652 13554 24686 13846
rect 24652 12460 24686 12752
rect 24652 11366 24686 11658
rect 24652 10272 24686 10564
rect 24652 9178 24686 9470
rect 25710 13554 25744 13846
rect 29048 15050 29082 15342
rect 30106 19426 30140 19718
rect 30106 18332 30140 18624
rect 30106 17238 30140 17530
rect 30106 16144 30140 16436
rect 30106 15050 30140 15342
rect 31164 19426 31198 19718
rect 31164 18332 31198 18624
rect 31164 17238 31198 17530
rect 31164 16144 31198 16436
rect 31164 15050 31198 15342
rect 32222 19426 32256 19718
rect 35558 20920 35592 21212
rect 36616 25296 36650 25588
rect 36616 24202 36650 24494
rect 36616 23108 36650 23400
rect 36616 22014 36650 22306
rect 36616 20920 36650 21212
rect 37674 25296 37708 25588
rect 37674 24202 37708 24494
rect 37674 23108 37708 23400
rect 37674 22014 37708 22306
rect 37674 20920 37708 21212
rect 38732 25296 38766 25588
rect 42048 26756 42082 27048
rect 43106 31132 43140 31424
rect 43106 30038 43140 30330
rect 43106 28944 43140 29236
rect 43106 27850 43140 28142
rect 43106 26756 43140 27048
rect 44164 31132 44198 31424
rect 44164 30038 44198 30330
rect 44164 28944 44198 29236
rect 44164 27850 44198 28142
rect 44164 26756 44198 27048
rect 45222 31132 45256 31424
rect 48636 32612 48670 32904
rect 49694 36988 49728 37280
rect 49694 35894 49728 36186
rect 49694 34800 49728 35092
rect 49694 33706 49728 33998
rect 49694 32612 49728 32904
rect 50752 36988 50786 37280
rect 50752 35894 50786 36186
rect 50752 34800 50786 35092
rect 50752 33706 50786 33998
rect 50752 32612 50786 32904
rect 51810 36988 51844 37280
rect 55150 38442 55184 38734
rect 56208 42818 56242 43110
rect 56208 41724 56242 42016
rect 56208 40630 56242 40922
rect 56208 39536 56242 39828
rect 56208 38442 56242 38734
rect 57266 42818 57300 43110
rect 57266 41724 57300 42016
rect 57266 40630 57300 40922
rect 57266 39536 57300 39828
rect 57266 38442 57300 38734
rect 58324 42818 58358 43110
rect 58324 41724 58358 42016
rect 58324 40630 58358 40922
rect 58324 39536 58358 39828
rect 58324 38442 58358 38734
rect 59382 42818 59416 43110
rect 62508 42936 62542 43108
rect 59382 41724 59416 42016
rect 59382 40630 59416 40922
rect 59572 40204 59836 41772
rect 62194 41028 62288 42532
rect 62508 42242 62542 42414
rect 62508 41548 62542 41720
rect 62508 40854 62542 41026
rect 62508 40160 62542 40332
rect 63166 42936 63200 43108
rect 67844 43482 68066 43584
rect 63166 42242 63200 42414
rect 63166 41548 63200 41720
rect 63166 40854 63200 41026
rect 63166 40160 63200 40332
rect 63824 42936 63858 43108
rect 63824 42242 63858 42414
rect 63824 41548 63858 41720
rect 63824 40854 63858 41026
rect 63824 40160 63858 40332
rect 64482 42936 64516 43108
rect 65140 42936 65174 43108
rect 65798 42936 65832 43108
rect 64482 42242 64516 42414
rect 64482 41548 64516 41720
rect 64482 40854 64516 41026
rect 64482 40160 64516 40332
rect 65140 42242 65174 42414
rect 65140 41548 65174 41720
rect 65140 40854 65174 41026
rect 65140 40160 65174 40332
rect 66302 42938 66336 43110
rect 65798 42242 65832 42414
rect 65798 41548 65832 41720
rect 65798 40854 65832 41026
rect 65988 41030 66082 42534
rect 66302 42244 66336 42416
rect 66302 41550 66336 41722
rect 66302 40856 66336 41028
rect 65798 40160 65832 40332
rect 66302 40162 66336 40334
rect 66960 42938 66994 43110
rect 66960 42244 66994 42416
rect 66960 41550 66994 41722
rect 66960 40856 66994 41028
rect 66960 40162 66994 40334
rect 67618 42938 67652 43110
rect 67618 42244 67652 42416
rect 67618 41550 67652 41722
rect 67618 40856 67652 41028
rect 67618 40162 67652 40334
rect 68276 42938 68310 43110
rect 68934 42938 68968 43110
rect 71644 43472 71790 43584
rect 69592 42938 69626 43110
rect 70110 42952 70144 43124
rect 68276 42244 68310 42416
rect 68276 41550 68310 41722
rect 68276 40856 68310 41028
rect 68276 40162 68310 40334
rect 68934 42244 68968 42416
rect 69592 42244 69626 42416
rect 68934 41550 68968 41722
rect 68934 40856 68968 41028
rect 68934 40162 68968 40334
rect 69592 41550 69626 41722
rect 69592 40856 69626 41028
rect 69796 41044 69890 42548
rect 70110 42258 70144 42430
rect 70110 41564 70144 41736
rect 70110 40870 70144 41042
rect 69592 40162 69626 40334
rect 70110 40176 70144 40348
rect 70768 42952 70802 43124
rect 70768 42258 70802 42430
rect 70768 41564 70802 41736
rect 70768 40870 70802 41042
rect 70768 40176 70802 40348
rect 71426 42952 71460 43124
rect 71426 42258 71460 42430
rect 71426 41564 71460 41736
rect 71426 40870 71460 41042
rect 71426 40176 71460 40348
rect 72084 42952 72118 43124
rect 72742 42952 72776 43124
rect 73400 42952 73434 43124
rect 72084 42258 72118 42430
rect 72084 41564 72118 41736
rect 72084 40870 72118 41042
rect 72084 40176 72118 40348
rect 72742 42258 72776 42430
rect 72742 41564 72776 41736
rect 72742 40870 72776 41042
rect 72742 40176 72776 40348
rect 73400 42258 73434 42430
rect 73400 41564 73434 41736
rect 73400 40870 73434 41042
rect 73646 40970 73876 42876
rect 73400 40176 73434 40348
rect 59382 39536 59416 39828
rect 78570 39416 78774 39506
rect 80908 39444 81068 39522
rect 85084 39420 85284 39516
rect 59382 38442 59416 38734
rect 51810 35894 51844 36186
rect 51810 34800 51844 35092
rect 51810 33706 51844 33998
rect 51810 32612 51844 32904
rect 52868 36988 52902 37280
rect 52868 35894 52902 36186
rect 54092 37002 54126 37294
rect 55150 37002 55184 37294
rect 54092 35908 54126 36200
rect 55150 35908 55184 36200
rect 52868 34800 52902 35092
rect 53460 34564 53554 35760
rect 54092 34814 54126 35106
rect 55150 34814 55184 35106
rect 52868 33706 52902 33998
rect 52868 32612 52902 32904
rect 54092 33720 54126 34012
rect 55150 33720 55184 34012
rect 54092 32626 54126 32918
rect 45222 30038 45256 30330
rect 45222 28944 45256 29236
rect 45222 27850 45256 28142
rect 45222 26756 45256 27048
rect 46280 31132 46314 31424
rect 46280 30038 46314 30330
rect 47578 31154 47612 31446
rect 48636 31154 48670 31446
rect 47578 30060 47612 30352
rect 48636 30060 48670 30352
rect 46280 28944 46314 29236
rect 46946 28716 47040 29912
rect 47578 28966 47612 29258
rect 48636 28966 48670 29258
rect 46280 27850 46314 28142
rect 47578 27872 47612 28164
rect 48636 27872 48670 28164
rect 46280 26756 46314 27048
rect 47578 26778 47612 27070
rect 38732 24202 38766 24494
rect 38732 23108 38766 23400
rect 38732 22014 38766 22306
rect 38732 20920 38766 21212
rect 39790 25296 39824 25588
rect 39790 24202 39824 24494
rect 40990 25296 41024 25588
rect 42048 25296 42082 25588
rect 40990 24202 41024 24494
rect 42048 24202 42082 24494
rect 39790 23108 39824 23400
rect 40358 22858 40452 24054
rect 40990 23108 41024 23400
rect 42048 23108 42082 23400
rect 39790 22014 39824 22306
rect 39790 20920 39824 21212
rect 40990 22014 41024 22306
rect 42048 22014 42082 22306
rect 40990 20920 41024 21212
rect 32222 18332 32256 18624
rect 32222 17238 32256 17530
rect 32222 16144 32256 16436
rect 32222 15050 32256 15342
rect 33280 19426 33314 19718
rect 33280 18332 33314 18624
rect 34500 19432 34534 19724
rect 35558 19432 35592 19724
rect 34500 18338 34534 18630
rect 35558 18338 35592 18630
rect 33280 17238 33314 17530
rect 33868 16994 33962 18190
rect 34500 17244 34534 17536
rect 35558 17244 35592 17536
rect 33280 16144 33314 16436
rect 33280 15050 33314 15342
rect 34500 16150 34534 16442
rect 35558 16150 35592 16442
rect 34500 15056 34534 15348
rect 25710 12460 25744 12752
rect 25710 11366 25744 11658
rect 25710 10272 25744 10564
rect 25710 9178 25744 9470
rect 26768 13554 26802 13846
rect 26768 12460 26802 12752
rect 28000 13570 28034 13862
rect 29058 13570 29092 13862
rect 28000 12476 28034 12768
rect 29058 12476 29092 12768
rect 26768 11366 26802 11658
rect 27368 11132 27462 12328
rect 28000 11382 28034 11674
rect 29058 11382 29092 11674
rect 26768 10272 26802 10564
rect 28000 10288 28034 10580
rect 29058 10288 29092 10580
rect 26768 9178 26802 9470
rect 28000 9194 28034 9486
rect 19238 6568 19272 6860
rect 19238 5474 19272 5766
rect 19238 4380 19272 4672
rect 19238 3286 19272 3578
rect 20296 7662 20330 7954
rect 20296 6568 20330 6860
rect 21496 7646 21530 7938
rect 22554 7646 22588 7938
rect 21496 6552 21530 6844
rect 22554 6552 22588 6844
rect 20296 5474 20330 5766
rect 20864 5208 20958 6404
rect 21496 5458 21530 5750
rect 22554 5458 22588 5750
rect 20296 4380 20330 4672
rect 20296 3286 20330 3578
rect 21496 4364 21530 4656
rect 22554 4364 22588 4656
rect 21496 3270 21530 3562
rect 22554 3270 22588 3562
rect 23612 7646 23646 7938
rect 23612 6552 23646 6844
rect 23612 5458 23646 5750
rect 23612 4364 23646 4656
rect 23612 3270 23646 3562
rect 24670 7646 24704 7938
rect 24670 6552 24704 6844
rect 24670 5458 24704 5750
rect 24670 4364 24704 4656
rect 24670 3270 24704 3562
rect 25728 7646 25762 7938
rect 29058 9194 29092 9486
rect 30116 13570 30150 13862
rect 30116 12476 30150 12768
rect 30116 11382 30150 11674
rect 30116 10288 30150 10580
rect 30116 9194 30150 9486
rect 31174 13570 31208 13862
rect 31174 12476 31208 12768
rect 31174 11382 31208 11674
rect 31174 10288 31208 10580
rect 31174 9194 31208 9486
rect 32232 13570 32266 13862
rect 35558 15056 35592 15348
rect 36616 19432 36650 19724
rect 36616 18338 36650 18630
rect 36616 17244 36650 17536
rect 36616 16150 36650 16442
rect 36616 15056 36650 15348
rect 37674 19432 37708 19724
rect 37674 18338 37708 18630
rect 37674 17244 37708 17536
rect 37674 16150 37708 16442
rect 37674 15056 37708 15348
rect 38732 19432 38766 19724
rect 42048 20920 42082 21212
rect 43106 25296 43140 25588
rect 43106 24202 43140 24494
rect 43106 23108 43140 23400
rect 43106 22014 43140 22306
rect 43106 20920 43140 21212
rect 44164 25296 44198 25588
rect 44164 24202 44198 24494
rect 44164 23108 44198 23400
rect 44164 22014 44198 22306
rect 44164 20920 44198 21212
rect 45222 25296 45256 25588
rect 48636 26778 48670 27070
rect 49694 31154 49728 31446
rect 49694 30060 49728 30352
rect 49694 28966 49728 29258
rect 49694 27872 49728 28164
rect 49694 26778 49728 27070
rect 50752 31154 50786 31446
rect 50752 30060 50786 30352
rect 50752 28966 50786 29258
rect 50752 27872 50786 28164
rect 50752 26778 50786 27070
rect 51810 31154 51844 31446
rect 55150 32626 55184 32918
rect 56208 37002 56242 37294
rect 56208 35908 56242 36200
rect 56208 34814 56242 35106
rect 56208 33720 56242 34012
rect 56208 32626 56242 32918
rect 57266 37002 57300 37294
rect 57266 35908 57300 36200
rect 57266 34814 57300 35106
rect 57266 33720 57300 34012
rect 57266 32626 57300 32918
rect 58324 37002 58358 37294
rect 58324 35908 58358 36200
rect 58324 34814 58358 35106
rect 58324 33720 58358 34012
rect 58324 32626 58358 32918
rect 59382 37002 59416 37294
rect 59382 35908 59416 36200
rect 59382 34814 59416 35106
rect 59684 34446 59892 35834
rect 76760 35694 76908 38916
rect 77170 38922 77204 39094
rect 77170 38228 77204 38400
rect 77170 37534 77204 37706
rect 77170 36840 77204 37012
rect 77170 36146 77204 36318
rect 77170 35452 77204 35624
rect 77828 38922 77862 39094
rect 77828 38228 77862 38400
rect 77828 37534 77862 37706
rect 77828 36840 77862 37012
rect 77828 36146 77862 36318
rect 77828 35452 77862 35624
rect 78486 38922 78520 39094
rect 78486 38228 78520 38400
rect 78486 37534 78520 37706
rect 78486 36840 78520 37012
rect 78486 36146 78520 36318
rect 78486 35452 78520 35624
rect 79144 38922 79178 39094
rect 79802 38922 79836 39094
rect 79144 38228 79178 38400
rect 79144 37534 79178 37706
rect 79144 36840 79178 37012
rect 79144 36146 79178 36318
rect 79144 35452 79178 35624
rect 79802 38228 79836 38400
rect 79802 37534 79836 37706
rect 79802 36840 79836 37012
rect 79802 36146 79836 36318
rect 79802 35452 79836 35624
rect 80086 35688 80234 38910
rect 80496 38916 80530 39088
rect 80496 38222 80530 38394
rect 80496 37528 80530 37700
rect 80496 36834 80530 37006
rect 80496 36140 80530 36312
rect 80496 35446 80530 35618
rect 81154 38916 81188 39088
rect 81154 38222 81188 38394
rect 81154 37528 81188 37700
rect 81154 36834 81188 37006
rect 81154 36140 81188 36312
rect 81154 35446 81188 35618
rect 81812 38916 81846 39088
rect 81812 38222 81846 38394
rect 81812 37528 81846 37700
rect 81812 36834 81846 37006
rect 81812 36140 81846 36312
rect 81812 35446 81846 35618
rect 82470 38916 82504 39088
rect 82470 38222 82504 38394
rect 82470 37528 82504 37700
rect 82470 36834 82504 37006
rect 82470 36140 82504 36312
rect 82470 35446 82504 35618
rect 83128 38916 83162 39088
rect 83128 38222 83162 38394
rect 83128 37528 83162 37700
rect 83128 36834 83162 37006
rect 83128 36140 83162 36312
rect 83128 35446 83162 35618
rect 83396 35688 83544 38910
rect 83806 38916 83840 39088
rect 83806 38222 83840 38394
rect 83806 37528 83840 37700
rect 83806 36834 83840 37006
rect 83806 36140 83840 36312
rect 83806 35446 83840 35618
rect 84464 38916 84498 39088
rect 84464 38222 84498 38394
rect 84464 37528 84498 37700
rect 84464 36834 84498 37006
rect 84464 36140 84498 36312
rect 84464 35446 84498 35618
rect 85122 38916 85156 39088
rect 85122 38222 85156 38394
rect 85122 37528 85156 37700
rect 85122 36834 85156 37006
rect 85122 36140 85156 36312
rect 85122 35446 85156 35618
rect 85780 38916 85814 39088
rect 86438 38916 86472 39088
rect 85780 38222 85814 38394
rect 85780 37528 85814 37700
rect 85780 36834 85814 37006
rect 85780 36140 85814 36312
rect 85780 35446 85814 35618
rect 86438 38222 86472 38394
rect 86438 37528 86472 37700
rect 86438 36834 86472 37006
rect 86438 36140 86472 36312
rect 86438 35446 86472 35618
rect 86786 35656 86904 38988
rect 59382 33720 59416 34012
rect 59382 32626 59416 32918
rect 51810 30060 51844 30352
rect 51810 28966 51844 29258
rect 51810 27872 51844 28164
rect 51810 26778 51844 27070
rect 52868 31154 52902 31446
rect 52868 30060 52902 30352
rect 54092 31168 54126 31460
rect 55150 31168 55184 31460
rect 54092 30074 54126 30366
rect 55150 30074 55184 30366
rect 52868 28966 52902 29258
rect 53460 28730 53554 29926
rect 54092 28980 54126 29272
rect 55150 28980 55184 29272
rect 52868 27872 52902 28164
rect 52868 26778 52902 27070
rect 54092 27886 54126 28178
rect 55150 27886 55184 28178
rect 54092 26792 54126 27084
rect 45222 24202 45256 24494
rect 45222 23108 45256 23400
rect 45222 22014 45256 22306
rect 45222 20920 45256 21212
rect 46280 25296 46314 25588
rect 46280 24202 46314 24494
rect 47578 25318 47612 25610
rect 48636 25318 48670 25610
rect 47578 24224 47612 24516
rect 48636 24224 48670 24516
rect 46280 23108 46314 23400
rect 46946 22880 47040 24076
rect 47578 23130 47612 23422
rect 48636 23130 48670 23422
rect 46280 22014 46314 22306
rect 46280 20920 46314 21212
rect 47578 22036 47612 22328
rect 48636 22036 48670 22328
rect 47578 20942 47612 21234
rect 38732 18338 38766 18630
rect 38732 17244 38766 17536
rect 38732 16150 38766 16442
rect 38732 15056 38766 15348
rect 39790 19432 39824 19724
rect 39790 18338 39824 18630
rect 40990 19432 41024 19724
rect 42048 19432 42082 19724
rect 40990 18338 41024 18630
rect 42048 18338 42082 18630
rect 39790 17244 39824 17536
rect 40358 16994 40452 18190
rect 40990 17244 41024 17536
rect 42048 17244 42082 17536
rect 39790 16150 39824 16442
rect 39790 15056 39824 15348
rect 40990 16150 41024 16442
rect 42048 16150 42082 16442
rect 40990 15056 41024 15348
rect 32232 12476 32266 12768
rect 32232 11382 32266 11674
rect 32232 10288 32266 10580
rect 32232 9194 32266 9486
rect 33290 13570 33324 13862
rect 33290 12476 33324 12768
rect 34510 13576 34544 13868
rect 35568 13576 35602 13868
rect 34510 12482 34544 12774
rect 35568 12482 35602 12774
rect 33290 11382 33324 11674
rect 33878 11138 33972 12334
rect 34510 11388 34544 11680
rect 35568 11388 35602 11680
rect 33290 10288 33324 10580
rect 33290 9194 33324 9486
rect 34510 10294 34544 10586
rect 35568 10294 35602 10586
rect 34510 9200 34544 9492
rect 25728 6552 25762 6844
rect 25728 5458 25762 5750
rect 25728 4364 25762 4656
rect 25728 3270 25762 3562
rect 26786 7646 26820 7938
rect 26786 6552 26820 6844
rect 28018 7662 28052 7954
rect 29076 7662 29110 7954
rect 28018 6568 28052 6860
rect 29076 6568 29110 6860
rect 26786 5458 26820 5750
rect 27386 5224 27480 6420
rect 28018 5474 28052 5766
rect 29076 5474 29110 5766
rect 26786 4364 26820 4656
rect 26786 3270 26820 3562
rect 28018 4380 28052 4672
rect 29076 4380 29110 4672
rect 28018 3286 28052 3578
rect 29076 3286 29110 3578
rect 30134 7662 30168 7954
rect 30134 6568 30168 6860
rect 30134 5474 30168 5766
rect 30134 4380 30168 4672
rect 30134 3286 30168 3578
rect 31192 7662 31226 7954
rect 31192 6568 31226 6860
rect 31192 5474 31226 5766
rect 31192 4380 31226 4672
rect 31192 3286 31226 3578
rect 32250 7662 32284 7954
rect 35568 9200 35602 9492
rect 36626 13576 36660 13868
rect 36626 12482 36660 12774
rect 36626 11388 36660 11680
rect 36626 10294 36660 10586
rect 36626 9200 36660 9492
rect 37684 13576 37718 13868
rect 37684 12482 37718 12774
rect 37684 11388 37718 11680
rect 37684 10294 37718 10586
rect 37684 9200 37718 9492
rect 38742 13576 38776 13868
rect 42048 15056 42082 15348
rect 43106 19432 43140 19724
rect 43106 18338 43140 18630
rect 43106 17244 43140 17536
rect 43106 16150 43140 16442
rect 43106 15056 43140 15348
rect 44164 19432 44198 19724
rect 44164 18338 44198 18630
rect 44164 17244 44198 17536
rect 44164 16150 44198 16442
rect 44164 15056 44198 15348
rect 45222 19432 45256 19724
rect 48636 20942 48670 21234
rect 49694 25318 49728 25610
rect 49694 24224 49728 24516
rect 49694 23130 49728 23422
rect 49694 22036 49728 22328
rect 49694 20942 49728 21234
rect 50752 25318 50786 25610
rect 50752 24224 50786 24516
rect 50752 23130 50786 23422
rect 50752 22036 50786 22328
rect 50752 20942 50786 21234
rect 51810 25318 51844 25610
rect 55150 26792 55184 27084
rect 56208 31168 56242 31460
rect 56208 30074 56242 30366
rect 56208 28980 56242 29272
rect 56208 27886 56242 28178
rect 56208 26792 56242 27084
rect 57266 31168 57300 31460
rect 57266 30074 57300 30366
rect 57266 28980 57300 29272
rect 57266 27886 57300 28178
rect 57266 26792 57300 27084
rect 58324 31168 58358 31460
rect 58324 30074 58358 30366
rect 58324 28980 58358 29272
rect 58324 27886 58358 28178
rect 58324 26792 58358 27084
rect 59382 31168 59416 31460
rect 59382 30074 59416 30366
rect 59382 28980 59416 29272
rect 59382 27886 59416 28178
rect 59642 28426 59974 29896
rect 59382 26792 59416 27084
rect 51810 24224 51844 24516
rect 51810 23130 51844 23422
rect 51810 22036 51844 22328
rect 51810 20942 51844 21234
rect 52868 25318 52902 25610
rect 52868 24224 52902 24516
rect 54092 25332 54126 25624
rect 55150 25332 55184 25624
rect 54092 24238 54126 24530
rect 55150 24238 55184 24530
rect 52868 23130 52902 23422
rect 53460 22894 53554 24090
rect 54092 23144 54126 23436
rect 55150 23144 55184 23436
rect 52868 22036 52902 22328
rect 52868 20942 52902 21234
rect 54092 22050 54126 22342
rect 55150 22050 55184 22342
rect 54092 20956 54126 21248
rect 45222 18338 45256 18630
rect 45222 17244 45256 17536
rect 45222 16150 45256 16442
rect 45222 15056 45256 15348
rect 46280 19432 46314 19724
rect 46280 18338 46314 18630
rect 47578 19454 47612 19746
rect 48636 19454 48670 19746
rect 47578 18360 47612 18652
rect 48636 18360 48670 18652
rect 46280 17244 46314 17536
rect 46946 17016 47040 18212
rect 47578 17266 47612 17558
rect 48636 17266 48670 17558
rect 46280 16150 46314 16442
rect 46280 15056 46314 15348
rect 47578 16172 47612 16464
rect 48636 16172 48670 16464
rect 47578 15078 47612 15370
rect 38742 12482 38776 12774
rect 38742 11388 38776 11680
rect 38742 10294 38776 10586
rect 38742 9200 38776 9492
rect 39800 13576 39834 13868
rect 39800 12482 39834 12774
rect 41000 13576 41034 13868
rect 42058 13576 42092 13868
rect 41000 12482 41034 12774
rect 42058 12482 42092 12774
rect 39800 11388 39834 11680
rect 40368 11138 40462 12334
rect 41000 11388 41034 11680
rect 42058 11388 42092 11680
rect 39800 10294 39834 10586
rect 39800 9200 39834 9492
rect 41000 10294 41034 10586
rect 42058 10294 42092 10586
rect 41000 9200 41034 9492
rect 32250 6568 32284 6860
rect 32250 5474 32284 5766
rect 32250 4380 32284 4672
rect 32250 3286 32284 3578
rect 33308 7662 33342 7954
rect 33308 6568 33342 6860
rect 34528 7668 34562 7960
rect 35586 7668 35620 7960
rect 34528 6574 34562 6866
rect 35586 6574 35620 6866
rect 33308 5474 33342 5766
rect 33896 5230 33990 6426
rect 34528 5480 34562 5772
rect 35586 5480 35620 5772
rect 33308 4380 33342 4672
rect 33308 3286 33342 3578
rect 34528 4386 34562 4678
rect 35586 4386 35620 4678
rect 34528 3292 34562 3584
rect 35586 3292 35620 3584
rect 36644 7668 36678 7960
rect 36644 6574 36678 6866
rect 36644 5480 36678 5772
rect 36644 4386 36678 4678
rect 36644 3292 36678 3584
rect 37702 7668 37736 7960
rect 37702 6574 37736 6866
rect 37702 5480 37736 5772
rect 37702 4386 37736 4678
rect 37702 3292 37736 3584
rect 38760 7668 38794 7960
rect 42058 9200 42092 9492
rect 43116 13576 43150 13868
rect 43116 12482 43150 12774
rect 43116 11388 43150 11680
rect 43116 10294 43150 10586
rect 43116 9200 43150 9492
rect 44174 13576 44208 13868
rect 44174 12482 44208 12774
rect 44174 11388 44208 11680
rect 44174 10294 44208 10586
rect 44174 9200 44208 9492
rect 45232 13576 45266 13868
rect 48636 15078 48670 15370
rect 49694 19454 49728 19746
rect 49694 18360 49728 18652
rect 49694 17266 49728 17558
rect 49694 16172 49728 16464
rect 49694 15078 49728 15370
rect 50752 19454 50786 19746
rect 50752 18360 50786 18652
rect 50752 17266 50786 17558
rect 50752 16172 50786 16464
rect 50752 15078 50786 15370
rect 51810 19454 51844 19746
rect 55150 20956 55184 21248
rect 56208 25332 56242 25624
rect 56208 24238 56242 24530
rect 56208 23144 56242 23436
rect 56208 22050 56242 22342
rect 56208 20956 56242 21248
rect 57266 25332 57300 25624
rect 57266 24238 57300 24530
rect 57266 23144 57300 23436
rect 57266 22050 57300 22342
rect 57266 20956 57300 21248
rect 58324 25332 58358 25624
rect 67700 26216 68180 26314
rect 94062 26190 94392 26270
rect 58324 24238 58358 24530
rect 58324 23144 58358 23436
rect 58324 22050 58358 22342
rect 58324 20956 58358 21248
rect 59382 25332 59416 25624
rect 59382 24238 59416 24530
rect 62112 25276 62146 25568
rect 63170 25276 63204 25568
rect 59382 23144 59416 23436
rect 59614 22696 59864 24250
rect 62112 24182 62146 24474
rect 63170 24182 63204 24474
rect 61480 22838 61574 24034
rect 62112 23088 62146 23380
rect 63170 23088 63204 23380
rect 59382 22050 59416 22342
rect 59382 20956 59416 21248
rect 62112 21994 62146 22286
rect 63170 21994 63204 22286
rect 62112 20900 62146 21192
rect 63170 20900 63204 21192
rect 64228 25276 64262 25568
rect 64228 24182 64262 24474
rect 64228 23088 64262 23380
rect 64228 21994 64262 22286
rect 64228 20900 64262 21192
rect 65286 25276 65320 25568
rect 65286 24182 65320 24474
rect 65286 23088 65320 23380
rect 65286 21994 65320 22286
rect 65286 20900 65320 21192
rect 66344 25276 66378 25568
rect 66344 24182 66378 24474
rect 66344 23088 66378 23380
rect 66344 21994 66378 22286
rect 66344 20900 66378 21192
rect 67402 25276 67436 25568
rect 67402 24182 67436 24474
rect 68574 25274 68608 25566
rect 69632 25274 69666 25566
rect 68574 24180 68608 24472
rect 69632 24180 69666 24472
rect 67402 23088 67436 23380
rect 67942 22836 68036 24032
rect 68574 23086 68608 23378
rect 69632 23086 69666 23378
rect 67402 21994 67436 22286
rect 67402 20900 67436 21192
rect 68574 21992 68608 22284
rect 69632 21992 69666 22284
rect 68574 20898 68608 21190
rect 69632 20898 69666 21190
rect 70690 25274 70724 25566
rect 70690 24180 70724 24472
rect 70690 23086 70724 23378
rect 70690 21992 70724 22284
rect 51810 18360 51844 18652
rect 51810 17266 51844 17558
rect 51810 16172 51844 16464
rect 51810 15078 51844 15370
rect 52868 19454 52902 19746
rect 52868 18360 52902 18652
rect 54092 19468 54126 19760
rect 55150 19468 55184 19760
rect 54092 18374 54126 18666
rect 55150 18374 55184 18666
rect 52868 17266 52902 17558
rect 53460 17030 53554 18226
rect 54092 17280 54126 17572
rect 55150 17280 55184 17572
rect 52868 16172 52902 16464
rect 52868 15078 52902 15370
rect 54092 16186 54126 16478
rect 55150 16186 55184 16478
rect 54092 15092 54126 15384
rect 45232 12482 45266 12774
rect 45232 11388 45266 11680
rect 45232 10294 45266 10586
rect 45232 9200 45266 9492
rect 46290 13576 46324 13868
rect 46290 12482 46324 12774
rect 47588 13598 47622 13890
rect 48646 13598 48680 13890
rect 47588 12504 47622 12796
rect 48646 12504 48680 12796
rect 46290 11388 46324 11680
rect 46956 11160 47050 12356
rect 47588 11410 47622 11702
rect 48646 11410 48680 11702
rect 46290 10294 46324 10586
rect 46290 9200 46324 9492
rect 47588 10316 47622 10608
rect 48646 10316 48680 10608
rect 47588 9222 47622 9514
rect 38760 6574 38794 6866
rect 38760 5480 38794 5772
rect 38760 4386 38794 4678
rect 38760 3292 38794 3584
rect 39818 7668 39852 7960
rect 39818 6574 39852 6866
rect 41018 7668 41052 7960
rect 42076 7668 42110 7960
rect 41018 6574 41052 6866
rect 42076 6574 42110 6866
rect 39818 5480 39852 5772
rect 39818 4386 39852 4678
rect 39818 3292 39852 3584
rect 40386 5230 40480 6426
rect 41018 5480 41052 5772
rect 42076 5480 42110 5772
rect 41018 4386 41052 4678
rect 42076 4386 42110 4678
rect 41018 3292 41052 3584
rect 42076 3292 42110 3584
rect 43134 7668 43168 7960
rect 43134 6574 43168 6866
rect 43134 5480 43168 5772
rect 43134 4386 43168 4678
rect 43134 3292 43168 3584
rect 44192 7668 44226 7960
rect 44192 6574 44226 6866
rect 44192 5480 44226 5772
rect 44192 4386 44226 4678
rect 44192 3292 44226 3584
rect 45250 7668 45284 7960
rect 48646 9222 48680 9514
rect 49704 13598 49738 13890
rect 49704 12504 49738 12796
rect 49704 11410 49738 11702
rect 49704 10316 49738 10608
rect 49704 9222 49738 9514
rect 50762 13598 50796 13890
rect 55150 15092 55184 15384
rect 56208 19468 56242 19760
rect 56208 18374 56242 18666
rect 56208 17280 56242 17572
rect 56208 16186 56242 16478
rect 56208 15092 56242 15384
rect 57266 19468 57300 19760
rect 57266 18374 57300 18666
rect 57266 17280 57300 17572
rect 57266 16186 57300 16478
rect 57266 15092 57300 15384
rect 58324 19468 58358 19760
rect 70690 20898 70724 21190
rect 71748 25274 71782 25566
rect 71748 24180 71782 24472
rect 71748 23086 71782 23378
rect 71748 21992 71782 22284
rect 71748 20898 71782 21190
rect 72806 25274 72840 25566
rect 72806 24180 72840 24472
rect 72806 23086 72840 23378
rect 72806 21992 72840 22284
rect 72806 20898 72840 21190
rect 73864 25274 73898 25566
rect 73864 24180 73898 24472
rect 75268 25248 75302 25540
rect 76326 25248 76360 25540
rect 75268 24154 75302 24446
rect 76326 24154 76360 24446
rect 73864 23086 73898 23378
rect 74636 22810 74730 24006
rect 75268 23060 75302 23352
rect 76326 23060 76360 23352
rect 73864 21992 73898 22284
rect 73864 20898 73898 21190
rect 75268 21966 75302 22258
rect 76326 21966 76360 22258
rect 75268 20872 75302 21164
rect 76326 20872 76360 21164
rect 77384 25248 77418 25540
rect 77384 24154 77418 24446
rect 77384 23060 77418 23352
rect 77384 21966 77418 22258
rect 77384 20872 77418 21164
rect 78442 25248 78476 25540
rect 78442 24154 78476 24446
rect 78442 23060 78476 23352
rect 78442 21966 78476 22258
rect 78442 20872 78476 21164
rect 79500 25248 79534 25540
rect 79500 24154 79534 24446
rect 79500 23060 79534 23352
rect 79500 21966 79534 22258
rect 79500 20872 79534 21164
rect 80558 25248 80592 25540
rect 80558 24154 80592 24446
rect 81730 25246 81764 25538
rect 82788 25246 82822 25538
rect 81730 24152 81764 24444
rect 82788 24152 82822 24444
rect 80558 23060 80592 23352
rect 81098 22808 81192 24004
rect 81730 23058 81764 23350
rect 82788 23058 82822 23350
rect 80558 21966 80592 22258
rect 80558 20872 80592 21164
rect 81730 21964 81764 22256
rect 82788 21964 82822 22256
rect 81730 20870 81764 21162
rect 82788 20870 82822 21162
rect 83846 25246 83880 25538
rect 83846 24152 83880 24444
rect 83846 23058 83880 23350
rect 83846 21964 83880 22256
rect 83846 20870 83880 21162
rect 84904 25246 84938 25538
rect 84904 24152 84938 24444
rect 84904 23058 84938 23350
rect 84904 21964 84938 22256
rect 84904 20870 84938 21162
rect 85962 25246 85996 25538
rect 85962 24152 85996 24444
rect 85962 23058 85996 23350
rect 85962 21964 85996 22256
rect 85962 20870 85996 21162
rect 87020 25246 87054 25538
rect 87020 24152 87054 24444
rect 88502 25240 88536 25532
rect 89560 25240 89594 25532
rect 88502 24146 88536 24438
rect 89560 24146 89594 24438
rect 87020 23058 87054 23350
rect 87870 22802 87964 23998
rect 88502 23052 88536 23344
rect 89560 23052 89594 23344
rect 87020 21964 87054 22256
rect 87020 20870 87054 21162
rect 88502 21958 88536 22250
rect 89560 21958 89594 22250
rect 88502 20864 88536 21156
rect 89560 20864 89594 21156
rect 90618 25240 90652 25532
rect 90618 24146 90652 24438
rect 90618 23052 90652 23344
rect 90618 21958 90652 22250
rect 90618 20864 90652 21156
rect 91676 25240 91710 25532
rect 91676 24146 91710 24438
rect 91676 23052 91710 23344
rect 91676 21958 91710 22250
rect 91676 20864 91710 21156
rect 92734 25240 92768 25532
rect 92734 24146 92768 24438
rect 92734 23052 92768 23344
rect 92734 21958 92768 22250
rect 92734 20864 92768 21156
rect 93792 25240 93826 25532
rect 93792 24146 93826 24438
rect 94964 25238 94998 25530
rect 96022 25238 96056 25530
rect 94964 24144 94998 24436
rect 96022 24144 96056 24436
rect 93792 23052 93826 23344
rect 94332 22800 94426 23996
rect 94964 23050 94998 23342
rect 96022 23050 96056 23342
rect 93792 21958 93826 22250
rect 93792 20864 93826 21156
rect 94964 21956 94998 22248
rect 96022 21956 96056 22248
rect 94964 20862 94998 21154
rect 96022 20862 96056 21154
rect 97080 25238 97114 25530
rect 97080 24144 97114 24436
rect 97080 23050 97114 23342
rect 97080 21956 97114 22248
rect 97080 20862 97114 21154
rect 98138 25238 98172 25530
rect 98138 24144 98172 24436
rect 98138 23050 98172 23342
rect 98138 21956 98172 22248
rect 98138 20862 98172 21154
rect 99196 25238 99230 25530
rect 99196 24144 99230 24436
rect 99196 23050 99230 23342
rect 99196 21956 99230 22248
rect 99196 20862 99230 21154
rect 100254 25238 100288 25530
rect 100254 24144 100288 24436
rect 100254 23050 100288 23342
rect 100254 21956 100288 22248
rect 100254 20862 100288 21154
rect 100786 21760 101232 25032
rect 101232 21760 101276 25032
rect 58324 18374 58358 18666
rect 58324 17280 58358 17572
rect 58324 16186 58358 16478
rect 58324 15092 58358 15384
rect 59382 19468 59416 19760
rect 62118 19438 62152 19730
rect 63176 19438 63210 19730
rect 59382 18374 59416 18666
rect 59382 17280 59416 17572
rect 59698 16980 59892 18464
rect 62118 18344 62152 18636
rect 63176 18344 63210 18636
rect 61486 17000 61580 18196
rect 62118 17250 62152 17542
rect 63176 17250 63210 17542
rect 59382 16186 59416 16478
rect 59382 15092 59416 15384
rect 62118 16156 62152 16448
rect 63176 16156 63210 16448
rect 62118 15062 62152 15354
rect 63176 15062 63210 15354
rect 64234 19438 64268 19730
rect 64234 18344 64268 18636
rect 64234 17250 64268 17542
rect 64234 16156 64268 16448
rect 64234 15062 64268 15354
rect 65292 19438 65326 19730
rect 65292 18344 65326 18636
rect 65292 17250 65326 17542
rect 65292 16156 65326 16448
rect 65292 15062 65326 15354
rect 66350 19438 66384 19730
rect 66350 18344 66384 18636
rect 66350 17250 66384 17542
rect 66350 16156 66384 16448
rect 66350 15062 66384 15354
rect 67408 19438 67442 19730
rect 67408 18344 67442 18636
rect 68582 19450 68616 19742
rect 69640 19450 69674 19742
rect 68582 18356 68616 18648
rect 69640 18356 69674 18648
rect 67408 17250 67442 17542
rect 67950 17012 68044 18208
rect 68582 17262 68616 17554
rect 69640 17262 69674 17554
rect 67408 16156 67442 16448
rect 67408 15062 67442 15354
rect 68582 16168 68616 16460
rect 69640 16168 69674 16460
rect 68582 15074 68616 15366
rect 69640 15074 69674 15366
rect 70698 19450 70732 19742
rect 70698 18356 70732 18648
rect 70698 17262 70732 17554
rect 70698 16168 70732 16460
rect 70698 15074 70732 15366
rect 71756 19450 71790 19742
rect 71756 18356 71790 18648
rect 71756 17262 71790 17554
rect 71756 16168 71790 16460
rect 71756 15074 71790 15366
rect 72814 19450 72848 19742
rect 72814 18356 72848 18648
rect 72814 17262 72848 17554
rect 72814 16168 72848 16460
rect 72814 15074 72848 15366
rect 73872 19450 73906 19742
rect 73872 18356 73906 18648
rect 75274 19410 75308 19702
rect 76332 19410 76366 19702
rect 75274 18316 75308 18608
rect 76332 18316 76366 18608
rect 73872 17262 73906 17554
rect 74642 16972 74736 18168
rect 75274 17222 75308 17514
rect 76332 17222 76366 17514
rect 73872 16168 73906 16460
rect 73872 15074 73906 15366
rect 75274 16128 75308 16420
rect 76332 16128 76366 16420
rect 75274 15034 75308 15326
rect 76332 15034 76366 15326
rect 77390 19410 77424 19702
rect 77390 18316 77424 18608
rect 77390 17222 77424 17514
rect 77390 16128 77424 16420
rect 50762 12504 50796 12796
rect 50762 11410 50796 11702
rect 50762 10316 50796 10608
rect 50762 9222 50796 9514
rect 51820 13598 51854 13890
rect 51820 12504 51854 12796
rect 51820 11410 51854 11702
rect 51820 10316 51854 10608
rect 51820 9222 51854 9514
rect 52878 13598 52912 13890
rect 52878 12504 52912 12796
rect 54102 13612 54136 13904
rect 55160 13612 55194 13904
rect 54102 12518 54136 12810
rect 55160 12518 55194 12810
rect 52878 11410 52912 11702
rect 53470 11174 53564 12370
rect 54102 11424 54136 11716
rect 55160 11424 55194 11716
rect 52878 10316 52912 10608
rect 52878 9222 52912 9514
rect 54102 10330 54136 10622
rect 55160 10330 55194 10622
rect 54102 9236 54136 9528
rect 45250 6574 45284 6866
rect 45250 5480 45284 5772
rect 45250 4386 45284 4678
rect 45250 3292 45284 3584
rect 46308 7668 46342 7960
rect 46308 6574 46342 6866
rect 47606 7690 47640 7982
rect 48664 7690 48698 7982
rect 47606 6596 47640 6888
rect 48664 6596 48698 6888
rect 46308 5480 46342 5772
rect 46974 5252 47068 6448
rect 47606 5502 47640 5794
rect 48664 5502 48698 5794
rect 46308 4386 46342 4678
rect 46308 3292 46342 3584
rect 47606 4408 47640 4700
rect 48664 4408 48698 4700
rect 47606 3314 47640 3606
rect 48664 3314 48698 3606
rect 49722 7690 49756 7982
rect 49722 6596 49756 6888
rect 49722 5502 49756 5794
rect 49722 4408 49756 4700
rect 49722 3314 49756 3606
rect 50780 7690 50814 7982
rect 50780 6596 50814 6888
rect 50780 5502 50814 5794
rect 50780 4408 50814 4700
rect 50780 3314 50814 3606
rect 51838 7690 51872 7982
rect 55160 9236 55194 9528
rect 56218 13612 56252 13904
rect 56218 12518 56252 12810
rect 56218 11424 56252 11716
rect 56218 10330 56252 10622
rect 56218 9236 56252 9528
rect 57276 13612 57310 13904
rect 57276 12518 57310 12810
rect 57276 11424 57310 11716
rect 57276 10330 57310 10622
rect 57276 9236 57310 9528
rect 58334 13612 58368 13904
rect 77390 15034 77424 15326
rect 78448 19410 78482 19702
rect 78448 18316 78482 18608
rect 78448 17222 78482 17514
rect 78448 16128 78482 16420
rect 78448 15034 78482 15326
rect 79506 19410 79540 19702
rect 79506 18316 79540 18608
rect 79506 17222 79540 17514
rect 79506 16128 79540 16420
rect 79506 15034 79540 15326
rect 80564 19410 80598 19702
rect 80564 18316 80598 18608
rect 81738 19422 81772 19714
rect 82796 19422 82830 19714
rect 81738 18328 81772 18620
rect 82796 18328 82830 18620
rect 80564 17222 80598 17514
rect 81106 16984 81200 18180
rect 81738 17234 81772 17526
rect 82796 17234 82830 17526
rect 80564 16128 80598 16420
rect 80564 15034 80598 15326
rect 81738 16140 81772 16432
rect 82796 16140 82830 16432
rect 81738 15046 81772 15338
rect 82796 15046 82830 15338
rect 83854 19422 83888 19714
rect 83854 18328 83888 18620
rect 83854 17234 83888 17526
rect 83854 16140 83888 16432
rect 83854 15046 83888 15338
rect 84912 19422 84946 19714
rect 84912 18328 84946 18620
rect 84912 17234 84946 17526
rect 84912 16140 84946 16432
rect 84912 15046 84946 15338
rect 85970 19422 86004 19714
rect 85970 18328 86004 18620
rect 85970 17234 86004 17526
rect 85970 16140 86004 16432
rect 85970 15046 86004 15338
rect 87028 19422 87062 19714
rect 87028 18328 87062 18620
rect 88508 19402 88542 19694
rect 89566 19402 89600 19694
rect 88508 18308 88542 18600
rect 89566 18308 89600 18600
rect 87028 17234 87062 17526
rect 87876 16964 87970 18160
rect 88508 17214 88542 17506
rect 89566 17214 89600 17506
rect 87028 16140 87062 16432
rect 87028 15046 87062 15338
rect 88508 16120 88542 16412
rect 89566 16120 89600 16412
rect 88508 15026 88542 15318
rect 89566 15026 89600 15318
rect 90624 19402 90658 19694
rect 90624 18308 90658 18600
rect 90624 17214 90658 17506
rect 90624 16120 90658 16412
rect 90624 15026 90658 15318
rect 91682 19402 91716 19694
rect 91682 18308 91716 18600
rect 91682 17214 91716 17506
rect 91682 16120 91716 16412
rect 91682 15026 91716 15318
rect 92740 19402 92774 19694
rect 92740 18308 92774 18600
rect 92740 17214 92774 17506
rect 92740 16120 92774 16412
rect 92740 15026 92774 15318
rect 93798 19402 93832 19694
rect 93798 18308 93832 18600
rect 94972 19414 95006 19706
rect 96030 19414 96064 19706
rect 94972 18320 95006 18612
rect 96030 18320 96064 18612
rect 93798 17214 93832 17506
rect 94340 16976 94434 18172
rect 94972 17226 95006 17518
rect 96030 17226 96064 17518
rect 93798 16120 93832 16412
rect 93798 15026 93832 15318
rect 94972 16132 95006 16424
rect 96030 16132 96064 16424
rect 94972 15038 95006 15330
rect 96030 15038 96064 15330
rect 97088 19414 97122 19706
rect 97088 18320 97122 18612
rect 97088 17226 97122 17518
rect 97088 16132 97122 16424
rect 97088 15038 97122 15330
rect 98146 19414 98180 19706
rect 98146 18320 98180 18612
rect 98146 17226 98180 17518
rect 98146 16132 98180 16424
rect 98146 15038 98180 15330
rect 99204 19414 99238 19706
rect 99204 18320 99238 18612
rect 99204 17226 99238 17518
rect 99204 16132 99238 16424
rect 99204 15038 99238 15330
rect 100262 19414 100296 19706
rect 100262 18320 100296 18612
rect 100262 17226 100296 17518
rect 100262 16132 100296 16424
rect 100262 15038 100296 15330
rect 100742 15392 101120 18976
rect 58334 12518 58368 12810
rect 58334 11424 58368 11716
rect 58334 10330 58368 10622
rect 58334 9236 58368 9528
rect 59392 13612 59426 13904
rect 59392 12518 59426 12810
rect 62118 13580 62152 13872
rect 63176 13580 63210 13872
rect 59392 11424 59426 11716
rect 59698 11168 59934 12542
rect 62118 12486 62152 12778
rect 63176 12486 63210 12778
rect 61486 11142 61580 12338
rect 62118 11392 62152 11684
rect 63176 11392 63210 11684
rect 59392 10330 59426 10622
rect 59392 9236 59426 9528
rect 62118 10298 62152 10590
rect 63176 10298 63210 10590
rect 62118 9204 62152 9496
rect 63176 9204 63210 9496
rect 64234 13580 64268 13872
rect 64234 12486 64268 12778
rect 64234 11392 64268 11684
rect 64234 10298 64268 10590
rect 64234 9204 64268 9496
rect 65292 13580 65326 13872
rect 65292 12486 65326 12778
rect 65292 11392 65326 11684
rect 65292 10298 65326 10590
rect 65292 9204 65326 9496
rect 66350 13580 66384 13872
rect 66350 12486 66384 12778
rect 66350 11392 66384 11684
rect 66350 10298 66384 10590
rect 66350 9204 66384 9496
rect 67408 13580 67442 13872
rect 67408 12486 67442 12778
rect 68586 13578 68620 13870
rect 69644 13578 69678 13870
rect 68586 12484 68620 12776
rect 69644 12484 69678 12776
rect 67408 11392 67442 11684
rect 67954 11140 68048 12336
rect 68586 11390 68620 11682
rect 69644 11390 69678 11682
rect 67408 10298 67442 10590
rect 67408 9204 67442 9496
rect 68586 10296 68620 10588
rect 69644 10296 69678 10588
rect 68586 9202 68620 9494
rect 69644 9202 69678 9494
rect 70702 13578 70736 13870
rect 70702 12484 70736 12776
rect 70702 11390 70736 11682
rect 70702 10296 70736 10588
rect 51838 6596 51872 6888
rect 51838 5502 51872 5794
rect 51838 4408 51872 4700
rect 51838 3314 51872 3606
rect 52896 7690 52930 7982
rect 52896 6596 52930 6888
rect 54120 7704 54154 7996
rect 55178 7704 55212 7996
rect 54120 6610 54154 6902
rect 55178 6610 55212 6902
rect 52896 5502 52930 5794
rect 53488 5266 53582 6462
rect 54120 5516 54154 5808
rect 55178 5516 55212 5808
rect 52896 4408 52930 4700
rect 52896 3314 52930 3606
rect 54120 4422 54154 4714
rect 55178 4422 55212 4714
rect 54120 3328 54154 3620
rect 55178 3328 55212 3620
rect 56236 7704 56270 7996
rect 56236 6610 56270 6902
rect 56236 5516 56270 5808
rect 56236 4422 56270 4714
rect 56236 3328 56270 3620
rect 57294 7704 57328 7996
rect 57294 6610 57328 6902
rect 57294 5516 57328 5808
rect 57294 4422 57328 4714
rect 57294 3328 57328 3620
rect 58352 7704 58386 7996
rect 70702 9202 70736 9494
rect 71760 13578 71794 13870
rect 71760 12484 71794 12776
rect 71760 11390 71794 11682
rect 71760 10296 71794 10588
rect 71760 9202 71794 9494
rect 72818 13578 72852 13870
rect 72818 12484 72852 12776
rect 72818 11390 72852 11682
rect 72818 10296 72852 10588
rect 72818 9202 72852 9494
rect 73876 13578 73910 13870
rect 73876 12484 73910 12776
rect 75274 13552 75308 13844
rect 76332 13552 76366 13844
rect 75274 12458 75308 12750
rect 76332 12458 76366 12750
rect 73876 11390 73910 11682
rect 74642 11114 74736 12310
rect 75274 11364 75308 11656
rect 76332 11364 76366 11656
rect 73876 10296 73910 10588
rect 73876 9202 73910 9494
rect 75274 10270 75308 10562
rect 76332 10270 76366 10562
rect 75274 9176 75308 9468
rect 76332 9176 76366 9468
rect 77390 13552 77424 13844
rect 77390 12458 77424 12750
rect 77390 11364 77424 11656
rect 77390 10270 77424 10562
rect 77390 9176 77424 9468
rect 78448 13552 78482 13844
rect 78448 12458 78482 12750
rect 78448 11364 78482 11656
rect 78448 10270 78482 10562
rect 78448 9176 78482 9468
rect 79506 13552 79540 13844
rect 79506 12458 79540 12750
rect 79506 11364 79540 11656
rect 79506 10270 79540 10562
rect 79506 9176 79540 9468
rect 80564 13552 80598 13844
rect 80564 12458 80598 12750
rect 81742 13550 81776 13842
rect 82800 13550 82834 13842
rect 81742 12456 81776 12748
rect 82800 12456 82834 12748
rect 80564 11364 80598 11656
rect 81110 11112 81204 12308
rect 81742 11362 81776 11654
rect 82800 11362 82834 11654
rect 80564 10270 80598 10562
rect 80564 9176 80598 9468
rect 81742 10268 81776 10560
rect 82800 10268 82834 10560
rect 81742 9174 81776 9466
rect 82800 9174 82834 9466
rect 83858 13550 83892 13842
rect 83858 12456 83892 12748
rect 83858 11362 83892 11654
rect 83858 10268 83892 10560
rect 83858 9174 83892 9466
rect 84916 13550 84950 13842
rect 84916 12456 84950 12748
rect 84916 11362 84950 11654
rect 84916 10268 84950 10560
rect 84916 9174 84950 9466
rect 85974 13550 86008 13842
rect 85974 12456 86008 12748
rect 85974 11362 86008 11654
rect 85974 10268 86008 10560
rect 85974 9174 86008 9466
rect 87032 13550 87066 13842
rect 87032 12456 87066 12748
rect 88508 13544 88542 13836
rect 89566 13544 89600 13836
rect 88508 12450 88542 12742
rect 89566 12450 89600 12742
rect 87032 11362 87066 11654
rect 87876 11106 87970 12302
rect 88508 11356 88542 11648
rect 89566 11356 89600 11648
rect 87032 10268 87066 10560
rect 87032 9174 87066 9466
rect 88508 10262 88542 10554
rect 89566 10262 89600 10554
rect 88508 9168 88542 9460
rect 89566 9168 89600 9460
rect 90624 13544 90658 13836
rect 90624 12450 90658 12742
rect 90624 11356 90658 11648
rect 90624 10262 90658 10554
rect 90624 9168 90658 9460
rect 91682 13544 91716 13836
rect 91682 12450 91716 12742
rect 91682 11356 91716 11648
rect 91682 10262 91716 10554
rect 91682 9168 91716 9460
rect 92740 13544 92774 13836
rect 92740 12450 92774 12742
rect 92740 11356 92774 11648
rect 92740 10262 92774 10554
rect 92740 9168 92774 9460
rect 93798 13544 93832 13836
rect 93798 12450 93832 12742
rect 94976 13542 95010 13834
rect 96034 13542 96068 13834
rect 94976 12448 95010 12740
rect 96034 12448 96068 12740
rect 93798 11356 93832 11648
rect 94344 11104 94438 12300
rect 94976 11354 95010 11646
rect 96034 11354 96068 11646
rect 93798 10262 93832 10554
rect 93798 9168 93832 9460
rect 94976 10260 95010 10552
rect 96034 10260 96068 10552
rect 94976 9166 95010 9458
rect 96034 9166 96068 9458
rect 97092 13542 97126 13834
rect 97092 12448 97126 12740
rect 97092 11354 97126 11646
rect 97092 10260 97126 10552
rect 97092 9166 97126 9458
rect 98150 13542 98184 13834
rect 98150 12448 98184 12740
rect 98150 11354 98184 11646
rect 98150 10260 98184 10552
rect 98150 9166 98184 9458
rect 99208 13542 99242 13834
rect 99208 12448 99242 12740
rect 99208 11354 99242 11646
rect 99208 10260 99242 10552
rect 99208 9166 99242 9458
rect 100266 13542 100300 13834
rect 100266 12448 100300 12740
rect 100266 11354 100300 11646
rect 100266 10260 100300 10552
rect 100266 9166 100300 9458
rect 100876 9760 101098 13456
rect 58352 6610 58386 6902
rect 58352 5516 58386 5808
rect 58352 4422 58386 4714
rect 58352 3328 58386 3620
rect 59410 7704 59444 7996
rect 59410 6610 59444 6902
rect 62118 7722 62152 8014
rect 63176 7722 63210 8014
rect 59410 5516 59444 5808
rect 59684 5340 59850 6714
rect 62118 6628 62152 6920
rect 63176 6628 63210 6920
rect 59410 4422 59444 4714
rect 59410 3328 59444 3620
rect 61486 5284 61580 6480
rect 62118 5534 62152 5826
rect 63176 5534 63210 5826
rect 62118 4440 62152 4732
rect 63176 4440 63210 4732
rect 62118 3346 62152 3638
rect 63176 3346 63210 3638
rect 64234 7722 64268 8014
rect 64234 6628 64268 6920
rect 64234 5534 64268 5826
rect 64234 4440 64268 4732
rect 64234 3346 64268 3638
rect 65292 7722 65326 8014
rect 65292 6628 65326 6920
rect 65292 5534 65326 5826
rect 65292 4440 65326 4732
rect 65292 3346 65326 3638
rect 66350 7722 66384 8014
rect 66350 6628 66384 6920
rect 66350 5534 66384 5826
rect 66350 4440 66384 4732
rect 66350 3346 66384 3638
rect 67408 7722 67442 8014
rect 67408 6628 67442 6920
rect 68590 7720 68624 8012
rect 69648 7720 69682 8012
rect 68590 6626 68624 6918
rect 69648 6626 69682 6918
rect 67408 5534 67442 5826
rect 67408 4440 67442 4732
rect 67408 3346 67442 3638
rect 67958 5282 68052 6478
rect 68590 5532 68624 5824
rect 69648 5532 69682 5824
rect 68590 4438 68624 4730
rect 69648 4438 69682 4730
rect 68590 3344 68624 3636
rect 69648 3344 69682 3636
rect 70706 7720 70740 8012
rect 70706 6626 70740 6918
rect 70706 5532 70740 5824
rect 70706 4438 70740 4730
rect 70706 3344 70740 3636
rect 71764 7720 71798 8012
rect 71764 6626 71798 6918
rect 71764 5532 71798 5824
rect 71764 4438 71798 4730
rect 71764 3344 71798 3636
rect 72822 7720 72856 8012
rect 72822 6626 72856 6918
rect 72822 5532 72856 5824
rect 72822 4438 72856 4730
rect 72822 3344 72856 3636
rect 73880 7720 73914 8012
rect 73880 6626 73914 6918
rect 75274 7694 75308 7986
rect 76332 7694 76366 7986
rect 75274 6600 75308 6892
rect 76332 6600 76366 6892
rect 73880 5532 73914 5824
rect 73880 4438 73914 4730
rect 73880 3344 73914 3636
rect 74642 5256 74736 6452
rect 39836 -1246 41558 -496
rect 59520 -682 60594 -184
rect 67080 -192 69254 840
rect 75274 5506 75308 5798
rect 76332 5506 76366 5798
rect 75274 4412 75308 4704
rect 76332 4412 76366 4704
rect 75274 3318 75308 3610
rect 76332 3318 76366 3610
rect 77390 7694 77424 7986
rect 77390 6600 77424 6892
rect 77390 5506 77424 5798
rect 77390 4412 77424 4704
rect 77390 3318 77424 3610
rect 78448 7694 78482 7986
rect 78448 6600 78482 6892
rect 78448 5506 78482 5798
rect 78448 4412 78482 4704
rect 78448 3318 78482 3610
rect 79506 7694 79540 7986
rect 79506 6600 79540 6892
rect 79506 5506 79540 5798
rect 79506 4412 79540 4704
rect 79506 3318 79540 3610
rect 80564 7694 80598 7986
rect 80564 6600 80598 6892
rect 81746 7692 81780 7984
rect 82804 7692 82838 7984
rect 81746 6598 81780 6890
rect 82804 6598 82838 6890
rect 80564 5506 80598 5798
rect 81114 5254 81208 6450
rect 81746 5504 81780 5796
rect 82804 5504 82838 5796
rect 80564 4412 80598 4704
rect 80564 3318 80598 3610
rect 81746 4410 81780 4702
rect 82804 4410 82838 4702
rect 81746 3316 81780 3608
rect 82804 3316 82838 3608
rect 83862 7692 83896 7984
rect 83862 6598 83896 6890
rect 83862 5504 83896 5796
rect 83862 4410 83896 4702
rect 83862 3316 83896 3608
rect 84920 7692 84954 7984
rect 84920 6598 84954 6890
rect 84920 5504 84954 5796
rect 84920 4410 84954 4702
rect 84920 3316 84954 3608
rect 85978 7692 86012 7984
rect 85978 6598 86012 6890
rect 85978 5504 86012 5796
rect 85978 4410 86012 4702
rect 85978 3316 86012 3608
rect 87036 7692 87070 7984
rect 87036 6598 87070 6890
rect 88508 7686 88542 7978
rect 89566 7686 89600 7978
rect 88508 6592 88542 6884
rect 89566 6592 89600 6884
rect 87036 5504 87070 5796
rect 87876 5248 87970 6444
rect 88508 5498 88542 5790
rect 89566 5498 89600 5790
rect 87036 4410 87070 4702
rect 87036 3316 87070 3608
rect 88508 4404 88542 4696
rect 89566 4404 89600 4696
rect 88508 3310 88542 3602
rect 89566 3310 89600 3602
rect 90624 7686 90658 7978
rect 90624 6592 90658 6884
rect 90624 5498 90658 5790
rect 90624 4404 90658 4696
rect 90624 3310 90658 3602
rect 91682 7686 91716 7978
rect 91682 6592 91716 6884
rect 91682 5498 91716 5790
rect 91682 4404 91716 4696
rect 91682 3310 91716 3602
rect 92740 7686 92774 7978
rect 92740 6592 92774 6884
rect 92740 5498 92774 5790
rect 92740 4404 92774 4696
rect 92740 3310 92774 3602
rect 93798 7686 93832 7978
rect 93798 6592 93832 6884
rect 94980 7684 95014 7976
rect 96038 7684 96072 7976
rect 94980 6590 95014 6882
rect 96038 6590 96072 6882
rect 93798 5498 93832 5790
rect 94348 5246 94442 6442
rect 94980 5496 95014 5788
rect 96038 5496 96072 5788
rect 93798 4404 93832 4696
rect 93798 3310 93832 3602
rect 94980 4402 95014 4694
rect 96038 4402 96072 4694
rect 94980 3308 95014 3600
rect 96038 3308 96072 3600
rect 97096 7684 97130 7976
rect 97096 6590 97130 6882
rect 97096 5496 97130 5788
rect 97096 4402 97130 4694
rect 97096 3308 97130 3600
rect 98154 7684 98188 7976
rect 98154 6590 98188 6882
rect 98154 5496 98188 5788
rect 98154 4402 98188 4694
rect 98154 3308 98188 3600
rect 99212 7684 99246 7976
rect 99212 6590 99246 6882
rect 99212 5496 99246 5788
rect 99212 4402 99246 4694
rect 99212 3308 99246 3600
rect 100270 7684 100304 7976
rect 100270 6590 100304 6882
rect 100270 5496 100304 5788
rect 100270 4402 100304 4694
rect 100270 3308 100304 3600
rect 100898 3594 101098 7268
rect 73674 -228 75848 804
<< metal1 >>
rect 58792 78708 94938 78714
rect 788 76048 94938 78708
rect 3778 69202 4576 76048
rect 42754 73680 45400 73768
rect 56220 73766 56604 76048
rect 58792 75912 94938 76048
rect 42754 73478 43052 73680
rect 45226 73478 45400 73680
rect 42754 73366 45400 73478
rect 46762 73678 49408 73766
rect 46762 73476 47060 73678
rect 49234 73476 49408 73678
rect 46762 73364 49408 73476
rect 50774 73678 53420 73766
rect 50774 73476 51072 73678
rect 53246 73476 53420 73678
rect 50774 73364 53420 73476
rect 54784 73678 57430 73766
rect 54784 73476 55082 73678
rect 57256 73476 57430 73678
rect 54784 73364 57430 73476
rect 42398 73228 42594 73234
rect 42398 73194 42410 73228
rect 42582 73194 42594 73228
rect 42398 73188 42594 73194
rect 43092 73228 43288 73234
rect 43092 73194 43104 73228
rect 43276 73194 43288 73228
rect 43092 73188 43288 73194
rect 43786 73228 43982 73234
rect 43786 73194 43798 73228
rect 43970 73194 43982 73228
rect 43786 73188 43982 73194
rect 44480 73228 44676 73234
rect 44480 73194 44492 73228
rect 44664 73194 44676 73228
rect 44480 73188 44676 73194
rect 45174 73228 45370 73234
rect 45174 73194 45186 73228
rect 45358 73194 45370 73228
rect 45174 73188 45370 73194
rect 46406 73226 46602 73232
rect 46406 73192 46418 73226
rect 46590 73192 46602 73226
rect 46406 73186 46602 73192
rect 47100 73226 47296 73232
rect 47100 73192 47112 73226
rect 47284 73192 47296 73226
rect 47100 73186 47296 73192
rect 47794 73226 47990 73232
rect 47794 73192 47806 73226
rect 47978 73192 47990 73226
rect 47794 73186 47990 73192
rect 48488 73226 48684 73232
rect 48488 73192 48500 73226
rect 48672 73192 48684 73226
rect 48488 73186 48684 73192
rect 49182 73226 49378 73232
rect 49182 73192 49194 73226
rect 49366 73192 49378 73226
rect 49182 73186 49378 73192
rect 50418 73226 50614 73232
rect 50418 73192 50430 73226
rect 50602 73192 50614 73226
rect 50418 73186 50614 73192
rect 51112 73226 51308 73232
rect 51112 73192 51124 73226
rect 51296 73192 51308 73226
rect 51112 73186 51308 73192
rect 51806 73226 52002 73232
rect 51806 73192 51818 73226
rect 51990 73192 52002 73226
rect 51806 73186 52002 73192
rect 52500 73226 52696 73232
rect 52500 73192 52512 73226
rect 52684 73192 52696 73226
rect 52500 73186 52696 73192
rect 53194 73226 53390 73232
rect 53194 73192 53206 73226
rect 53378 73192 53390 73226
rect 53194 73186 53390 73192
rect 54428 73226 54624 73232
rect 54428 73192 54440 73226
rect 54612 73192 54624 73226
rect 54428 73186 54624 73192
rect 55122 73226 55318 73232
rect 55122 73192 55134 73226
rect 55306 73192 55318 73226
rect 55122 73186 55318 73192
rect 55816 73226 56012 73232
rect 55816 73192 55828 73226
rect 56000 73192 56012 73226
rect 55816 73186 56012 73192
rect 56510 73226 56706 73232
rect 56510 73192 56522 73226
rect 56694 73192 56706 73226
rect 56510 73186 56706 73192
rect 57204 73226 57400 73232
rect 57204 73192 57216 73226
rect 57388 73192 57400 73226
rect 57204 73186 57400 73192
rect 70984 72980 71248 75912
rect 72564 74482 72908 74538
rect 72564 74380 72632 74482
rect 72838 74380 72908 74482
rect 72564 74328 72908 74380
rect 71332 74040 71378 74052
rect 71332 73868 71338 74040
rect 71372 73868 71378 74040
rect 71332 73856 71378 73868
rect 71990 74040 72036 74052
rect 71990 73868 71996 74040
rect 72030 73868 72036 74040
rect 71990 73856 72036 73868
rect 72648 74040 72694 74052
rect 72648 73868 72654 74040
rect 72688 73868 72694 74040
rect 73306 74040 73352 74052
rect 73306 73924 73312 74040
rect 72648 73856 72694 73868
rect 73240 73868 73312 73924
rect 73346 73924 73352 74040
rect 73964 74040 74010 74052
rect 73346 73868 73366 73924
rect 73240 73532 73366 73868
rect 73964 73868 73970 74040
rect 74004 73868 74010 74040
rect 73964 73856 74010 73868
rect 75196 74020 75242 74032
rect 75196 73848 75202 74020
rect 75236 73848 75242 74020
rect 75196 73836 75242 73848
rect 75854 74020 75900 74032
rect 75854 73848 75860 74020
rect 75894 73848 75900 74020
rect 75854 73836 75900 73848
rect 76512 74020 76558 74032
rect 76512 73848 76518 74020
rect 76552 73848 76558 74020
rect 77170 74020 77216 74032
rect 77170 73904 77176 74020
rect 76512 73836 76558 73848
rect 77104 73848 77176 73904
rect 77210 73904 77216 74020
rect 77770 74020 77930 75912
rect 80314 74572 80914 74608
rect 80314 74422 80464 74572
rect 80754 74422 80914 74572
rect 80314 74366 80914 74422
rect 77770 73944 77834 74020
rect 77210 73848 77230 73904
rect 73238 73500 73366 73532
rect 77104 73512 77230 73848
rect 77828 73848 77834 73944
rect 77868 73944 77930 74020
rect 79046 74034 79092 74046
rect 77868 73848 77874 73944
rect 79046 73862 79052 74034
rect 79086 73862 79092 74034
rect 79046 73850 79092 73862
rect 79704 74034 79750 74046
rect 79704 73862 79710 74034
rect 79744 73862 79750 74034
rect 79704 73850 79750 73862
rect 80362 74034 80408 74046
rect 80362 73862 80368 74034
rect 80402 73862 80408 74034
rect 81020 74034 81066 74046
rect 81020 73918 81026 74034
rect 80362 73850 80408 73862
rect 80954 73862 81026 73918
rect 81060 73918 81066 74034
rect 81678 74034 81724 74046
rect 81060 73862 81080 73918
rect 77828 73836 77874 73848
rect 80954 73526 81080 73862
rect 81678 73862 81684 74034
rect 81718 73862 81724 74034
rect 81678 73850 81724 73862
rect 73238 73466 73338 73500
rect 70984 72778 71066 72980
rect 42398 72570 42594 72576
rect 42398 72536 42410 72570
rect 42582 72536 42594 72570
rect 42398 72530 42594 72536
rect 43092 72570 43288 72576
rect 43092 72536 43104 72570
rect 43276 72536 43288 72570
rect 43092 72530 43288 72536
rect 43786 72570 43982 72576
rect 43786 72536 43798 72570
rect 43970 72536 43982 72570
rect 43786 72530 43982 72536
rect 44480 72570 44676 72576
rect 44480 72536 44492 72570
rect 44664 72536 44676 72570
rect 44480 72530 44676 72536
rect 45174 72570 45370 72576
rect 45174 72536 45186 72570
rect 45358 72536 45370 72570
rect 45174 72530 45370 72536
rect 46406 72568 46602 72574
rect 46406 72534 46418 72568
rect 46590 72534 46602 72568
rect 46406 72528 46602 72534
rect 47100 72568 47296 72574
rect 47100 72534 47112 72568
rect 47284 72534 47296 72568
rect 47100 72528 47296 72534
rect 47794 72568 47990 72574
rect 47794 72534 47806 72568
rect 47978 72534 47990 72568
rect 47794 72528 47990 72534
rect 48488 72568 48684 72574
rect 48488 72534 48500 72568
rect 48672 72534 48684 72568
rect 48488 72528 48684 72534
rect 49182 72568 49378 72574
rect 49182 72534 49194 72568
rect 49366 72534 49378 72568
rect 49182 72528 49378 72534
rect 50418 72568 50614 72574
rect 50418 72534 50430 72568
rect 50602 72534 50614 72568
rect 50418 72528 50614 72534
rect 51112 72568 51308 72574
rect 51112 72534 51124 72568
rect 51296 72534 51308 72568
rect 51112 72528 51308 72534
rect 51806 72568 52002 72574
rect 51806 72534 51818 72568
rect 51990 72534 52002 72568
rect 51806 72528 52002 72534
rect 52500 72568 52696 72574
rect 52500 72534 52512 72568
rect 52684 72534 52696 72568
rect 52500 72528 52696 72534
rect 53194 72568 53390 72574
rect 53194 72534 53206 72568
rect 53378 72534 53390 72568
rect 53194 72528 53390 72534
rect 54428 72568 54624 72574
rect 54428 72534 54440 72568
rect 54612 72534 54624 72568
rect 54428 72528 54624 72534
rect 55122 72568 55318 72574
rect 55122 72534 55134 72568
rect 55306 72534 55318 72568
rect 55122 72528 55318 72534
rect 55816 72568 56012 72574
rect 55816 72534 55828 72568
rect 56000 72534 56012 72568
rect 55816 72528 56012 72534
rect 56510 72568 56706 72574
rect 56510 72534 56522 72568
rect 56694 72534 56706 72568
rect 56510 72528 56706 72534
rect 57204 72568 57400 72574
rect 57204 72534 57216 72568
rect 57388 72534 57400 72568
rect 57204 72528 57400 72534
rect 42398 71912 42594 71918
rect 42398 71878 42410 71912
rect 42582 71878 42594 71912
rect 42398 71872 42594 71878
rect 43092 71912 43288 71918
rect 43092 71878 43104 71912
rect 43276 71878 43288 71912
rect 43092 71872 43288 71878
rect 43786 71912 43982 71918
rect 43786 71878 43798 71912
rect 43970 71878 43982 71912
rect 43786 71872 43982 71878
rect 44480 71912 44676 71918
rect 44480 71878 44492 71912
rect 44664 71878 44676 71912
rect 44480 71872 44676 71878
rect 45174 71912 45370 71918
rect 45174 71878 45186 71912
rect 45358 71878 45370 71912
rect 45174 71872 45370 71878
rect 46406 71910 46602 71916
rect 46406 71876 46418 71910
rect 46590 71876 46602 71910
rect 46406 71870 46602 71876
rect 47100 71910 47296 71916
rect 47100 71876 47112 71910
rect 47284 71876 47296 71910
rect 47100 71870 47296 71876
rect 47794 71910 47990 71916
rect 47794 71876 47806 71910
rect 47978 71876 47990 71910
rect 47794 71870 47990 71876
rect 48488 71910 48684 71916
rect 48488 71876 48500 71910
rect 48672 71876 48684 71910
rect 48488 71870 48684 71876
rect 49182 71910 49378 71916
rect 49182 71876 49194 71910
rect 49366 71876 49378 71910
rect 49182 71870 49378 71876
rect 50418 71910 50614 71916
rect 50418 71876 50430 71910
rect 50602 71876 50614 71910
rect 50418 71870 50614 71876
rect 51112 71910 51308 71916
rect 51112 71876 51124 71910
rect 51296 71876 51308 71910
rect 51112 71870 51308 71876
rect 51806 71910 52002 71916
rect 51806 71876 51818 71910
rect 51990 71876 52002 71910
rect 51806 71870 52002 71876
rect 52500 71910 52696 71916
rect 52500 71876 52512 71910
rect 52684 71876 52696 71910
rect 52500 71870 52696 71876
rect 53194 71910 53390 71916
rect 53194 71876 53206 71910
rect 53378 71876 53390 71910
rect 53194 71870 53390 71876
rect 54428 71910 54624 71916
rect 54428 71876 54440 71910
rect 54612 71876 54624 71910
rect 54428 71870 54624 71876
rect 55122 71910 55318 71916
rect 55122 71876 55134 71910
rect 55306 71876 55318 71910
rect 55122 71870 55318 71876
rect 55816 71910 56012 71916
rect 55816 71876 55828 71910
rect 56000 71876 56012 71910
rect 55816 71870 56012 71876
rect 56510 71910 56706 71916
rect 56510 71876 56522 71910
rect 56694 71876 56706 71910
rect 56510 71870 56706 71876
rect 57204 71910 57400 71916
rect 57204 71876 57216 71910
rect 57388 71876 57400 71910
rect 57204 71870 57400 71876
rect 42398 71254 42594 71260
rect 42398 71220 42410 71254
rect 42582 71220 42594 71254
rect 42398 71214 42594 71220
rect 43092 71254 43288 71260
rect 43092 71220 43104 71254
rect 43276 71220 43288 71254
rect 43092 71214 43288 71220
rect 43786 71254 43982 71260
rect 43786 71220 43798 71254
rect 43970 71220 43982 71254
rect 43786 71214 43982 71220
rect 44480 71254 44676 71260
rect 44480 71220 44492 71254
rect 44664 71220 44676 71254
rect 44480 71214 44676 71220
rect 45174 71254 45370 71260
rect 45174 71220 45186 71254
rect 45358 71220 45370 71254
rect 45174 71214 45370 71220
rect 46406 71252 46602 71258
rect 46406 71218 46418 71252
rect 46590 71218 46602 71252
rect 46406 71212 46602 71218
rect 47100 71252 47296 71258
rect 47100 71218 47112 71252
rect 47284 71218 47296 71252
rect 47100 71212 47296 71218
rect 47794 71252 47990 71258
rect 47794 71218 47806 71252
rect 47978 71218 47990 71252
rect 47794 71212 47990 71218
rect 48488 71252 48684 71258
rect 48488 71218 48500 71252
rect 48672 71218 48684 71252
rect 48488 71212 48684 71218
rect 49182 71252 49378 71258
rect 49182 71218 49194 71252
rect 49366 71218 49378 71252
rect 49182 71212 49378 71218
rect 50418 71252 50614 71258
rect 50418 71218 50430 71252
rect 50602 71218 50614 71252
rect 50418 71212 50614 71218
rect 51112 71252 51308 71258
rect 51112 71218 51124 71252
rect 51296 71218 51308 71252
rect 51112 71212 51308 71218
rect 51806 71252 52002 71258
rect 51806 71218 51818 71252
rect 51990 71218 52002 71252
rect 51806 71212 52002 71218
rect 52500 71252 52696 71258
rect 52500 71218 52512 71252
rect 52684 71218 52696 71252
rect 52500 71212 52696 71218
rect 53194 71252 53390 71258
rect 53194 71218 53206 71252
rect 53378 71218 53390 71252
rect 53194 71212 53390 71218
rect 54428 71252 54624 71258
rect 54428 71218 54440 71252
rect 54612 71218 54624 71252
rect 54428 71212 54624 71218
rect 55122 71252 55318 71258
rect 55122 71218 55134 71252
rect 55306 71218 55318 71252
rect 55122 71212 55318 71218
rect 55816 71252 56012 71258
rect 55816 71218 55828 71252
rect 56000 71218 56012 71252
rect 55816 71212 56012 71218
rect 56510 71252 56706 71258
rect 56510 71218 56522 71252
rect 56694 71218 56706 71252
rect 56510 71212 56706 71218
rect 57204 71252 57400 71258
rect 57204 71218 57216 71252
rect 57388 71218 57400 71252
rect 57204 71212 57400 71218
rect 42398 70596 42594 70602
rect 42398 70562 42410 70596
rect 42582 70562 42594 70596
rect 42398 70556 42594 70562
rect 43092 70596 43288 70602
rect 43092 70562 43104 70596
rect 43276 70562 43288 70596
rect 43092 70556 43288 70562
rect 43786 70596 43982 70602
rect 43786 70562 43798 70596
rect 43970 70562 43982 70596
rect 43786 70556 43982 70562
rect 44480 70596 44676 70602
rect 44480 70562 44492 70596
rect 44664 70562 44676 70596
rect 44480 70556 44676 70562
rect 45174 70596 45370 70602
rect 45174 70562 45186 70596
rect 45358 70562 45370 70596
rect 45174 70556 45370 70562
rect 46406 70594 46602 70600
rect 46406 70560 46418 70594
rect 46590 70560 46602 70594
rect 46406 70554 46602 70560
rect 47100 70594 47296 70600
rect 47100 70560 47112 70594
rect 47284 70560 47296 70594
rect 47100 70554 47296 70560
rect 47794 70594 47990 70600
rect 47794 70560 47806 70594
rect 47978 70560 47990 70594
rect 47794 70554 47990 70560
rect 48488 70594 48684 70600
rect 48488 70560 48500 70594
rect 48672 70560 48684 70594
rect 48488 70554 48684 70560
rect 49182 70594 49378 70600
rect 49182 70560 49194 70594
rect 49366 70560 49378 70594
rect 49182 70554 49378 70560
rect 50418 70594 50614 70600
rect 50418 70560 50430 70594
rect 50602 70560 50614 70594
rect 50418 70554 50614 70560
rect 51112 70594 51308 70600
rect 51112 70560 51124 70594
rect 51296 70560 51308 70594
rect 51112 70554 51308 70560
rect 51806 70594 52002 70600
rect 51806 70560 51818 70594
rect 51990 70560 52002 70594
rect 51806 70554 52002 70560
rect 52500 70594 52696 70600
rect 52500 70560 52512 70594
rect 52684 70560 52696 70594
rect 52500 70554 52696 70560
rect 53194 70594 53390 70600
rect 53194 70560 53206 70594
rect 53378 70560 53390 70594
rect 53194 70554 53390 70560
rect 54428 70594 54624 70600
rect 54428 70560 54440 70594
rect 54612 70560 54624 70594
rect 54428 70554 54624 70560
rect 55122 70594 55318 70600
rect 55122 70560 55134 70594
rect 55306 70560 55318 70594
rect 55122 70554 55318 70560
rect 55816 70594 56012 70600
rect 55816 70560 55828 70594
rect 56000 70560 56012 70594
rect 55816 70554 56012 70560
rect 56510 70594 56706 70600
rect 56510 70560 56522 70594
rect 56694 70560 56706 70594
rect 56510 70554 56706 70560
rect 57204 70594 57400 70600
rect 57204 70560 57216 70594
rect 57388 70560 57400 70594
rect 57204 70554 57400 70560
rect 71012 70412 71066 72778
rect 71150 72778 71248 72980
rect 71304 73126 71350 73138
rect 71304 72954 71310 73126
rect 71344 72954 71350 73126
rect 71304 72942 71350 72954
rect 71962 73126 72008 73138
rect 71962 72954 71968 73126
rect 72002 72954 72008 73126
rect 71962 72942 72008 72954
rect 72620 73126 72666 73138
rect 72620 72954 72626 73126
rect 72660 72954 72666 73126
rect 73240 73126 73338 73466
rect 77102 73480 77230 73512
rect 80952 73494 81080 73526
rect 77102 73446 77202 73480
rect 80952 73460 81052 73494
rect 73240 73072 73284 73126
rect 73266 73070 73284 73072
rect 72620 72942 72666 72954
rect 73278 72954 73284 73070
rect 73318 73070 73338 73126
rect 73936 73126 73982 73138
rect 73318 72954 73324 73070
rect 73278 72942 73324 72954
rect 73936 72954 73942 73126
rect 73976 72954 73982 73126
rect 75168 73106 75214 73118
rect 73936 72942 73982 72954
rect 74876 72960 75092 73106
rect 71150 70412 71228 72778
rect 71304 72432 71350 72444
rect 71304 72260 71310 72432
rect 71344 72260 71350 72432
rect 71304 72248 71350 72260
rect 71962 72432 72008 72444
rect 71962 72260 71968 72432
rect 72002 72260 72008 72432
rect 71962 72248 72008 72260
rect 72620 72432 72666 72444
rect 72620 72260 72626 72432
rect 72660 72260 72666 72432
rect 72620 72248 72666 72260
rect 73278 72432 73324 72444
rect 73278 72260 73284 72432
rect 73318 72260 73324 72432
rect 73278 72248 73324 72260
rect 73936 72432 73982 72444
rect 73936 72260 73942 72432
rect 73976 72260 73982 72432
rect 73936 72248 73982 72260
rect 71304 71738 71350 71750
rect 71304 71566 71310 71738
rect 71344 71566 71350 71738
rect 71304 71554 71350 71566
rect 71962 71738 72008 71750
rect 71962 71566 71968 71738
rect 72002 71566 72008 71738
rect 71962 71554 72008 71566
rect 72620 71738 72666 71750
rect 72620 71566 72626 71738
rect 72660 71566 72666 71738
rect 72620 71554 72666 71566
rect 73278 71738 73324 71750
rect 73278 71566 73284 71738
rect 73318 71566 73324 71738
rect 73278 71554 73324 71566
rect 73936 71738 73982 71750
rect 73936 71566 73942 71738
rect 73976 71566 73982 71738
rect 73936 71554 73982 71566
rect 71304 71044 71350 71056
rect 71304 70872 71310 71044
rect 71344 70872 71350 71044
rect 71304 70860 71350 70872
rect 71962 71044 72008 71056
rect 71962 70872 71968 71044
rect 72002 70872 72008 71044
rect 71962 70860 72008 70872
rect 72620 71044 72666 71056
rect 72620 70872 72626 71044
rect 72660 70872 72666 71044
rect 72620 70860 72666 70872
rect 73278 71044 73324 71056
rect 73278 70872 73284 71044
rect 73318 70872 73324 71044
rect 73278 70860 73324 70872
rect 73936 71044 73982 71056
rect 73936 70872 73942 71044
rect 73976 70872 73982 71044
rect 73936 70860 73982 70872
rect 71012 70266 71228 70412
rect 74876 70392 74930 72960
rect 75014 70392 75092 72960
rect 75168 72934 75174 73106
rect 75208 72934 75214 73106
rect 75168 72922 75214 72934
rect 75826 73106 75872 73118
rect 75826 72934 75832 73106
rect 75866 72934 75872 73106
rect 75826 72922 75872 72934
rect 76484 73106 76530 73118
rect 76484 72934 76490 73106
rect 76524 72934 76530 73106
rect 77104 73106 77202 73446
rect 79018 73120 79064 73132
rect 77104 73052 77148 73106
rect 77130 73050 77148 73052
rect 76484 72922 76530 72934
rect 77142 72934 77148 73050
rect 77182 73050 77202 73106
rect 77800 73106 77846 73118
rect 77182 72934 77188 73050
rect 77142 72922 77188 72934
rect 77800 72934 77806 73106
rect 77840 72934 77846 73106
rect 77800 72922 77846 72934
rect 78726 72974 78942 73120
rect 75168 72412 75214 72424
rect 75168 72240 75174 72412
rect 75208 72240 75214 72412
rect 75168 72228 75214 72240
rect 75826 72412 75872 72424
rect 75826 72240 75832 72412
rect 75866 72240 75872 72412
rect 75826 72228 75872 72240
rect 76484 72412 76530 72424
rect 76484 72240 76490 72412
rect 76524 72240 76530 72412
rect 76484 72228 76530 72240
rect 77142 72412 77188 72424
rect 77142 72240 77148 72412
rect 77182 72240 77188 72412
rect 77142 72228 77188 72240
rect 77800 72412 77846 72424
rect 77800 72240 77806 72412
rect 77840 72240 77846 72412
rect 77800 72228 77846 72240
rect 75168 71718 75214 71730
rect 75168 71546 75174 71718
rect 75208 71546 75214 71718
rect 75168 71534 75214 71546
rect 75826 71718 75872 71730
rect 75826 71546 75832 71718
rect 75866 71546 75872 71718
rect 75826 71534 75872 71546
rect 76484 71718 76530 71730
rect 76484 71546 76490 71718
rect 76524 71546 76530 71718
rect 76484 71534 76530 71546
rect 77142 71718 77188 71730
rect 77142 71546 77148 71718
rect 77182 71546 77188 71718
rect 77142 71534 77188 71546
rect 77800 71718 77846 71730
rect 77800 71546 77806 71718
rect 77840 71546 77846 71718
rect 77800 71534 77846 71546
rect 75168 71024 75214 71036
rect 75168 70852 75174 71024
rect 75208 70852 75214 71024
rect 75168 70840 75214 70852
rect 75826 71024 75872 71036
rect 75826 70852 75832 71024
rect 75866 70852 75872 71024
rect 75826 70840 75872 70852
rect 76484 71024 76530 71036
rect 76484 70852 76490 71024
rect 76524 70852 76530 71024
rect 76484 70840 76530 70852
rect 77142 71024 77188 71036
rect 77142 70852 77148 71024
rect 77182 70852 77188 71024
rect 77142 70840 77188 70852
rect 77800 71024 77846 71036
rect 77800 70852 77806 71024
rect 77840 70852 77846 71024
rect 77800 70840 77846 70852
rect 71304 70350 71350 70362
rect 71304 70178 71310 70350
rect 71344 70178 71350 70350
rect 71304 70166 71350 70178
rect 71962 70350 72008 70362
rect 71962 70178 71968 70350
rect 72002 70178 72008 70350
rect 71962 70166 72008 70178
rect 72620 70350 72666 70362
rect 72620 70178 72626 70350
rect 72660 70178 72666 70350
rect 73278 70350 73324 70362
rect 73278 70236 73284 70350
rect 72620 70166 72666 70178
rect 73262 70178 73284 70236
rect 73318 70236 73324 70350
rect 73936 70350 73982 70362
rect 73318 70178 73346 70236
rect 42398 69938 42594 69944
rect 42398 69904 42410 69938
rect 42582 69904 42594 69938
rect 42398 69898 42594 69904
rect 43092 69938 43288 69944
rect 43092 69904 43104 69938
rect 43276 69904 43288 69938
rect 43092 69898 43288 69904
rect 43786 69938 43982 69944
rect 43786 69904 43798 69938
rect 43970 69904 43982 69938
rect 43786 69898 43982 69904
rect 44480 69938 44676 69944
rect 44480 69904 44492 69938
rect 44664 69904 44676 69938
rect 44480 69898 44676 69904
rect 45174 69938 45370 69944
rect 45174 69904 45186 69938
rect 45358 69904 45370 69938
rect 45174 69898 45370 69904
rect 46406 69936 46602 69942
rect 46406 69902 46418 69936
rect 46590 69902 46602 69936
rect 46406 69896 46602 69902
rect 47100 69936 47296 69942
rect 47100 69902 47112 69936
rect 47284 69902 47296 69936
rect 47100 69896 47296 69902
rect 47794 69936 47990 69942
rect 47794 69902 47806 69936
rect 47978 69902 47990 69936
rect 47794 69896 47990 69902
rect 48488 69936 48684 69942
rect 48488 69902 48500 69936
rect 48672 69902 48684 69936
rect 48488 69896 48684 69902
rect 49182 69936 49378 69942
rect 49182 69902 49194 69936
rect 49366 69902 49378 69936
rect 49182 69896 49378 69902
rect 50418 69936 50614 69942
rect 50418 69902 50430 69936
rect 50602 69902 50614 69936
rect 50418 69896 50614 69902
rect 51112 69936 51308 69942
rect 51112 69902 51124 69936
rect 51296 69902 51308 69936
rect 51112 69896 51308 69902
rect 51806 69936 52002 69942
rect 51806 69902 51818 69936
rect 51990 69902 52002 69936
rect 51806 69896 52002 69902
rect 52500 69936 52696 69942
rect 52500 69902 52512 69936
rect 52684 69902 52696 69936
rect 52500 69896 52696 69902
rect 53194 69936 53390 69942
rect 53194 69902 53206 69936
rect 53378 69902 53390 69936
rect 53194 69896 53390 69902
rect 54428 69936 54624 69942
rect 54428 69902 54440 69936
rect 54612 69902 54624 69936
rect 54428 69896 54624 69902
rect 55122 69936 55318 69942
rect 55122 69902 55134 69936
rect 55306 69902 55318 69936
rect 55122 69896 55318 69902
rect 55816 69936 56012 69942
rect 55816 69902 55828 69936
rect 56000 69902 56012 69936
rect 55816 69896 56012 69902
rect 56510 69936 56706 69942
rect 56510 69902 56522 69936
rect 56694 69902 56706 69936
rect 56510 69896 56706 69902
rect 57204 69936 57400 69942
rect 57204 69902 57216 69936
rect 57388 69902 57400 69936
rect 57204 69896 57400 69902
rect 57692 69662 57870 69752
rect 42746 69482 45392 69570
rect 42746 69280 43044 69482
rect 45218 69280 45392 69482
rect 3778 68604 4600 69202
rect 42746 69168 45392 69280
rect 46740 69482 49386 69570
rect 46740 69280 47038 69482
rect 49212 69280 49386 69482
rect 46740 69168 49386 69280
rect 50762 69482 53408 69570
rect 50762 69280 51060 69482
rect 53234 69280 53408 69482
rect 50762 69168 53408 69280
rect 54784 69482 57430 69570
rect 54784 69280 55082 69482
rect 57256 69280 57430 69482
rect 57692 69482 57740 69662
rect 57844 69482 57870 69662
rect 57692 69408 57870 69482
rect 71300 69350 71346 69362
rect 54784 69168 57430 69280
rect 71008 69204 71224 69350
rect 42390 69030 42586 69036
rect 42390 68996 42402 69030
rect 42574 68996 42586 69030
rect 42390 68990 42586 68996
rect 43084 69030 43280 69036
rect 43084 68996 43096 69030
rect 43268 68996 43280 69030
rect 43084 68990 43280 68996
rect 43778 69030 43974 69036
rect 43778 68996 43790 69030
rect 43962 68996 43974 69030
rect 43778 68990 43974 68996
rect 44472 69030 44668 69036
rect 44472 68996 44484 69030
rect 44656 68996 44668 69030
rect 44472 68990 44668 68996
rect 45166 69030 45362 69036
rect 45166 68996 45178 69030
rect 45350 68996 45362 69030
rect 45166 68990 45362 68996
rect 46384 69030 46580 69036
rect 46384 68996 46396 69030
rect 46568 68996 46580 69030
rect 46384 68990 46580 68996
rect 47078 69030 47274 69036
rect 47078 68996 47090 69030
rect 47262 68996 47274 69030
rect 47078 68990 47274 68996
rect 47772 69030 47968 69036
rect 47772 68996 47784 69030
rect 47956 68996 47968 69030
rect 47772 68990 47968 68996
rect 48466 69030 48662 69036
rect 48466 68996 48478 69030
rect 48650 68996 48662 69030
rect 48466 68990 48662 68996
rect 49160 69030 49356 69036
rect 49160 68996 49172 69030
rect 49344 68996 49356 69030
rect 49160 68990 49356 68996
rect 50406 69030 50602 69036
rect 50406 68996 50418 69030
rect 50590 68996 50602 69030
rect 50406 68990 50602 68996
rect 51100 69030 51296 69036
rect 51100 68996 51112 69030
rect 51284 68996 51296 69030
rect 51100 68990 51296 68996
rect 51794 69030 51990 69036
rect 51794 68996 51806 69030
rect 51978 68996 51990 69030
rect 51794 68990 51990 68996
rect 52488 69030 52684 69036
rect 52488 68996 52500 69030
rect 52672 68996 52684 69030
rect 52488 68990 52684 68996
rect 53182 69030 53378 69036
rect 53182 68996 53194 69030
rect 53366 68996 53378 69030
rect 53182 68990 53378 68996
rect 54428 69030 54624 69036
rect 54428 68996 54440 69030
rect 54612 68996 54624 69030
rect 54428 68990 54624 68996
rect 55122 69030 55318 69036
rect 55122 68996 55134 69030
rect 55306 68996 55318 69030
rect 55122 68990 55318 68996
rect 55816 69030 56012 69036
rect 55816 68996 55828 69030
rect 56000 68996 56012 69030
rect 55816 68990 56012 68996
rect 56510 69030 56706 69036
rect 56510 68996 56522 69030
rect 56694 68996 56706 69030
rect 56510 68990 56706 68996
rect 57204 69030 57400 69036
rect 57204 68996 57216 69030
rect 57388 68996 57400 69030
rect 57204 68990 57400 68996
rect 972 65904 2604 65962
rect 3878 65958 4600 68604
rect 42390 68372 42586 68378
rect 42390 68338 42402 68372
rect 42574 68338 42586 68372
rect 42390 68332 42586 68338
rect 43084 68372 43280 68378
rect 43084 68338 43096 68372
rect 43268 68338 43280 68372
rect 43084 68332 43280 68338
rect 43778 68372 43974 68378
rect 43778 68338 43790 68372
rect 43962 68338 43974 68372
rect 43778 68332 43974 68338
rect 44472 68372 44668 68378
rect 44472 68338 44484 68372
rect 44656 68338 44668 68372
rect 44472 68332 44668 68338
rect 45166 68372 45362 68378
rect 45166 68338 45178 68372
rect 45350 68338 45362 68372
rect 45166 68332 45362 68338
rect 46384 68372 46580 68378
rect 46384 68338 46396 68372
rect 46568 68338 46580 68372
rect 46384 68332 46580 68338
rect 47078 68372 47274 68378
rect 47078 68338 47090 68372
rect 47262 68338 47274 68372
rect 47078 68332 47274 68338
rect 47772 68372 47968 68378
rect 47772 68338 47784 68372
rect 47956 68338 47968 68372
rect 47772 68332 47968 68338
rect 48466 68372 48662 68378
rect 48466 68338 48478 68372
rect 48650 68338 48662 68372
rect 48466 68332 48662 68338
rect 49160 68372 49356 68378
rect 49160 68338 49172 68372
rect 49344 68338 49356 68372
rect 49160 68332 49356 68338
rect 50406 68372 50602 68378
rect 50406 68338 50418 68372
rect 50590 68338 50602 68372
rect 50406 68332 50602 68338
rect 51100 68372 51296 68378
rect 51100 68338 51112 68372
rect 51284 68338 51296 68372
rect 51100 68332 51296 68338
rect 51794 68372 51990 68378
rect 51794 68338 51806 68372
rect 51978 68338 51990 68372
rect 51794 68332 51990 68338
rect 52488 68372 52684 68378
rect 52488 68338 52500 68372
rect 52672 68338 52684 68372
rect 52488 68332 52684 68338
rect 53182 68372 53378 68378
rect 53182 68338 53194 68372
rect 53366 68338 53378 68372
rect 53182 68332 53378 68338
rect 54428 68372 54624 68378
rect 54428 68338 54440 68372
rect 54612 68338 54624 68372
rect 54428 68332 54624 68338
rect 55122 68372 55318 68378
rect 55122 68338 55134 68372
rect 55306 68338 55318 68372
rect 55122 68332 55318 68338
rect 55816 68372 56012 68378
rect 55816 68338 55828 68372
rect 56000 68338 56012 68372
rect 55816 68332 56012 68338
rect 56510 68372 56706 68378
rect 56510 68338 56522 68372
rect 56694 68338 56706 68372
rect 56510 68332 56706 68338
rect 57204 68372 57400 68378
rect 57204 68338 57216 68372
rect 57388 68338 57400 68372
rect 57204 68332 57400 68338
rect 42390 67714 42586 67720
rect 42390 67680 42402 67714
rect 42574 67680 42586 67714
rect 42390 67674 42586 67680
rect 43084 67714 43280 67720
rect 43084 67680 43096 67714
rect 43268 67680 43280 67714
rect 43084 67674 43280 67680
rect 43778 67714 43974 67720
rect 43778 67680 43790 67714
rect 43962 67680 43974 67714
rect 43778 67674 43974 67680
rect 44472 67714 44668 67720
rect 44472 67680 44484 67714
rect 44656 67680 44668 67714
rect 44472 67674 44668 67680
rect 45166 67714 45362 67720
rect 45166 67680 45178 67714
rect 45350 67680 45362 67714
rect 45166 67674 45362 67680
rect 46384 67714 46580 67720
rect 46384 67680 46396 67714
rect 46568 67680 46580 67714
rect 46384 67674 46580 67680
rect 47078 67714 47274 67720
rect 47078 67680 47090 67714
rect 47262 67680 47274 67714
rect 47078 67674 47274 67680
rect 47772 67714 47968 67720
rect 47772 67680 47784 67714
rect 47956 67680 47968 67714
rect 47772 67674 47968 67680
rect 48466 67714 48662 67720
rect 48466 67680 48478 67714
rect 48650 67680 48662 67714
rect 48466 67674 48662 67680
rect 49160 67714 49356 67720
rect 49160 67680 49172 67714
rect 49344 67680 49356 67714
rect 49160 67674 49356 67680
rect 50406 67714 50602 67720
rect 50406 67680 50418 67714
rect 50590 67680 50602 67714
rect 50406 67674 50602 67680
rect 51100 67714 51296 67720
rect 51100 67680 51112 67714
rect 51284 67680 51296 67714
rect 51100 67674 51296 67680
rect 51794 67714 51990 67720
rect 51794 67680 51806 67714
rect 51978 67680 51990 67714
rect 51794 67674 51990 67680
rect 52488 67714 52684 67720
rect 52488 67680 52500 67714
rect 52672 67680 52684 67714
rect 52488 67674 52684 67680
rect 53182 67714 53378 67720
rect 53182 67680 53194 67714
rect 53366 67680 53378 67714
rect 53182 67674 53378 67680
rect 54428 67714 54624 67720
rect 54428 67680 54440 67714
rect 54612 67680 54624 67714
rect 54428 67674 54624 67680
rect 55122 67714 55318 67720
rect 55122 67680 55134 67714
rect 55306 67680 55318 67714
rect 55122 67674 55318 67680
rect 55816 67714 56012 67720
rect 55816 67680 55828 67714
rect 56000 67680 56012 67714
rect 55816 67674 56012 67680
rect 56510 67714 56706 67720
rect 56510 67680 56522 67714
rect 56694 67680 56706 67714
rect 56510 67674 56706 67680
rect 57204 67714 57400 67720
rect 57204 67680 57216 67714
rect 57388 67680 57400 67714
rect 57204 67674 57400 67680
rect 42390 67056 42586 67062
rect 42390 67022 42402 67056
rect 42574 67022 42586 67056
rect 42390 67016 42586 67022
rect 43084 67056 43280 67062
rect 43084 67022 43096 67056
rect 43268 67022 43280 67056
rect 43084 67016 43280 67022
rect 43778 67056 43974 67062
rect 43778 67022 43790 67056
rect 43962 67022 43974 67056
rect 43778 67016 43974 67022
rect 44472 67056 44668 67062
rect 44472 67022 44484 67056
rect 44656 67022 44668 67056
rect 44472 67016 44668 67022
rect 45166 67056 45362 67062
rect 45166 67022 45178 67056
rect 45350 67022 45362 67056
rect 45166 67016 45362 67022
rect 46384 67056 46580 67062
rect 46384 67022 46396 67056
rect 46568 67022 46580 67056
rect 46384 67016 46580 67022
rect 47078 67056 47274 67062
rect 47078 67022 47090 67056
rect 47262 67022 47274 67056
rect 47078 67016 47274 67022
rect 47772 67056 47968 67062
rect 47772 67022 47784 67056
rect 47956 67022 47968 67056
rect 47772 67016 47968 67022
rect 48466 67056 48662 67062
rect 48466 67022 48478 67056
rect 48650 67022 48662 67056
rect 48466 67016 48662 67022
rect 49160 67056 49356 67062
rect 49160 67022 49172 67056
rect 49344 67022 49356 67056
rect 49160 67016 49356 67022
rect 50406 67056 50602 67062
rect 50406 67022 50418 67056
rect 50590 67022 50602 67056
rect 50406 67016 50602 67022
rect 51100 67056 51296 67062
rect 51100 67022 51112 67056
rect 51284 67022 51296 67056
rect 51100 67016 51296 67022
rect 51794 67056 51990 67062
rect 51794 67022 51806 67056
rect 51978 67022 51990 67056
rect 51794 67016 51990 67022
rect 52488 67056 52684 67062
rect 52488 67022 52500 67056
rect 52672 67022 52684 67056
rect 52488 67016 52684 67022
rect 53182 67056 53378 67062
rect 53182 67022 53194 67056
rect 53366 67022 53378 67056
rect 53182 67016 53378 67022
rect 54428 67056 54624 67062
rect 54428 67022 54440 67056
rect 54612 67022 54624 67056
rect 54428 67016 54624 67022
rect 55122 67056 55318 67062
rect 55122 67022 55134 67056
rect 55306 67022 55318 67056
rect 55122 67016 55318 67022
rect 55816 67056 56012 67062
rect 55816 67022 55828 67056
rect 56000 67022 56012 67056
rect 55816 67016 56012 67022
rect 56510 67056 56706 67062
rect 56510 67022 56522 67056
rect 56694 67022 56706 67056
rect 56510 67016 56706 67022
rect 57204 67056 57400 67062
rect 57204 67022 57216 67056
rect 57388 67022 57400 67056
rect 57204 67016 57400 67022
rect 71008 66636 71062 69204
rect 71146 66636 71224 69204
rect 71300 69178 71306 69350
rect 71340 69178 71346 69350
rect 71300 69166 71346 69178
rect 71958 69350 72004 69362
rect 71958 69178 71964 69350
rect 71998 69178 72004 69350
rect 71958 69166 72004 69178
rect 72616 69350 72662 69362
rect 72616 69178 72622 69350
rect 72656 69178 72662 69350
rect 73262 69350 73346 70178
rect 73936 70178 73942 70350
rect 73976 70178 73982 70350
rect 74876 70246 75092 70392
rect 78726 70406 78780 72974
rect 78864 70406 78942 72974
rect 79018 72948 79024 73120
rect 79058 72948 79064 73120
rect 79018 72936 79064 72948
rect 79676 73120 79722 73132
rect 79676 72948 79682 73120
rect 79716 72948 79722 73120
rect 79676 72936 79722 72948
rect 80334 73120 80380 73132
rect 80334 72948 80340 73120
rect 80374 72948 80380 73120
rect 80954 73120 81052 73460
rect 80954 73066 80998 73120
rect 80980 73064 80998 73066
rect 80334 72936 80380 72948
rect 80992 72948 80998 73064
rect 81032 73064 81052 73120
rect 81650 73120 81696 73132
rect 81032 72948 81038 73064
rect 80992 72936 81038 72948
rect 81650 72948 81656 73120
rect 81690 72948 81696 73120
rect 81650 72936 81696 72948
rect 79018 72426 79064 72438
rect 79018 72254 79024 72426
rect 79058 72254 79064 72426
rect 79018 72242 79064 72254
rect 79676 72426 79722 72438
rect 79676 72254 79682 72426
rect 79716 72254 79722 72426
rect 79676 72242 79722 72254
rect 80334 72426 80380 72438
rect 80334 72254 80340 72426
rect 80374 72254 80380 72426
rect 80334 72242 80380 72254
rect 80992 72426 81038 72438
rect 80992 72254 80998 72426
rect 81032 72254 81038 72426
rect 80992 72242 81038 72254
rect 81650 72426 81696 72438
rect 81650 72254 81656 72426
rect 81690 72254 81696 72426
rect 81650 72242 81696 72254
rect 79018 71732 79064 71744
rect 79018 71560 79024 71732
rect 79058 71560 79064 71732
rect 79018 71548 79064 71560
rect 79676 71732 79722 71744
rect 79676 71560 79682 71732
rect 79716 71560 79722 71732
rect 79676 71548 79722 71560
rect 80334 71732 80380 71744
rect 80334 71560 80340 71732
rect 80374 71560 80380 71732
rect 80334 71548 80380 71560
rect 80992 71732 81038 71744
rect 80992 71560 80998 71732
rect 81032 71560 81038 71732
rect 80992 71548 81038 71560
rect 81650 71732 81696 71744
rect 81650 71560 81656 71732
rect 81690 71560 81696 71732
rect 81650 71548 81696 71560
rect 79018 71038 79064 71050
rect 79018 70866 79024 71038
rect 79058 70866 79064 71038
rect 79018 70854 79064 70866
rect 79676 71038 79722 71050
rect 79676 70866 79682 71038
rect 79716 70866 79722 71038
rect 79676 70854 79722 70866
rect 80334 71038 80380 71050
rect 80334 70866 80340 71038
rect 80374 70866 80380 71038
rect 80334 70854 80380 70866
rect 80992 71038 81038 71050
rect 80992 70866 80998 71038
rect 81032 70866 81038 71038
rect 80992 70854 81038 70866
rect 81650 71038 81696 71050
rect 81650 70866 81656 71038
rect 81690 70866 81696 71038
rect 81650 70854 81696 70866
rect 75168 70330 75214 70342
rect 73936 70166 73982 70178
rect 75168 70158 75174 70330
rect 75208 70158 75214 70330
rect 75168 70146 75214 70158
rect 75826 70330 75872 70342
rect 75826 70158 75832 70330
rect 75866 70158 75872 70330
rect 75826 70146 75872 70158
rect 76484 70330 76530 70342
rect 76484 70158 76490 70330
rect 76524 70158 76530 70330
rect 77142 70330 77188 70342
rect 77142 70216 77148 70330
rect 76484 70146 76530 70158
rect 77126 70158 77148 70216
rect 77182 70216 77188 70330
rect 77800 70330 77846 70342
rect 77182 70158 77210 70216
rect 73262 69290 73280 69350
rect 72616 69166 72662 69178
rect 73274 69178 73280 69290
rect 73314 69290 73346 69350
rect 73932 69350 73978 69362
rect 73314 69178 73320 69290
rect 73274 69166 73320 69178
rect 73932 69178 73938 69350
rect 73972 69178 73978 69350
rect 75164 69330 75210 69342
rect 73932 69166 73978 69178
rect 74872 69184 75088 69330
rect 71300 68656 71346 68668
rect 71300 68484 71306 68656
rect 71340 68484 71346 68656
rect 71300 68472 71346 68484
rect 71958 68656 72004 68668
rect 71958 68484 71964 68656
rect 71998 68484 72004 68656
rect 71958 68472 72004 68484
rect 72616 68656 72662 68668
rect 72616 68484 72622 68656
rect 72656 68484 72662 68656
rect 72616 68472 72662 68484
rect 73274 68656 73320 68668
rect 73274 68484 73280 68656
rect 73314 68484 73320 68656
rect 73274 68472 73320 68484
rect 73932 68656 73978 68668
rect 73932 68484 73938 68656
rect 73972 68484 73978 68656
rect 73932 68472 73978 68484
rect 71300 67962 71346 67974
rect 71300 67790 71306 67962
rect 71340 67790 71346 67962
rect 71300 67778 71346 67790
rect 71958 67962 72004 67974
rect 71958 67790 71964 67962
rect 71998 67790 72004 67962
rect 71958 67778 72004 67790
rect 72616 67962 72662 67974
rect 72616 67790 72622 67962
rect 72656 67790 72662 67962
rect 72616 67778 72662 67790
rect 73274 67962 73320 67974
rect 73274 67790 73280 67962
rect 73314 67790 73320 67962
rect 73274 67778 73320 67790
rect 73932 67962 73978 67974
rect 73932 67790 73938 67962
rect 73972 67790 73978 67962
rect 73932 67778 73978 67790
rect 71300 67268 71346 67280
rect 71300 67096 71306 67268
rect 71340 67096 71346 67268
rect 71300 67084 71346 67096
rect 71958 67268 72004 67280
rect 71958 67096 71964 67268
rect 71998 67096 72004 67268
rect 71958 67084 72004 67096
rect 72616 67268 72662 67280
rect 72616 67096 72622 67268
rect 72656 67096 72662 67268
rect 72616 67084 72662 67096
rect 73274 67268 73320 67280
rect 73274 67096 73280 67268
rect 73314 67096 73320 67268
rect 73274 67084 73320 67096
rect 73932 67268 73978 67280
rect 73932 67096 73938 67268
rect 73972 67096 73978 67268
rect 73932 67084 73978 67096
rect 71008 66490 71224 66636
rect 74872 66616 74926 69184
rect 75010 66616 75088 69184
rect 75164 69158 75170 69330
rect 75204 69158 75210 69330
rect 75164 69146 75210 69158
rect 75822 69330 75868 69342
rect 75822 69158 75828 69330
rect 75862 69158 75868 69330
rect 75822 69146 75868 69158
rect 76480 69330 76526 69342
rect 76480 69158 76486 69330
rect 76520 69158 76526 69330
rect 77126 69330 77210 70158
rect 77800 70158 77806 70330
rect 77840 70158 77846 70330
rect 78726 70260 78942 70406
rect 79018 70344 79064 70356
rect 79018 70172 79024 70344
rect 79058 70172 79064 70344
rect 79018 70160 79064 70172
rect 79676 70344 79722 70356
rect 79676 70172 79682 70344
rect 79716 70172 79722 70344
rect 79676 70160 79722 70172
rect 80334 70344 80380 70356
rect 80334 70172 80340 70344
rect 80374 70172 80380 70344
rect 80992 70344 81038 70356
rect 80992 70230 80998 70344
rect 80334 70160 80380 70172
rect 80976 70172 80998 70230
rect 81032 70230 81038 70344
rect 81650 70344 81696 70356
rect 81032 70172 81060 70230
rect 77800 70146 77846 70158
rect 79014 69344 79060 69356
rect 77126 69270 77144 69330
rect 76480 69146 76526 69158
rect 77138 69158 77144 69270
rect 77178 69270 77210 69330
rect 77796 69330 77842 69342
rect 77178 69158 77184 69270
rect 77138 69146 77184 69158
rect 77796 69158 77802 69330
rect 77836 69158 77842 69330
rect 77796 69146 77842 69158
rect 78722 69198 78938 69344
rect 75164 68636 75210 68648
rect 75164 68464 75170 68636
rect 75204 68464 75210 68636
rect 75164 68452 75210 68464
rect 75822 68636 75868 68648
rect 75822 68464 75828 68636
rect 75862 68464 75868 68636
rect 75822 68452 75868 68464
rect 76480 68636 76526 68648
rect 76480 68464 76486 68636
rect 76520 68464 76526 68636
rect 76480 68452 76526 68464
rect 77138 68636 77184 68648
rect 77138 68464 77144 68636
rect 77178 68464 77184 68636
rect 77138 68452 77184 68464
rect 77796 68636 77842 68648
rect 77796 68464 77802 68636
rect 77836 68464 77842 68636
rect 77796 68452 77842 68464
rect 75164 67942 75210 67954
rect 75164 67770 75170 67942
rect 75204 67770 75210 67942
rect 75164 67758 75210 67770
rect 75822 67942 75868 67954
rect 75822 67770 75828 67942
rect 75862 67770 75868 67942
rect 75822 67758 75868 67770
rect 76480 67942 76526 67954
rect 76480 67770 76486 67942
rect 76520 67770 76526 67942
rect 76480 67758 76526 67770
rect 77138 67942 77184 67954
rect 77138 67770 77144 67942
rect 77178 67770 77184 67942
rect 77138 67758 77184 67770
rect 77796 67942 77842 67954
rect 77796 67770 77802 67942
rect 77836 67770 77842 67942
rect 77796 67758 77842 67770
rect 75164 67248 75210 67260
rect 75164 67076 75170 67248
rect 75204 67076 75210 67248
rect 75164 67064 75210 67076
rect 75822 67248 75868 67260
rect 75822 67076 75828 67248
rect 75862 67076 75868 67248
rect 75822 67064 75868 67076
rect 76480 67248 76526 67260
rect 76480 67076 76486 67248
rect 76520 67076 76526 67248
rect 76480 67064 76526 67076
rect 77138 67248 77184 67260
rect 77138 67076 77144 67248
rect 77178 67076 77184 67248
rect 77138 67064 77184 67076
rect 77796 67248 77842 67260
rect 77796 67076 77802 67248
rect 77836 67076 77842 67248
rect 77796 67064 77842 67076
rect 71300 66574 71346 66586
rect 42390 66398 42586 66404
rect 42390 66364 42402 66398
rect 42574 66364 42586 66398
rect 42390 66358 42586 66364
rect 43084 66398 43280 66404
rect 43084 66364 43096 66398
rect 43268 66364 43280 66398
rect 43084 66358 43280 66364
rect 43778 66398 43974 66404
rect 43778 66364 43790 66398
rect 43962 66364 43974 66398
rect 43778 66358 43974 66364
rect 44472 66398 44668 66404
rect 44472 66364 44484 66398
rect 44656 66364 44668 66398
rect 44472 66358 44668 66364
rect 45166 66398 45362 66404
rect 45166 66364 45178 66398
rect 45350 66364 45362 66398
rect 45166 66358 45362 66364
rect 46384 66398 46580 66404
rect 46384 66364 46396 66398
rect 46568 66364 46580 66398
rect 46384 66358 46580 66364
rect 47078 66398 47274 66404
rect 47078 66364 47090 66398
rect 47262 66364 47274 66398
rect 47078 66358 47274 66364
rect 47772 66398 47968 66404
rect 47772 66364 47784 66398
rect 47956 66364 47968 66398
rect 47772 66358 47968 66364
rect 48466 66398 48662 66404
rect 48466 66364 48478 66398
rect 48650 66364 48662 66398
rect 48466 66358 48662 66364
rect 49160 66398 49356 66404
rect 49160 66364 49172 66398
rect 49344 66364 49356 66398
rect 49160 66358 49356 66364
rect 50406 66398 50602 66404
rect 50406 66364 50418 66398
rect 50590 66364 50602 66398
rect 50406 66358 50602 66364
rect 51100 66398 51296 66404
rect 51100 66364 51112 66398
rect 51284 66364 51296 66398
rect 51100 66358 51296 66364
rect 51794 66398 51990 66404
rect 51794 66364 51806 66398
rect 51978 66364 51990 66398
rect 51794 66358 51990 66364
rect 52488 66398 52684 66404
rect 52488 66364 52500 66398
rect 52672 66364 52684 66398
rect 52488 66358 52684 66364
rect 53182 66398 53378 66404
rect 53182 66364 53194 66398
rect 53366 66364 53378 66398
rect 53182 66358 53378 66364
rect 54428 66398 54624 66404
rect 54428 66364 54440 66398
rect 54612 66364 54624 66398
rect 54428 66358 54624 66364
rect 55122 66398 55318 66404
rect 55122 66364 55134 66398
rect 55306 66364 55318 66398
rect 55122 66358 55318 66364
rect 55816 66398 56012 66404
rect 55816 66364 55828 66398
rect 56000 66364 56012 66398
rect 55816 66358 56012 66364
rect 56510 66398 56706 66404
rect 56510 66364 56522 66398
rect 56694 66364 56706 66398
rect 56510 66358 56706 66364
rect 57204 66398 57400 66404
rect 57204 66364 57216 66398
rect 57388 66364 57400 66398
rect 71300 66402 71306 66574
rect 71340 66402 71346 66574
rect 71300 66390 71346 66402
rect 71958 66574 72004 66586
rect 71958 66402 71964 66574
rect 71998 66402 72004 66574
rect 71958 66390 72004 66402
rect 72616 66574 72662 66586
rect 72616 66402 72622 66574
rect 72656 66402 72662 66574
rect 73274 66574 73320 66586
rect 73274 66476 73280 66574
rect 72616 66390 72662 66402
rect 73238 66402 73280 66476
rect 73314 66476 73320 66574
rect 73932 66574 73978 66586
rect 73314 66402 73362 66476
rect 57204 66358 57400 66364
rect 972 65834 1086 65904
rect 2490 65834 2604 65904
rect 972 65758 2604 65834
rect 3640 65900 5272 65958
rect 3640 65830 3754 65900
rect 5158 65830 5272 65900
rect 3640 65754 5272 65830
rect 6314 65906 7946 65964
rect 6314 65836 6428 65906
rect 7832 65836 7946 65906
rect 6314 65760 7946 65836
rect 8960 65906 10592 65964
rect 8960 65836 9074 65906
rect 10478 65836 10592 65906
rect 8960 65760 10592 65836
rect 11614 65900 13246 65958
rect 11614 65830 11728 65900
rect 13132 65830 13246 65900
rect 11614 65754 13246 65830
rect 14268 65906 15900 65964
rect 14268 65836 14382 65906
rect 15786 65836 15900 65906
rect 14268 65760 15900 65836
rect 16894 65910 18526 65968
rect 16894 65840 17008 65910
rect 18412 65840 18526 65910
rect 16894 65764 18526 65840
rect 19392 65924 20628 65994
rect 19392 65816 19562 65924
rect 20520 65816 20628 65924
rect 19392 65724 20628 65816
rect 19560 65620 19756 65626
rect 19560 65586 19572 65620
rect 19744 65586 19756 65620
rect 954 65570 1150 65576
rect 954 65536 966 65570
rect 1138 65536 1150 65570
rect 954 65530 1150 65536
rect 1648 65570 1844 65576
rect 1648 65536 1660 65570
rect 1832 65536 1844 65570
rect 1648 65530 1844 65536
rect 2342 65570 2538 65576
rect 6296 65572 6492 65578
rect 2342 65536 2354 65570
rect 2526 65536 2538 65570
rect 2342 65530 2538 65536
rect 3622 65566 3818 65572
rect 3622 65532 3634 65566
rect 3806 65532 3818 65566
rect 3622 65526 3818 65532
rect 4316 65566 4512 65572
rect 4316 65532 4328 65566
rect 4500 65532 4512 65566
rect 4316 65526 4512 65532
rect 5010 65566 5206 65572
rect 5010 65532 5022 65566
rect 5194 65532 5206 65566
rect 6296 65538 6308 65572
rect 6480 65538 6492 65572
rect 6296 65532 6492 65538
rect 6990 65572 7186 65578
rect 6990 65538 7002 65572
rect 7174 65538 7186 65572
rect 6990 65532 7186 65538
rect 7684 65572 7880 65578
rect 7684 65538 7696 65572
rect 7868 65538 7880 65572
rect 7684 65532 7880 65538
rect 8942 65572 9138 65578
rect 8942 65538 8954 65572
rect 9126 65538 9138 65572
rect 8942 65532 9138 65538
rect 9636 65572 9832 65578
rect 9636 65538 9648 65572
rect 9820 65538 9832 65572
rect 9636 65532 9832 65538
rect 10330 65572 10526 65578
rect 14250 65572 14446 65578
rect 10330 65538 10342 65572
rect 10514 65538 10526 65572
rect 10330 65532 10526 65538
rect 11596 65566 11792 65572
rect 11596 65532 11608 65566
rect 11780 65532 11792 65566
rect 5010 65526 5206 65532
rect 11596 65526 11792 65532
rect 12290 65566 12486 65572
rect 12290 65532 12302 65566
rect 12474 65532 12486 65566
rect 12290 65526 12486 65532
rect 12984 65566 13180 65572
rect 12984 65532 12996 65566
rect 13168 65532 13180 65566
rect 14250 65538 14262 65572
rect 14434 65538 14446 65572
rect 14250 65532 14446 65538
rect 14944 65572 15140 65578
rect 14944 65538 14956 65572
rect 15128 65538 15140 65572
rect 14944 65532 15140 65538
rect 15638 65572 15834 65578
rect 15638 65538 15650 65572
rect 15822 65538 15834 65572
rect 15638 65532 15834 65538
rect 16876 65576 17072 65582
rect 16876 65542 16888 65576
rect 17060 65542 17072 65576
rect 16876 65536 17072 65542
rect 17570 65576 17766 65582
rect 17570 65542 17582 65576
rect 17754 65542 17766 65576
rect 17570 65536 17766 65542
rect 18264 65576 18460 65582
rect 19560 65580 19756 65586
rect 20254 65620 20450 65626
rect 20254 65586 20266 65620
rect 20438 65586 20450 65620
rect 20254 65580 20450 65586
rect 18264 65542 18276 65576
rect 18448 65542 18460 65576
rect 18264 65536 18460 65542
rect 12984 65526 13180 65532
rect 38838 65126 38848 65882
rect 39974 65126 39984 65882
rect 42390 65740 42586 65746
rect 42390 65706 42402 65740
rect 42574 65706 42586 65740
rect 42390 65700 42586 65706
rect 43084 65740 43280 65746
rect 43084 65706 43096 65740
rect 43268 65706 43280 65740
rect 43084 65700 43280 65706
rect 43778 65740 43974 65746
rect 43778 65706 43790 65740
rect 43962 65706 43974 65740
rect 43778 65700 43974 65706
rect 44472 65740 44668 65746
rect 44472 65706 44484 65740
rect 44656 65706 44668 65740
rect 44472 65700 44668 65706
rect 45166 65740 45362 65746
rect 45166 65706 45178 65740
rect 45350 65706 45362 65740
rect 45166 65700 45362 65706
rect 46384 65740 46580 65746
rect 46384 65706 46396 65740
rect 46568 65706 46580 65740
rect 46384 65700 46580 65706
rect 47078 65740 47274 65746
rect 47078 65706 47090 65740
rect 47262 65706 47274 65740
rect 47078 65700 47274 65706
rect 47772 65740 47968 65746
rect 47772 65706 47784 65740
rect 47956 65706 47968 65740
rect 47772 65700 47968 65706
rect 48466 65740 48662 65746
rect 48466 65706 48478 65740
rect 48650 65706 48662 65740
rect 48466 65700 48662 65706
rect 49160 65740 49356 65746
rect 49160 65706 49172 65740
rect 49344 65706 49356 65740
rect 49160 65700 49356 65706
rect 50406 65740 50602 65746
rect 50406 65706 50418 65740
rect 50590 65706 50602 65740
rect 50406 65700 50602 65706
rect 51100 65740 51296 65746
rect 51100 65706 51112 65740
rect 51284 65706 51296 65740
rect 51100 65700 51296 65706
rect 51794 65740 51990 65746
rect 51794 65706 51806 65740
rect 51978 65706 51990 65740
rect 51794 65700 51990 65706
rect 52488 65740 52684 65746
rect 52488 65706 52500 65740
rect 52672 65706 52684 65740
rect 52488 65700 52684 65706
rect 53182 65740 53378 65746
rect 53182 65706 53194 65740
rect 53366 65706 53378 65740
rect 53182 65700 53378 65706
rect 54428 65740 54624 65746
rect 54428 65706 54440 65740
rect 54612 65706 54624 65740
rect 54428 65700 54624 65706
rect 55122 65740 55318 65746
rect 55122 65706 55134 65740
rect 55306 65706 55318 65740
rect 55122 65700 55318 65706
rect 55816 65740 56012 65746
rect 55816 65706 55828 65740
rect 56000 65706 56012 65740
rect 55816 65700 56012 65706
rect 56510 65740 56706 65746
rect 56510 65706 56522 65740
rect 56694 65706 56706 65740
rect 56510 65700 56706 65706
rect 57204 65740 57400 65746
rect 57204 65706 57216 65740
rect 57388 65706 57400 65740
rect 57204 65700 57400 65706
rect 71300 65580 71346 65592
rect 71008 65434 71224 65580
rect 19560 64962 19756 64968
rect 19560 64928 19572 64962
rect 19744 64928 19756 64962
rect 954 64912 1150 64918
rect 954 64878 966 64912
rect 1138 64878 1150 64912
rect 954 64872 1150 64878
rect 1648 64912 1844 64918
rect 1648 64878 1660 64912
rect 1832 64878 1844 64912
rect 1648 64872 1844 64878
rect 2342 64912 2538 64918
rect 6296 64914 6492 64920
rect 2342 64878 2354 64912
rect 2526 64878 2538 64912
rect 2342 64872 2538 64878
rect 3622 64908 3818 64914
rect 3622 64874 3634 64908
rect 3806 64874 3818 64908
rect 3622 64868 3818 64874
rect 4316 64908 4512 64914
rect 4316 64874 4328 64908
rect 4500 64874 4512 64908
rect 4316 64868 4512 64874
rect 5010 64908 5206 64914
rect 5010 64874 5022 64908
rect 5194 64874 5206 64908
rect 6296 64880 6308 64914
rect 6480 64880 6492 64914
rect 6296 64874 6492 64880
rect 6990 64914 7186 64920
rect 6990 64880 7002 64914
rect 7174 64880 7186 64914
rect 6990 64874 7186 64880
rect 7684 64914 7880 64920
rect 7684 64880 7696 64914
rect 7868 64880 7880 64914
rect 7684 64874 7880 64880
rect 8942 64914 9138 64920
rect 8942 64880 8954 64914
rect 9126 64880 9138 64914
rect 8942 64874 9138 64880
rect 9636 64914 9832 64920
rect 9636 64880 9648 64914
rect 9820 64880 9832 64914
rect 9636 64874 9832 64880
rect 10330 64914 10526 64920
rect 14250 64914 14446 64920
rect 10330 64880 10342 64914
rect 10514 64880 10526 64914
rect 10330 64874 10526 64880
rect 11596 64908 11792 64914
rect 11596 64874 11608 64908
rect 11780 64874 11792 64908
rect 5010 64868 5206 64874
rect 11596 64868 11792 64874
rect 12290 64908 12486 64914
rect 12290 64874 12302 64908
rect 12474 64874 12486 64908
rect 12290 64868 12486 64874
rect 12984 64908 13180 64914
rect 12984 64874 12996 64908
rect 13168 64874 13180 64908
rect 14250 64880 14262 64914
rect 14434 64880 14446 64914
rect 14250 64874 14446 64880
rect 14944 64914 15140 64920
rect 14944 64880 14956 64914
rect 15128 64880 15140 64914
rect 14944 64874 15140 64880
rect 15638 64914 15834 64920
rect 15638 64880 15650 64914
rect 15822 64880 15834 64914
rect 15638 64874 15834 64880
rect 16876 64918 17072 64924
rect 16876 64884 16888 64918
rect 17060 64884 17072 64918
rect 16876 64878 17072 64884
rect 17570 64918 17766 64924
rect 17570 64884 17582 64918
rect 17754 64884 17766 64918
rect 17570 64878 17766 64884
rect 18264 64918 18460 64924
rect 19560 64922 19756 64928
rect 20254 64962 20450 64968
rect 20254 64928 20266 64962
rect 20438 64928 20450 64962
rect 20254 64922 20450 64928
rect 18264 64884 18276 64918
rect 18448 64884 18460 64918
rect 18264 64878 18460 64884
rect 12984 64868 13180 64874
rect 19560 64304 19756 64310
rect 19560 64270 19572 64304
rect 19744 64270 19756 64304
rect 954 64254 1150 64260
rect 954 64220 966 64254
rect 1138 64220 1150 64254
rect 954 64214 1150 64220
rect 1648 64254 1844 64260
rect 1648 64220 1660 64254
rect 1832 64220 1844 64254
rect 1648 64214 1844 64220
rect 2342 64254 2538 64260
rect 6296 64256 6492 64262
rect 2342 64220 2354 64254
rect 2526 64220 2538 64254
rect 2342 64214 2538 64220
rect 3622 64250 3818 64256
rect 3622 64216 3634 64250
rect 3806 64216 3818 64250
rect 3622 64210 3818 64216
rect 4316 64250 4512 64256
rect 4316 64216 4328 64250
rect 4500 64216 4512 64250
rect 4316 64210 4512 64216
rect 5010 64250 5206 64256
rect 5010 64216 5022 64250
rect 5194 64216 5206 64250
rect 6296 64222 6308 64256
rect 6480 64222 6492 64256
rect 6296 64216 6492 64222
rect 6990 64256 7186 64262
rect 6990 64222 7002 64256
rect 7174 64222 7186 64256
rect 6990 64216 7186 64222
rect 7684 64256 7880 64262
rect 7684 64222 7696 64256
rect 7868 64222 7880 64256
rect 7684 64216 7880 64222
rect 8942 64256 9138 64262
rect 8942 64222 8954 64256
rect 9126 64222 9138 64256
rect 8942 64216 9138 64222
rect 9636 64256 9832 64262
rect 9636 64222 9648 64256
rect 9820 64222 9832 64256
rect 9636 64216 9832 64222
rect 10330 64256 10526 64262
rect 14250 64256 14446 64262
rect 10330 64222 10342 64256
rect 10514 64222 10526 64256
rect 10330 64216 10526 64222
rect 11596 64250 11792 64256
rect 11596 64216 11608 64250
rect 11780 64216 11792 64250
rect 5010 64210 5206 64216
rect 11596 64210 11792 64216
rect 12290 64250 12486 64256
rect 12290 64216 12302 64250
rect 12474 64216 12486 64250
rect 12290 64210 12486 64216
rect 12984 64250 13180 64256
rect 12984 64216 12996 64250
rect 13168 64216 13180 64250
rect 14250 64222 14262 64256
rect 14434 64222 14446 64256
rect 14250 64216 14446 64222
rect 14944 64256 15140 64262
rect 14944 64222 14956 64256
rect 15128 64222 15140 64256
rect 14944 64216 15140 64222
rect 15638 64256 15834 64262
rect 15638 64222 15650 64256
rect 15822 64222 15834 64256
rect 15638 64216 15834 64222
rect 16876 64260 17072 64266
rect 16876 64226 16888 64260
rect 17060 64226 17072 64260
rect 16876 64220 17072 64226
rect 17570 64260 17766 64266
rect 17570 64226 17582 64260
rect 17754 64226 17766 64260
rect 17570 64220 17766 64226
rect 18264 64260 18460 64266
rect 19560 64264 19756 64270
rect 20254 64304 20450 64310
rect 20254 64270 20266 64304
rect 20438 64270 20450 64304
rect 20254 64264 20450 64270
rect 39286 64292 39472 65126
rect 42734 65008 45380 65096
rect 42734 64806 43032 65008
rect 45206 64806 45380 65008
rect 42734 64694 45380 64806
rect 46742 65006 49388 65094
rect 46742 64804 47040 65006
rect 49214 64804 49388 65006
rect 46742 64692 49388 64804
rect 50754 65006 53400 65094
rect 50754 64804 51052 65006
rect 53226 64804 53400 65006
rect 50754 64692 53400 64804
rect 54764 65006 57410 65094
rect 54764 64804 55062 65006
rect 57236 64804 57410 65006
rect 54764 64692 57410 64804
rect 42378 64556 42574 64562
rect 42378 64522 42390 64556
rect 42562 64522 42574 64556
rect 42378 64516 42574 64522
rect 43072 64556 43268 64562
rect 43072 64522 43084 64556
rect 43256 64522 43268 64556
rect 43072 64516 43268 64522
rect 43766 64556 43962 64562
rect 43766 64522 43778 64556
rect 43950 64522 43962 64556
rect 43766 64516 43962 64522
rect 44460 64556 44656 64562
rect 44460 64522 44472 64556
rect 44644 64522 44656 64556
rect 44460 64516 44656 64522
rect 45154 64556 45350 64562
rect 45154 64522 45166 64556
rect 45338 64522 45350 64556
rect 45154 64516 45350 64522
rect 46386 64554 46582 64560
rect 46386 64520 46398 64554
rect 46570 64520 46582 64554
rect 46386 64514 46582 64520
rect 47080 64554 47276 64560
rect 47080 64520 47092 64554
rect 47264 64520 47276 64554
rect 47080 64514 47276 64520
rect 47774 64554 47970 64560
rect 47774 64520 47786 64554
rect 47958 64520 47970 64554
rect 47774 64514 47970 64520
rect 48468 64554 48664 64560
rect 48468 64520 48480 64554
rect 48652 64520 48664 64554
rect 48468 64514 48664 64520
rect 49162 64554 49358 64560
rect 49162 64520 49174 64554
rect 49346 64520 49358 64554
rect 49162 64514 49358 64520
rect 50398 64554 50594 64560
rect 50398 64520 50410 64554
rect 50582 64520 50594 64554
rect 50398 64514 50594 64520
rect 51092 64554 51288 64560
rect 51092 64520 51104 64554
rect 51276 64520 51288 64554
rect 51092 64514 51288 64520
rect 51786 64554 51982 64560
rect 51786 64520 51798 64554
rect 51970 64520 51982 64554
rect 51786 64514 51982 64520
rect 52480 64554 52676 64560
rect 52480 64520 52492 64554
rect 52664 64520 52676 64554
rect 52480 64514 52676 64520
rect 53174 64554 53370 64560
rect 53174 64520 53186 64554
rect 53358 64520 53370 64554
rect 53174 64514 53370 64520
rect 54408 64554 54604 64560
rect 54408 64520 54420 64554
rect 54592 64520 54604 64554
rect 54408 64514 54604 64520
rect 55102 64554 55298 64560
rect 55102 64520 55114 64554
rect 55286 64520 55298 64554
rect 55102 64514 55298 64520
rect 55796 64554 55992 64560
rect 55796 64520 55808 64554
rect 55980 64520 55992 64554
rect 55796 64514 55992 64520
rect 56490 64554 56686 64560
rect 56490 64520 56502 64554
rect 56674 64520 56686 64554
rect 56490 64514 56686 64520
rect 57184 64554 57380 64560
rect 57184 64520 57196 64554
rect 57368 64520 57380 64554
rect 57184 64514 57380 64520
rect 41772 64304 42106 64372
rect 41772 64292 41840 64304
rect 18264 64226 18276 64260
rect 18448 64226 18460 64260
rect 18264 64220 18460 64226
rect 12984 64210 13180 64216
rect 39286 64162 41840 64292
rect 20692 64112 20810 64144
rect 20692 64074 20732 64112
rect 20782 64074 20810 64112
rect 41772 64136 41840 64162
rect 42022 64136 42106 64304
rect 41772 64076 42106 64136
rect 20692 64032 20810 64074
rect 42378 63898 42574 63904
rect 42378 63864 42390 63898
rect 42562 63864 42574 63898
rect 42378 63858 42574 63864
rect 43072 63898 43268 63904
rect 43072 63864 43084 63898
rect 43256 63864 43268 63898
rect 43072 63858 43268 63864
rect 43766 63898 43962 63904
rect 43766 63864 43778 63898
rect 43950 63864 43962 63898
rect 43766 63858 43962 63864
rect 44460 63898 44656 63904
rect 44460 63864 44472 63898
rect 44644 63864 44656 63898
rect 44460 63858 44656 63864
rect 45154 63898 45350 63904
rect 45154 63864 45166 63898
rect 45338 63864 45350 63898
rect 45154 63858 45350 63864
rect 46386 63896 46582 63902
rect 46386 63862 46398 63896
rect 46570 63862 46582 63896
rect 46386 63856 46582 63862
rect 47080 63896 47276 63902
rect 47080 63862 47092 63896
rect 47264 63862 47276 63896
rect 47080 63856 47276 63862
rect 47774 63896 47970 63902
rect 47774 63862 47786 63896
rect 47958 63862 47970 63896
rect 47774 63856 47970 63862
rect 48468 63896 48664 63902
rect 48468 63862 48480 63896
rect 48652 63862 48664 63896
rect 48468 63856 48664 63862
rect 49162 63896 49358 63902
rect 49162 63862 49174 63896
rect 49346 63862 49358 63896
rect 49162 63856 49358 63862
rect 50398 63896 50594 63902
rect 50398 63862 50410 63896
rect 50582 63862 50594 63896
rect 50398 63856 50594 63862
rect 51092 63896 51288 63902
rect 51092 63862 51104 63896
rect 51276 63862 51288 63896
rect 51092 63856 51288 63862
rect 51786 63896 51982 63902
rect 51786 63862 51798 63896
rect 51970 63862 51982 63896
rect 51786 63856 51982 63862
rect 52480 63896 52676 63902
rect 52480 63862 52492 63896
rect 52664 63862 52676 63896
rect 52480 63856 52676 63862
rect 53174 63896 53370 63902
rect 53174 63862 53186 63896
rect 53358 63862 53370 63896
rect 53174 63856 53370 63862
rect 54408 63896 54604 63902
rect 54408 63862 54420 63896
rect 54592 63862 54604 63896
rect 54408 63856 54604 63862
rect 55102 63896 55298 63902
rect 55102 63862 55114 63896
rect 55286 63862 55298 63896
rect 55102 63856 55298 63862
rect 55796 63896 55992 63902
rect 55796 63862 55808 63896
rect 55980 63862 55992 63896
rect 55796 63856 55992 63862
rect 56490 63896 56686 63902
rect 56490 63862 56502 63896
rect 56674 63862 56686 63896
rect 56490 63856 56686 63862
rect 57184 63896 57380 63902
rect 57184 63862 57196 63896
rect 57368 63862 57380 63896
rect 57184 63856 57380 63862
rect 19560 63646 19756 63652
rect 19560 63612 19572 63646
rect 19744 63612 19756 63646
rect 954 63596 1150 63602
rect 954 63562 966 63596
rect 1138 63562 1150 63596
rect 954 63556 1150 63562
rect 1648 63596 1844 63602
rect 1648 63562 1660 63596
rect 1832 63562 1844 63596
rect 1648 63556 1844 63562
rect 2342 63596 2538 63602
rect 6296 63598 6492 63604
rect 2342 63562 2354 63596
rect 2526 63562 2538 63596
rect 2342 63556 2538 63562
rect 3622 63592 3818 63598
rect 3622 63558 3634 63592
rect 3806 63558 3818 63592
rect 3622 63552 3818 63558
rect 4316 63592 4512 63598
rect 4316 63558 4328 63592
rect 4500 63558 4512 63592
rect 4316 63552 4512 63558
rect 5010 63592 5206 63598
rect 5010 63558 5022 63592
rect 5194 63558 5206 63592
rect 6296 63564 6308 63598
rect 6480 63564 6492 63598
rect 6296 63558 6492 63564
rect 6990 63598 7186 63604
rect 6990 63564 7002 63598
rect 7174 63564 7186 63598
rect 6990 63558 7186 63564
rect 7684 63598 7880 63604
rect 7684 63564 7696 63598
rect 7868 63564 7880 63598
rect 7684 63558 7880 63564
rect 8942 63598 9138 63604
rect 8942 63564 8954 63598
rect 9126 63564 9138 63598
rect 8942 63558 9138 63564
rect 9636 63598 9832 63604
rect 9636 63564 9648 63598
rect 9820 63564 9832 63598
rect 9636 63558 9832 63564
rect 10330 63598 10526 63604
rect 14250 63598 14446 63604
rect 10330 63564 10342 63598
rect 10514 63564 10526 63598
rect 10330 63558 10526 63564
rect 11596 63592 11792 63598
rect 11596 63558 11608 63592
rect 11780 63558 11792 63592
rect 5010 63552 5206 63558
rect 11596 63552 11792 63558
rect 12290 63592 12486 63598
rect 12290 63558 12302 63592
rect 12474 63558 12486 63592
rect 12290 63552 12486 63558
rect 12984 63592 13180 63598
rect 12984 63558 12996 63592
rect 13168 63558 13180 63592
rect 14250 63564 14262 63598
rect 14434 63564 14446 63598
rect 14250 63558 14446 63564
rect 14944 63598 15140 63604
rect 14944 63564 14956 63598
rect 15128 63564 15140 63598
rect 14944 63558 15140 63564
rect 15638 63598 15834 63604
rect 15638 63564 15650 63598
rect 15822 63564 15834 63598
rect 15638 63558 15834 63564
rect 16876 63602 17072 63608
rect 16876 63568 16888 63602
rect 17060 63568 17072 63602
rect 16876 63562 17072 63568
rect 17570 63602 17766 63608
rect 17570 63568 17582 63602
rect 17754 63568 17766 63602
rect 17570 63562 17766 63568
rect 18264 63602 18460 63608
rect 19560 63606 19756 63612
rect 20254 63646 20450 63652
rect 20254 63612 20266 63646
rect 20438 63612 20450 63646
rect 20254 63606 20450 63612
rect 18264 63568 18276 63602
rect 18448 63568 18460 63602
rect 18264 63562 18460 63568
rect 12984 63552 13180 63558
rect 42378 63240 42574 63246
rect 42378 63206 42390 63240
rect 42562 63206 42574 63240
rect 42378 63200 42574 63206
rect 43072 63240 43268 63246
rect 43072 63206 43084 63240
rect 43256 63206 43268 63240
rect 43072 63200 43268 63206
rect 43766 63240 43962 63246
rect 43766 63206 43778 63240
rect 43950 63206 43962 63240
rect 43766 63200 43962 63206
rect 44460 63240 44656 63246
rect 44460 63206 44472 63240
rect 44644 63206 44656 63240
rect 44460 63200 44656 63206
rect 45154 63240 45350 63246
rect 45154 63206 45166 63240
rect 45338 63206 45350 63240
rect 45154 63200 45350 63206
rect 46386 63238 46582 63244
rect 46386 63204 46398 63238
rect 46570 63204 46582 63238
rect 46386 63198 46582 63204
rect 47080 63238 47276 63244
rect 47080 63204 47092 63238
rect 47264 63204 47276 63238
rect 47080 63198 47276 63204
rect 47774 63238 47970 63244
rect 47774 63204 47786 63238
rect 47958 63204 47970 63238
rect 47774 63198 47970 63204
rect 48468 63238 48664 63244
rect 48468 63204 48480 63238
rect 48652 63204 48664 63238
rect 48468 63198 48664 63204
rect 49162 63238 49358 63244
rect 49162 63204 49174 63238
rect 49346 63204 49358 63238
rect 49162 63198 49358 63204
rect 50398 63238 50594 63244
rect 50398 63204 50410 63238
rect 50582 63204 50594 63238
rect 50398 63198 50594 63204
rect 51092 63238 51288 63244
rect 51092 63204 51104 63238
rect 51276 63204 51288 63238
rect 51092 63198 51288 63204
rect 51786 63238 51982 63244
rect 51786 63204 51798 63238
rect 51970 63204 51982 63238
rect 51786 63198 51982 63204
rect 52480 63238 52676 63244
rect 52480 63204 52492 63238
rect 52664 63204 52676 63238
rect 52480 63198 52676 63204
rect 53174 63238 53370 63244
rect 53174 63204 53186 63238
rect 53358 63204 53370 63238
rect 53174 63198 53370 63204
rect 54408 63238 54604 63244
rect 54408 63204 54420 63238
rect 54592 63204 54604 63238
rect 54408 63198 54604 63204
rect 55102 63238 55298 63244
rect 55102 63204 55114 63238
rect 55286 63204 55298 63238
rect 55102 63198 55298 63204
rect 55796 63238 55992 63244
rect 55796 63204 55808 63238
rect 55980 63204 55992 63238
rect 55796 63198 55992 63204
rect 56490 63238 56686 63244
rect 56490 63204 56502 63238
rect 56674 63204 56686 63238
rect 56490 63198 56686 63204
rect 57184 63238 57380 63244
rect 57184 63204 57196 63238
rect 57368 63204 57380 63238
rect 57184 63198 57380 63204
rect 19560 62988 19756 62994
rect 19560 62954 19572 62988
rect 19744 62954 19756 62988
rect 954 62938 1150 62944
rect 954 62904 966 62938
rect 1138 62904 1150 62938
rect 954 62898 1150 62904
rect 1648 62938 1844 62944
rect 1648 62904 1660 62938
rect 1832 62904 1844 62938
rect 1648 62898 1844 62904
rect 2342 62938 2538 62944
rect 6296 62940 6492 62946
rect 2342 62904 2354 62938
rect 2526 62904 2538 62938
rect 2342 62898 2538 62904
rect 3622 62934 3818 62940
rect 3622 62900 3634 62934
rect 3806 62900 3818 62934
rect 3622 62894 3818 62900
rect 4316 62934 4512 62940
rect 4316 62900 4328 62934
rect 4500 62900 4512 62934
rect 4316 62894 4512 62900
rect 5010 62934 5206 62940
rect 5010 62900 5022 62934
rect 5194 62900 5206 62934
rect 6296 62906 6308 62940
rect 6480 62906 6492 62940
rect 6296 62900 6492 62906
rect 6990 62940 7186 62946
rect 6990 62906 7002 62940
rect 7174 62906 7186 62940
rect 6990 62900 7186 62906
rect 7684 62940 7880 62946
rect 7684 62906 7696 62940
rect 7868 62906 7880 62940
rect 7684 62900 7880 62906
rect 8942 62940 9138 62946
rect 8942 62906 8954 62940
rect 9126 62906 9138 62940
rect 8942 62900 9138 62906
rect 9636 62940 9832 62946
rect 9636 62906 9648 62940
rect 9820 62906 9832 62940
rect 9636 62900 9832 62906
rect 10330 62940 10526 62946
rect 14250 62940 14446 62946
rect 10330 62906 10342 62940
rect 10514 62906 10526 62940
rect 10330 62900 10526 62906
rect 11596 62934 11792 62940
rect 11596 62900 11608 62934
rect 11780 62900 11792 62934
rect 5010 62894 5206 62900
rect 11596 62894 11792 62900
rect 12290 62934 12486 62940
rect 12290 62900 12302 62934
rect 12474 62900 12486 62934
rect 12290 62894 12486 62900
rect 12984 62934 13180 62940
rect 12984 62900 12996 62934
rect 13168 62900 13180 62934
rect 14250 62906 14262 62940
rect 14434 62906 14446 62940
rect 14250 62900 14446 62906
rect 14944 62940 15140 62946
rect 14944 62906 14956 62940
rect 15128 62906 15140 62940
rect 14944 62900 15140 62906
rect 15638 62940 15834 62946
rect 15638 62906 15650 62940
rect 15822 62906 15834 62940
rect 15638 62900 15834 62906
rect 16876 62944 17072 62950
rect 16876 62910 16888 62944
rect 17060 62910 17072 62944
rect 16876 62904 17072 62910
rect 17570 62944 17766 62950
rect 17570 62910 17582 62944
rect 17754 62910 17766 62944
rect 17570 62904 17766 62910
rect 18264 62944 18460 62950
rect 19560 62948 19756 62954
rect 20254 62988 20450 62994
rect 20254 62954 20266 62988
rect 20438 62954 20450 62988
rect 20254 62948 20450 62954
rect 18264 62910 18276 62944
rect 18448 62910 18460 62944
rect 18264 62904 18460 62910
rect 12984 62894 13180 62900
rect 71008 62866 71062 65434
rect 71146 62866 71224 65434
rect 71300 65408 71306 65580
rect 71340 65408 71346 65580
rect 71300 65396 71346 65408
rect 71958 65580 72004 65592
rect 71958 65408 71964 65580
rect 71998 65408 72004 65580
rect 71958 65396 72004 65408
rect 72616 65580 72662 65592
rect 72616 65408 72622 65580
rect 72656 65408 72662 65580
rect 73238 65580 73362 66402
rect 73932 66402 73938 66574
rect 73972 66402 73978 66574
rect 74872 66470 75088 66616
rect 78722 66630 78776 69198
rect 78860 66630 78938 69198
rect 79014 69172 79020 69344
rect 79054 69172 79060 69344
rect 79014 69160 79060 69172
rect 79672 69344 79718 69356
rect 79672 69172 79678 69344
rect 79712 69172 79718 69344
rect 79672 69160 79718 69172
rect 80330 69344 80376 69356
rect 80330 69172 80336 69344
rect 80370 69172 80376 69344
rect 80976 69344 81060 70172
rect 81650 70172 81656 70344
rect 81690 70172 81696 70344
rect 81650 70160 81696 70172
rect 80976 69284 80994 69344
rect 80330 69160 80376 69172
rect 80988 69172 80994 69284
rect 81028 69284 81060 69344
rect 81646 69344 81692 69356
rect 81028 69172 81034 69284
rect 80988 69160 81034 69172
rect 81646 69172 81652 69344
rect 81686 69172 81692 69344
rect 81646 69160 81692 69172
rect 79014 68650 79060 68662
rect 79014 68478 79020 68650
rect 79054 68478 79060 68650
rect 79014 68466 79060 68478
rect 79672 68650 79718 68662
rect 79672 68478 79678 68650
rect 79712 68478 79718 68650
rect 79672 68466 79718 68478
rect 80330 68650 80376 68662
rect 80330 68478 80336 68650
rect 80370 68478 80376 68650
rect 80330 68466 80376 68478
rect 80988 68650 81034 68662
rect 80988 68478 80994 68650
rect 81028 68478 81034 68650
rect 80988 68466 81034 68478
rect 81646 68650 81692 68662
rect 81646 68478 81652 68650
rect 81686 68478 81692 68650
rect 81646 68466 81692 68478
rect 79014 67956 79060 67968
rect 79014 67784 79020 67956
rect 79054 67784 79060 67956
rect 79014 67772 79060 67784
rect 79672 67956 79718 67968
rect 79672 67784 79678 67956
rect 79712 67784 79718 67956
rect 79672 67772 79718 67784
rect 80330 67956 80376 67968
rect 80330 67784 80336 67956
rect 80370 67784 80376 67956
rect 80330 67772 80376 67784
rect 80988 67956 81034 67968
rect 80988 67784 80994 67956
rect 81028 67784 81034 67956
rect 80988 67772 81034 67784
rect 81646 67956 81692 67968
rect 81646 67784 81652 67956
rect 81686 67784 81692 67956
rect 81646 67772 81692 67784
rect 79014 67262 79060 67274
rect 79014 67090 79020 67262
rect 79054 67090 79060 67262
rect 79014 67078 79060 67090
rect 79672 67262 79718 67274
rect 79672 67090 79678 67262
rect 79712 67090 79718 67262
rect 79672 67078 79718 67090
rect 80330 67262 80376 67274
rect 80330 67090 80336 67262
rect 80370 67090 80376 67262
rect 80330 67078 80376 67090
rect 80988 67262 81034 67274
rect 80988 67090 80994 67262
rect 81028 67090 81034 67262
rect 80988 67078 81034 67090
rect 81646 67262 81692 67274
rect 81646 67090 81652 67262
rect 81686 67090 81692 67262
rect 81646 67078 81692 67090
rect 75164 66554 75210 66566
rect 73932 66390 73978 66402
rect 75164 66382 75170 66554
rect 75204 66382 75210 66554
rect 75164 66370 75210 66382
rect 75822 66554 75868 66566
rect 75822 66382 75828 66554
rect 75862 66382 75868 66554
rect 75822 66370 75868 66382
rect 76480 66554 76526 66566
rect 76480 66382 76486 66554
rect 76520 66382 76526 66554
rect 77138 66554 77184 66566
rect 77138 66456 77144 66554
rect 76480 66370 76526 66382
rect 77102 66382 77144 66456
rect 77178 66456 77184 66554
rect 77796 66554 77842 66566
rect 77178 66382 77226 66456
rect 73238 65478 73280 65580
rect 72616 65396 72662 65408
rect 73274 65408 73280 65478
rect 73314 65478 73362 65580
rect 73932 65580 73978 65592
rect 73314 65408 73320 65478
rect 73274 65396 73320 65408
rect 73932 65408 73938 65580
rect 73972 65408 73978 65580
rect 75164 65560 75210 65572
rect 73932 65396 73978 65408
rect 74872 65414 75088 65560
rect 71300 64886 71346 64898
rect 71300 64714 71306 64886
rect 71340 64714 71346 64886
rect 71300 64702 71346 64714
rect 71958 64886 72004 64898
rect 71958 64714 71964 64886
rect 71998 64714 72004 64886
rect 71958 64702 72004 64714
rect 72616 64886 72662 64898
rect 72616 64714 72622 64886
rect 72656 64714 72662 64886
rect 72616 64702 72662 64714
rect 73274 64886 73320 64898
rect 73274 64714 73280 64886
rect 73314 64714 73320 64886
rect 73274 64702 73320 64714
rect 73932 64886 73978 64898
rect 73932 64714 73938 64886
rect 73972 64714 73978 64886
rect 73932 64702 73978 64714
rect 71300 64192 71346 64204
rect 71300 64020 71306 64192
rect 71340 64020 71346 64192
rect 71300 64008 71346 64020
rect 71958 64192 72004 64204
rect 71958 64020 71964 64192
rect 71998 64020 72004 64192
rect 71958 64008 72004 64020
rect 72616 64192 72662 64204
rect 72616 64020 72622 64192
rect 72656 64020 72662 64192
rect 72616 64008 72662 64020
rect 73274 64192 73320 64204
rect 73274 64020 73280 64192
rect 73314 64020 73320 64192
rect 73274 64008 73320 64020
rect 73932 64192 73978 64204
rect 73932 64020 73938 64192
rect 73972 64020 73978 64192
rect 73932 64008 73978 64020
rect 71300 63498 71346 63510
rect 71300 63326 71306 63498
rect 71340 63326 71346 63498
rect 71300 63314 71346 63326
rect 71958 63498 72004 63510
rect 71958 63326 71964 63498
rect 71998 63326 72004 63498
rect 71958 63314 72004 63326
rect 72616 63498 72662 63510
rect 72616 63326 72622 63498
rect 72656 63326 72662 63498
rect 72616 63314 72662 63326
rect 73274 63498 73320 63510
rect 73274 63326 73280 63498
rect 73314 63326 73320 63498
rect 73274 63314 73320 63326
rect 73932 63498 73978 63510
rect 73932 63326 73938 63498
rect 73972 63326 73978 63498
rect 73932 63314 73978 63326
rect 71008 62720 71224 62866
rect 74872 62846 74926 65414
rect 75010 62846 75088 65414
rect 75164 65388 75170 65560
rect 75204 65388 75210 65560
rect 75164 65376 75210 65388
rect 75822 65560 75868 65572
rect 75822 65388 75828 65560
rect 75862 65388 75868 65560
rect 75822 65376 75868 65388
rect 76480 65560 76526 65572
rect 76480 65388 76486 65560
rect 76520 65388 76526 65560
rect 77102 65560 77226 66382
rect 77796 66382 77802 66554
rect 77836 66382 77842 66554
rect 78722 66484 78938 66630
rect 79014 66568 79060 66580
rect 79014 66396 79020 66568
rect 79054 66396 79060 66568
rect 79014 66384 79060 66396
rect 79672 66568 79718 66580
rect 79672 66396 79678 66568
rect 79712 66396 79718 66568
rect 79672 66384 79718 66396
rect 80330 66568 80376 66580
rect 80330 66396 80336 66568
rect 80370 66396 80376 66568
rect 80988 66568 81034 66580
rect 80988 66470 80994 66568
rect 80330 66384 80376 66396
rect 80952 66396 80994 66470
rect 81028 66470 81034 66568
rect 81646 66568 81692 66580
rect 81028 66396 81076 66470
rect 77796 66370 77842 66382
rect 79014 65574 79060 65586
rect 77102 65458 77144 65560
rect 76480 65376 76526 65388
rect 77138 65388 77144 65458
rect 77178 65458 77226 65560
rect 77796 65560 77842 65572
rect 77178 65388 77184 65458
rect 77138 65376 77184 65388
rect 77796 65388 77802 65560
rect 77836 65388 77842 65560
rect 77796 65376 77842 65388
rect 78722 65428 78938 65574
rect 75164 64866 75210 64878
rect 75164 64694 75170 64866
rect 75204 64694 75210 64866
rect 75164 64682 75210 64694
rect 75822 64866 75868 64878
rect 75822 64694 75828 64866
rect 75862 64694 75868 64866
rect 75822 64682 75868 64694
rect 76480 64866 76526 64878
rect 76480 64694 76486 64866
rect 76520 64694 76526 64866
rect 76480 64682 76526 64694
rect 77138 64866 77184 64878
rect 77138 64694 77144 64866
rect 77178 64694 77184 64866
rect 77138 64682 77184 64694
rect 77796 64866 77842 64878
rect 77796 64694 77802 64866
rect 77836 64694 77842 64866
rect 77796 64682 77842 64694
rect 75164 64172 75210 64184
rect 75164 64000 75170 64172
rect 75204 64000 75210 64172
rect 75164 63988 75210 64000
rect 75822 64172 75868 64184
rect 75822 64000 75828 64172
rect 75862 64000 75868 64172
rect 75822 63988 75868 64000
rect 76480 64172 76526 64184
rect 76480 64000 76486 64172
rect 76520 64000 76526 64172
rect 76480 63988 76526 64000
rect 77138 64172 77184 64184
rect 77138 64000 77144 64172
rect 77178 64000 77184 64172
rect 77138 63988 77184 64000
rect 77796 64172 77842 64184
rect 77796 64000 77802 64172
rect 77836 64000 77842 64172
rect 77796 63988 77842 64000
rect 75164 63478 75210 63490
rect 75164 63306 75170 63478
rect 75204 63306 75210 63478
rect 75164 63294 75210 63306
rect 75822 63478 75868 63490
rect 75822 63306 75828 63478
rect 75862 63306 75868 63478
rect 75822 63294 75868 63306
rect 76480 63478 76526 63490
rect 76480 63306 76486 63478
rect 76520 63306 76526 63478
rect 76480 63294 76526 63306
rect 77138 63478 77184 63490
rect 77138 63306 77144 63478
rect 77178 63306 77184 63478
rect 77138 63294 77184 63306
rect 77796 63478 77842 63490
rect 77796 63306 77802 63478
rect 77836 63306 77842 63478
rect 77796 63294 77842 63306
rect 71300 62804 71346 62816
rect 71300 62632 71306 62804
rect 71340 62632 71346 62804
rect 71300 62620 71346 62632
rect 71958 62804 72004 62816
rect 71958 62632 71964 62804
rect 71998 62632 72004 62804
rect 71958 62620 72004 62632
rect 72616 62804 72662 62816
rect 72616 62632 72622 62804
rect 72656 62632 72662 62804
rect 73274 62804 73320 62816
rect 73274 62776 73280 62804
rect 72616 62620 72662 62632
rect 73260 62632 73280 62776
rect 73314 62776 73320 62804
rect 73932 62804 73978 62816
rect 73314 62632 73336 62776
rect 42378 62582 42574 62588
rect 42378 62548 42390 62582
rect 42562 62548 42574 62582
rect 42378 62542 42574 62548
rect 43072 62582 43268 62588
rect 43072 62548 43084 62582
rect 43256 62548 43268 62582
rect 43072 62542 43268 62548
rect 43766 62582 43962 62588
rect 43766 62548 43778 62582
rect 43950 62548 43962 62582
rect 43766 62542 43962 62548
rect 44460 62582 44656 62588
rect 44460 62548 44472 62582
rect 44644 62548 44656 62582
rect 44460 62542 44656 62548
rect 45154 62582 45350 62588
rect 45154 62548 45166 62582
rect 45338 62548 45350 62582
rect 45154 62542 45350 62548
rect 46386 62580 46582 62586
rect 46386 62546 46398 62580
rect 46570 62546 46582 62580
rect 46386 62540 46582 62546
rect 47080 62580 47276 62586
rect 47080 62546 47092 62580
rect 47264 62546 47276 62580
rect 47080 62540 47276 62546
rect 47774 62580 47970 62586
rect 47774 62546 47786 62580
rect 47958 62546 47970 62580
rect 47774 62540 47970 62546
rect 48468 62580 48664 62586
rect 48468 62546 48480 62580
rect 48652 62546 48664 62580
rect 48468 62540 48664 62546
rect 49162 62580 49358 62586
rect 49162 62546 49174 62580
rect 49346 62546 49358 62580
rect 49162 62540 49358 62546
rect 50398 62580 50594 62586
rect 50398 62546 50410 62580
rect 50582 62546 50594 62580
rect 50398 62540 50594 62546
rect 51092 62580 51288 62586
rect 51092 62546 51104 62580
rect 51276 62546 51288 62580
rect 51092 62540 51288 62546
rect 51786 62580 51982 62586
rect 51786 62546 51798 62580
rect 51970 62546 51982 62580
rect 51786 62540 51982 62546
rect 52480 62580 52676 62586
rect 52480 62546 52492 62580
rect 52664 62546 52676 62580
rect 52480 62540 52676 62546
rect 53174 62580 53370 62586
rect 53174 62546 53186 62580
rect 53358 62546 53370 62580
rect 53174 62540 53370 62546
rect 54408 62580 54604 62586
rect 54408 62546 54420 62580
rect 54592 62546 54604 62580
rect 54408 62540 54604 62546
rect 55102 62580 55298 62586
rect 55102 62546 55114 62580
rect 55286 62546 55298 62580
rect 55102 62540 55298 62546
rect 55796 62580 55992 62586
rect 55796 62546 55808 62580
rect 55980 62546 55992 62580
rect 55796 62540 55992 62546
rect 56490 62580 56686 62586
rect 56490 62546 56502 62580
rect 56674 62546 56686 62580
rect 56490 62540 56686 62546
rect 57184 62580 57380 62586
rect 57184 62546 57196 62580
rect 57368 62546 57380 62580
rect 57184 62540 57380 62546
rect 19560 62330 19756 62336
rect 19560 62296 19572 62330
rect 19744 62296 19756 62330
rect 954 62280 1150 62286
rect 954 62246 966 62280
rect 1138 62246 1150 62280
rect 954 62240 1150 62246
rect 1648 62280 1844 62286
rect 1648 62246 1660 62280
rect 1832 62246 1844 62280
rect 1648 62240 1844 62246
rect 2342 62280 2538 62286
rect 6296 62282 6492 62288
rect 2342 62246 2354 62280
rect 2526 62246 2538 62280
rect 2342 62240 2538 62246
rect 3622 62276 3818 62282
rect 3622 62242 3634 62276
rect 3806 62242 3818 62276
rect 3622 62236 3818 62242
rect 4316 62276 4512 62282
rect 4316 62242 4328 62276
rect 4500 62242 4512 62276
rect 4316 62236 4512 62242
rect 5010 62276 5206 62282
rect 5010 62242 5022 62276
rect 5194 62242 5206 62276
rect 6296 62248 6308 62282
rect 6480 62248 6492 62282
rect 6296 62242 6492 62248
rect 6990 62282 7186 62288
rect 6990 62248 7002 62282
rect 7174 62248 7186 62282
rect 6990 62242 7186 62248
rect 7684 62282 7880 62288
rect 7684 62248 7696 62282
rect 7868 62248 7880 62282
rect 7684 62242 7880 62248
rect 8942 62282 9138 62288
rect 8942 62248 8954 62282
rect 9126 62248 9138 62282
rect 8942 62242 9138 62248
rect 9636 62282 9832 62288
rect 9636 62248 9648 62282
rect 9820 62248 9832 62282
rect 9636 62242 9832 62248
rect 10330 62282 10526 62288
rect 14250 62282 14446 62288
rect 10330 62248 10342 62282
rect 10514 62248 10526 62282
rect 10330 62242 10526 62248
rect 11596 62276 11792 62282
rect 11596 62242 11608 62276
rect 11780 62242 11792 62276
rect 5010 62236 5206 62242
rect 11596 62236 11792 62242
rect 12290 62276 12486 62282
rect 12290 62242 12302 62276
rect 12474 62242 12486 62276
rect 12290 62236 12486 62242
rect 12984 62276 13180 62282
rect 12984 62242 12996 62276
rect 13168 62242 13180 62276
rect 14250 62248 14262 62282
rect 14434 62248 14446 62282
rect 14250 62242 14446 62248
rect 14944 62282 15140 62288
rect 14944 62248 14956 62282
rect 15128 62248 15140 62282
rect 14944 62242 15140 62248
rect 15638 62282 15834 62288
rect 15638 62248 15650 62282
rect 15822 62248 15834 62282
rect 15638 62242 15834 62248
rect 16876 62286 17072 62292
rect 16876 62252 16888 62286
rect 17060 62252 17072 62286
rect 16876 62246 17072 62252
rect 17570 62286 17766 62292
rect 17570 62252 17582 62286
rect 17754 62252 17766 62286
rect 17570 62246 17766 62252
rect 18264 62286 18460 62292
rect 19560 62290 19756 62296
rect 20254 62330 20450 62336
rect 20254 62296 20266 62330
rect 20438 62296 20450 62330
rect 20254 62290 20450 62296
rect 18264 62252 18276 62286
rect 18448 62252 18460 62286
rect 18264 62246 18460 62252
rect 12984 62236 13180 62242
rect 42378 61924 42574 61930
rect 42378 61890 42390 61924
rect 42562 61890 42574 61924
rect 42378 61884 42574 61890
rect 43072 61924 43268 61930
rect 43072 61890 43084 61924
rect 43256 61890 43268 61924
rect 43072 61884 43268 61890
rect 43766 61924 43962 61930
rect 43766 61890 43778 61924
rect 43950 61890 43962 61924
rect 43766 61884 43962 61890
rect 44460 61924 44656 61930
rect 44460 61890 44472 61924
rect 44644 61890 44656 61924
rect 44460 61884 44656 61890
rect 45154 61924 45350 61930
rect 45154 61890 45166 61924
rect 45338 61890 45350 61924
rect 45154 61884 45350 61890
rect 46386 61922 46582 61928
rect 46386 61888 46398 61922
rect 46570 61888 46582 61922
rect 46386 61882 46582 61888
rect 47080 61922 47276 61928
rect 47080 61888 47092 61922
rect 47264 61888 47276 61922
rect 47080 61882 47276 61888
rect 47774 61922 47970 61928
rect 47774 61888 47786 61922
rect 47958 61888 47970 61922
rect 47774 61882 47970 61888
rect 48468 61922 48664 61928
rect 48468 61888 48480 61922
rect 48652 61888 48664 61922
rect 48468 61882 48664 61888
rect 49162 61922 49358 61928
rect 49162 61888 49174 61922
rect 49346 61888 49358 61922
rect 49162 61882 49358 61888
rect 50398 61922 50594 61928
rect 50398 61888 50410 61922
rect 50582 61888 50594 61922
rect 50398 61882 50594 61888
rect 51092 61922 51288 61928
rect 51092 61888 51104 61922
rect 51276 61888 51288 61922
rect 51092 61882 51288 61888
rect 51786 61922 51982 61928
rect 51786 61888 51798 61922
rect 51970 61888 51982 61922
rect 51786 61882 51982 61888
rect 52480 61922 52676 61928
rect 52480 61888 52492 61922
rect 52664 61888 52676 61922
rect 52480 61882 52676 61888
rect 53174 61922 53370 61928
rect 53174 61888 53186 61922
rect 53358 61888 53370 61922
rect 53174 61882 53370 61888
rect 54408 61922 54604 61928
rect 54408 61888 54420 61922
rect 54592 61888 54604 61922
rect 54408 61882 54604 61888
rect 55102 61922 55298 61928
rect 55102 61888 55114 61922
rect 55286 61888 55298 61922
rect 55102 61882 55298 61888
rect 55796 61922 55992 61928
rect 55796 61888 55808 61922
rect 55980 61888 55992 61922
rect 55796 61882 55992 61888
rect 56490 61922 56686 61928
rect 56490 61888 56502 61922
rect 56674 61888 56686 61922
rect 56490 61882 56686 61888
rect 57184 61922 57380 61928
rect 57184 61888 57196 61922
rect 57368 61888 57380 61922
rect 57184 61882 57380 61888
rect 71300 61816 71346 61828
rect 19560 61672 19756 61678
rect 19560 61638 19572 61672
rect 19744 61638 19756 61672
rect 954 61622 1150 61628
rect 954 61588 966 61622
rect 1138 61588 1150 61622
rect 954 61582 1150 61588
rect 1648 61622 1844 61628
rect 1648 61588 1660 61622
rect 1832 61588 1844 61622
rect 1648 61582 1844 61588
rect 2342 61622 2538 61628
rect 6296 61624 6492 61630
rect 2342 61588 2354 61622
rect 2526 61588 2538 61622
rect 2342 61582 2538 61588
rect 3622 61618 3818 61624
rect 3622 61584 3634 61618
rect 3806 61584 3818 61618
rect 3622 61578 3818 61584
rect 4316 61618 4512 61624
rect 4316 61584 4328 61618
rect 4500 61584 4512 61618
rect 4316 61578 4512 61584
rect 5010 61618 5206 61624
rect 5010 61584 5022 61618
rect 5194 61584 5206 61618
rect 6296 61590 6308 61624
rect 6480 61590 6492 61624
rect 6296 61584 6492 61590
rect 6990 61624 7186 61630
rect 6990 61590 7002 61624
rect 7174 61590 7186 61624
rect 6990 61584 7186 61590
rect 7684 61624 7880 61630
rect 7684 61590 7696 61624
rect 7868 61590 7880 61624
rect 7684 61584 7880 61590
rect 8942 61624 9138 61630
rect 8942 61590 8954 61624
rect 9126 61590 9138 61624
rect 8942 61584 9138 61590
rect 9636 61624 9832 61630
rect 9636 61590 9648 61624
rect 9820 61590 9832 61624
rect 9636 61584 9832 61590
rect 10330 61624 10526 61630
rect 14250 61624 14446 61630
rect 10330 61590 10342 61624
rect 10514 61590 10526 61624
rect 10330 61584 10526 61590
rect 11596 61618 11792 61624
rect 11596 61584 11608 61618
rect 11780 61584 11792 61618
rect 5010 61578 5206 61584
rect 11596 61578 11792 61584
rect 12290 61618 12486 61624
rect 12290 61584 12302 61618
rect 12474 61584 12486 61618
rect 12290 61578 12486 61584
rect 12984 61618 13180 61624
rect 12984 61584 12996 61618
rect 13168 61584 13180 61618
rect 14250 61590 14262 61624
rect 14434 61590 14446 61624
rect 14250 61584 14446 61590
rect 14944 61624 15140 61630
rect 14944 61590 14956 61624
rect 15128 61590 15140 61624
rect 14944 61584 15140 61590
rect 15638 61624 15834 61630
rect 15638 61590 15650 61624
rect 15822 61590 15834 61624
rect 15638 61584 15834 61590
rect 16876 61628 17072 61634
rect 16876 61594 16888 61628
rect 17060 61594 17072 61628
rect 16876 61588 17072 61594
rect 17570 61628 17766 61634
rect 17570 61594 17582 61628
rect 17754 61594 17766 61628
rect 17570 61588 17766 61594
rect 18264 61628 18460 61634
rect 19560 61632 19756 61638
rect 20254 61672 20450 61678
rect 20254 61638 20266 61672
rect 20438 61638 20450 61672
rect 20254 61632 20450 61638
rect 71008 61670 71224 61816
rect 18264 61594 18276 61628
rect 18448 61594 18460 61628
rect 18264 61588 18460 61594
rect 12984 61578 13180 61584
rect 42378 61266 42574 61272
rect 42378 61232 42390 61266
rect 42562 61232 42574 61266
rect 42378 61226 42574 61232
rect 43072 61266 43268 61272
rect 43072 61232 43084 61266
rect 43256 61232 43268 61266
rect 43072 61226 43268 61232
rect 43766 61266 43962 61272
rect 43766 61232 43778 61266
rect 43950 61232 43962 61266
rect 43766 61226 43962 61232
rect 44460 61266 44656 61272
rect 44460 61232 44472 61266
rect 44644 61232 44656 61266
rect 44460 61226 44656 61232
rect 45154 61266 45350 61272
rect 45154 61232 45166 61266
rect 45338 61232 45350 61266
rect 45154 61226 45350 61232
rect 46386 61264 46582 61270
rect 46386 61230 46398 61264
rect 46570 61230 46582 61264
rect 46386 61224 46582 61230
rect 47080 61264 47276 61270
rect 47080 61230 47092 61264
rect 47264 61230 47276 61264
rect 47080 61224 47276 61230
rect 47774 61264 47970 61270
rect 47774 61230 47786 61264
rect 47958 61230 47970 61264
rect 47774 61224 47970 61230
rect 48468 61264 48664 61270
rect 48468 61230 48480 61264
rect 48652 61230 48664 61264
rect 48468 61224 48664 61230
rect 49162 61264 49358 61270
rect 49162 61230 49174 61264
rect 49346 61230 49358 61264
rect 49162 61224 49358 61230
rect 50398 61264 50594 61270
rect 50398 61230 50410 61264
rect 50582 61230 50594 61264
rect 50398 61224 50594 61230
rect 51092 61264 51288 61270
rect 51092 61230 51104 61264
rect 51276 61230 51288 61264
rect 51092 61224 51288 61230
rect 51786 61264 51982 61270
rect 51786 61230 51798 61264
rect 51970 61230 51982 61264
rect 51786 61224 51982 61230
rect 52480 61264 52676 61270
rect 52480 61230 52492 61264
rect 52664 61230 52676 61264
rect 52480 61224 52676 61230
rect 53174 61264 53370 61270
rect 53174 61230 53186 61264
rect 53358 61230 53370 61264
rect 53174 61224 53370 61230
rect 54408 61264 54604 61270
rect 54408 61230 54420 61264
rect 54592 61230 54604 61264
rect 54408 61224 54604 61230
rect 55102 61264 55298 61270
rect 55102 61230 55114 61264
rect 55286 61230 55298 61264
rect 55102 61224 55298 61230
rect 55796 61264 55992 61270
rect 55796 61230 55808 61264
rect 55980 61230 55992 61264
rect 55796 61224 55992 61230
rect 56490 61264 56686 61270
rect 56490 61230 56502 61264
rect 56674 61230 56686 61264
rect 56490 61224 56686 61230
rect 57184 61264 57380 61270
rect 57184 61230 57196 61264
rect 57368 61230 57380 61264
rect 57184 61224 57380 61230
rect 8374 61180 8588 61192
rect 5714 61104 5962 61116
rect 3080 61070 3310 61082
rect 3080 61020 3086 61070
rect 2396 60970 3086 61020
rect 954 60964 1150 60970
rect 954 60930 966 60964
rect 1138 60930 1150 60964
rect 954 60924 1150 60930
rect 1648 60964 1844 60970
rect 1648 60930 1660 60964
rect 1832 60930 1844 60964
rect 1648 60924 1844 60930
rect 2342 60964 3086 60970
rect 2342 60930 2354 60964
rect 2526 60930 3086 60964
rect 2342 60924 3086 60930
rect 2396 60860 3086 60924
rect 3080 60716 3086 60860
rect 3304 60716 3310 61070
rect 5714 61020 5720 61104
rect 5106 60966 5720 61020
rect 3622 60960 3818 60966
rect 3622 60926 3634 60960
rect 3806 60926 3818 60960
rect 3622 60920 3818 60926
rect 4316 60960 4512 60966
rect 4316 60926 4328 60960
rect 4500 60926 4512 60960
rect 4316 60920 4512 60926
rect 5010 60960 5720 60966
rect 5010 60926 5022 60960
rect 5194 60926 5720 60960
rect 5010 60920 5720 60926
rect 5106 60852 5720 60920
rect 5714 60742 5720 60852
rect 5956 60742 5962 61104
rect 8374 61062 8380 61180
rect 7748 60972 8380 61062
rect 6296 60966 6492 60972
rect 6296 60932 6308 60966
rect 6480 60932 6492 60966
rect 6296 60926 6492 60932
rect 6990 60966 7186 60972
rect 6990 60932 7002 60966
rect 7174 60932 7186 60966
rect 6990 60926 7186 60932
rect 7684 60966 8380 60972
rect 7684 60932 7696 60966
rect 7868 60932 8380 60966
rect 7684 60926 8380 60932
rect 7748 60826 8380 60926
rect 5714 60730 5962 60742
rect 3080 60704 3310 60716
rect 8374 60692 8380 60826
rect 8582 60692 8588 61180
rect 18866 61162 19088 61174
rect 13700 61128 13880 61140
rect 11050 61096 11280 61108
rect 11050 61010 11056 61096
rect 10408 60972 11056 61010
rect 8942 60966 9138 60972
rect 8942 60932 8954 60966
rect 9126 60932 9138 60966
rect 8942 60926 9138 60932
rect 9636 60966 9832 60972
rect 9636 60932 9648 60966
rect 9820 60932 9832 60966
rect 9636 60926 9832 60932
rect 10330 60966 11056 60972
rect 10330 60932 10342 60966
rect 10514 60932 11056 60966
rect 10330 60926 11056 60932
rect 10408 60818 11056 60926
rect 8374 60680 8588 60692
rect 11050 60658 11056 60818
rect 11274 60658 11280 61096
rect 13700 61002 13706 61128
rect 13016 60966 13706 61002
rect 11596 60960 11792 60966
rect 11596 60926 11608 60960
rect 11780 60926 11792 60960
rect 11596 60920 11792 60926
rect 12290 60960 12486 60966
rect 12290 60926 12302 60960
rect 12474 60926 12486 60960
rect 12290 60920 12486 60926
rect 12984 60960 13706 60966
rect 12984 60926 12996 60960
rect 13168 60926 13706 60960
rect 12984 60920 13706 60926
rect 13016 60884 13706 60920
rect 13700 60700 13706 60884
rect 13874 60700 13880 61128
rect 16316 61070 16582 61082
rect 16316 61028 16322 61070
rect 15692 60972 16322 61028
rect 14250 60966 14446 60972
rect 14250 60932 14262 60966
rect 14434 60932 14446 60966
rect 14250 60926 14446 60932
rect 14944 60966 15140 60972
rect 14944 60932 14956 60966
rect 15128 60932 15140 60966
rect 14944 60926 15140 60932
rect 15638 60966 16322 60972
rect 15638 60932 15650 60966
rect 15822 60932 16322 60966
rect 15638 60926 16322 60932
rect 15692 60910 16322 60926
rect 16316 60800 16322 60910
rect 16576 60800 16582 61070
rect 18866 61052 18872 61162
rect 18318 60976 18872 61052
rect 16876 60970 17072 60976
rect 16876 60936 16888 60970
rect 17060 60936 17072 60970
rect 16876 60930 17072 60936
rect 17570 60970 17766 60976
rect 17570 60936 17582 60970
rect 17754 60936 17766 60970
rect 17570 60930 17766 60936
rect 18264 60970 18872 60976
rect 18264 60936 18276 60970
rect 18448 60936 18872 60970
rect 18264 60930 18872 60936
rect 18318 60894 18872 60930
rect 18866 60816 18872 60894
rect 19082 60816 19088 61162
rect 57706 61090 58040 61298
rect 19560 61014 19756 61020
rect 19560 60980 19572 61014
rect 19744 60980 19756 61014
rect 19560 60974 19756 60980
rect 20254 61014 20450 61020
rect 20254 60980 20266 61014
rect 20438 60980 20450 61014
rect 20254 60974 20450 60980
rect 18866 60804 19088 60816
rect 42726 60810 45372 60898
rect 16316 60788 16582 60800
rect 13700 60688 13880 60700
rect 11050 60646 11280 60658
rect 42726 60608 43024 60810
rect 45198 60608 45372 60810
rect 42726 60496 45372 60608
rect 46720 60810 49366 60898
rect 46720 60608 47018 60810
rect 49192 60608 49366 60810
rect 46720 60496 49366 60608
rect 50742 60810 53388 60898
rect 50742 60608 51040 60810
rect 53214 60608 53388 60810
rect 50742 60496 53388 60608
rect 54764 60810 57410 60898
rect 54764 60608 55062 60810
rect 57236 60608 57410 60810
rect 54764 60496 57410 60608
rect 57706 60588 57798 61090
rect 57940 60948 58040 61090
rect 59906 60948 60318 60972
rect 57940 60764 60318 60948
rect 57940 60588 58040 60764
rect 57706 60396 58040 60588
rect 19560 60356 19756 60362
rect 19560 60322 19572 60356
rect 19744 60322 19756 60356
rect 954 60306 1150 60312
rect 954 60272 966 60306
rect 1138 60272 1150 60306
rect 954 60266 1150 60272
rect 1648 60306 1844 60312
rect 1648 60272 1660 60306
rect 1832 60272 1844 60306
rect 1648 60266 1844 60272
rect 2342 60306 2538 60312
rect 6296 60308 6492 60314
rect 2342 60272 2354 60306
rect 2526 60272 2538 60306
rect 2342 60266 2538 60272
rect 3622 60302 3818 60308
rect 3622 60268 3634 60302
rect 3806 60268 3818 60302
rect 3622 60262 3818 60268
rect 4316 60302 4512 60308
rect 4316 60268 4328 60302
rect 4500 60268 4512 60302
rect 4316 60262 4512 60268
rect 5010 60302 5206 60308
rect 5010 60268 5022 60302
rect 5194 60268 5206 60302
rect 6296 60274 6308 60308
rect 6480 60274 6492 60308
rect 6296 60268 6492 60274
rect 6990 60308 7186 60314
rect 6990 60274 7002 60308
rect 7174 60274 7186 60308
rect 6990 60268 7186 60274
rect 7684 60308 7880 60314
rect 7684 60274 7696 60308
rect 7868 60274 7880 60308
rect 7684 60268 7880 60274
rect 8942 60308 9138 60314
rect 8942 60274 8954 60308
rect 9126 60274 9138 60308
rect 8942 60268 9138 60274
rect 9636 60308 9832 60314
rect 9636 60274 9648 60308
rect 9820 60274 9832 60308
rect 9636 60268 9832 60274
rect 10330 60308 10526 60314
rect 14250 60308 14446 60314
rect 10330 60274 10342 60308
rect 10514 60274 10526 60308
rect 10330 60268 10526 60274
rect 11596 60302 11792 60308
rect 11596 60268 11608 60302
rect 11780 60268 11792 60302
rect 5010 60262 5206 60268
rect 11596 60262 11792 60268
rect 12290 60302 12486 60308
rect 12290 60268 12302 60302
rect 12474 60268 12486 60302
rect 12290 60262 12486 60268
rect 12984 60302 13180 60308
rect 12984 60268 12996 60302
rect 13168 60268 13180 60302
rect 14250 60274 14262 60308
rect 14434 60274 14446 60308
rect 14250 60268 14446 60274
rect 14944 60308 15140 60314
rect 14944 60274 14956 60308
rect 15128 60274 15140 60308
rect 14944 60268 15140 60274
rect 15638 60308 15834 60314
rect 15638 60274 15650 60308
rect 15822 60274 15834 60308
rect 15638 60268 15834 60274
rect 16876 60312 17072 60318
rect 16876 60278 16888 60312
rect 17060 60278 17072 60312
rect 16876 60272 17072 60278
rect 17570 60312 17766 60318
rect 17570 60278 17582 60312
rect 17754 60278 17766 60312
rect 17570 60272 17766 60278
rect 18264 60312 18460 60318
rect 19560 60316 19756 60322
rect 20254 60356 20450 60362
rect 20254 60322 20266 60356
rect 20438 60322 20450 60356
rect 20254 60316 20450 60322
rect 42370 60358 42566 60364
rect 42370 60324 42382 60358
rect 42554 60324 42566 60358
rect 42370 60318 42566 60324
rect 43064 60358 43260 60364
rect 43064 60324 43076 60358
rect 43248 60324 43260 60358
rect 43064 60318 43260 60324
rect 43758 60358 43954 60364
rect 43758 60324 43770 60358
rect 43942 60324 43954 60358
rect 43758 60318 43954 60324
rect 44452 60358 44648 60364
rect 44452 60324 44464 60358
rect 44636 60324 44648 60358
rect 44452 60318 44648 60324
rect 45146 60358 45342 60364
rect 45146 60324 45158 60358
rect 45330 60324 45342 60358
rect 45146 60318 45342 60324
rect 46364 60358 46560 60364
rect 46364 60324 46376 60358
rect 46548 60324 46560 60358
rect 46364 60318 46560 60324
rect 47058 60358 47254 60364
rect 47058 60324 47070 60358
rect 47242 60324 47254 60358
rect 47058 60318 47254 60324
rect 47752 60358 47948 60364
rect 47752 60324 47764 60358
rect 47936 60324 47948 60358
rect 47752 60318 47948 60324
rect 48446 60358 48642 60364
rect 48446 60324 48458 60358
rect 48630 60324 48642 60358
rect 48446 60318 48642 60324
rect 49140 60358 49336 60364
rect 49140 60324 49152 60358
rect 49324 60324 49336 60358
rect 49140 60318 49336 60324
rect 50386 60358 50582 60364
rect 50386 60324 50398 60358
rect 50570 60324 50582 60358
rect 50386 60318 50582 60324
rect 51080 60358 51276 60364
rect 51080 60324 51092 60358
rect 51264 60324 51276 60358
rect 51080 60318 51276 60324
rect 51774 60358 51970 60364
rect 51774 60324 51786 60358
rect 51958 60324 51970 60358
rect 51774 60318 51970 60324
rect 52468 60358 52664 60364
rect 52468 60324 52480 60358
rect 52652 60324 52664 60358
rect 52468 60318 52664 60324
rect 53162 60358 53358 60364
rect 53162 60324 53174 60358
rect 53346 60324 53358 60358
rect 53162 60318 53358 60324
rect 54408 60358 54604 60364
rect 54408 60324 54420 60358
rect 54592 60324 54604 60358
rect 54408 60318 54604 60324
rect 55102 60358 55298 60364
rect 55102 60324 55114 60358
rect 55286 60324 55298 60358
rect 55102 60318 55298 60324
rect 55796 60358 55992 60364
rect 55796 60324 55808 60358
rect 55980 60324 55992 60358
rect 55796 60318 55992 60324
rect 56490 60358 56686 60364
rect 56490 60324 56502 60358
rect 56674 60324 56686 60358
rect 56490 60318 56686 60324
rect 57184 60358 57380 60364
rect 57184 60324 57196 60358
rect 57368 60324 57380 60358
rect 57184 60318 57380 60324
rect 18264 60278 18276 60312
rect 18448 60278 18460 60312
rect 18264 60272 18460 60278
rect 12984 60262 13180 60268
rect 944 59636 2576 59694
rect 944 59566 1058 59636
rect 2462 59566 2576 59636
rect 944 59490 2576 59566
rect 3612 59632 5244 59690
rect 3612 59562 3726 59632
rect 5130 59562 5244 59632
rect 3612 59486 5244 59562
rect 6286 59638 7918 59696
rect 6286 59568 6400 59638
rect 7804 59568 7918 59638
rect 6286 59492 7918 59568
rect 8932 59638 10564 59696
rect 8932 59568 9046 59638
rect 10450 59568 10564 59638
rect 8932 59492 10564 59568
rect 11586 59632 13218 59690
rect 11586 59562 11700 59632
rect 13104 59562 13218 59632
rect 11586 59486 13218 59562
rect 14240 59638 15872 59696
rect 14240 59568 14354 59638
rect 15758 59568 15872 59638
rect 14240 59492 15872 59568
rect 16866 59642 18498 59700
rect 16866 59572 16980 59642
rect 18384 59572 18498 59642
rect 16866 59496 18498 59572
rect 19364 59656 20600 59726
rect 42370 59700 42566 59706
rect 42370 59666 42382 59700
rect 42554 59666 42566 59700
rect 42370 59660 42566 59666
rect 43064 59700 43260 59706
rect 43064 59666 43076 59700
rect 43248 59666 43260 59700
rect 43064 59660 43260 59666
rect 43758 59700 43954 59706
rect 43758 59666 43770 59700
rect 43942 59666 43954 59700
rect 43758 59660 43954 59666
rect 44452 59700 44648 59706
rect 44452 59666 44464 59700
rect 44636 59666 44648 59700
rect 44452 59660 44648 59666
rect 45146 59700 45342 59706
rect 45146 59666 45158 59700
rect 45330 59666 45342 59700
rect 45146 59660 45342 59666
rect 46364 59700 46560 59706
rect 46364 59666 46376 59700
rect 46548 59666 46560 59700
rect 46364 59660 46560 59666
rect 47058 59700 47254 59706
rect 47058 59666 47070 59700
rect 47242 59666 47254 59700
rect 47058 59660 47254 59666
rect 47752 59700 47948 59706
rect 47752 59666 47764 59700
rect 47936 59666 47948 59700
rect 47752 59660 47948 59666
rect 48446 59700 48642 59706
rect 48446 59666 48458 59700
rect 48630 59666 48642 59700
rect 48446 59660 48642 59666
rect 49140 59700 49336 59706
rect 49140 59666 49152 59700
rect 49324 59666 49336 59700
rect 49140 59660 49336 59666
rect 50386 59700 50582 59706
rect 50386 59666 50398 59700
rect 50570 59666 50582 59700
rect 50386 59660 50582 59666
rect 51080 59700 51276 59706
rect 51080 59666 51092 59700
rect 51264 59666 51276 59700
rect 51080 59660 51276 59666
rect 51774 59700 51970 59706
rect 51774 59666 51786 59700
rect 51958 59666 51970 59700
rect 51774 59660 51970 59666
rect 52468 59700 52664 59706
rect 52468 59666 52480 59700
rect 52652 59666 52664 59700
rect 52468 59660 52664 59666
rect 53162 59700 53358 59706
rect 53162 59666 53174 59700
rect 53346 59666 53358 59700
rect 53162 59660 53358 59666
rect 54408 59700 54604 59706
rect 54408 59666 54420 59700
rect 54592 59666 54604 59700
rect 54408 59660 54604 59666
rect 55102 59700 55298 59706
rect 55102 59666 55114 59700
rect 55286 59666 55298 59700
rect 55102 59660 55298 59666
rect 55796 59700 55992 59706
rect 55796 59666 55808 59700
rect 55980 59666 55992 59700
rect 55796 59660 55992 59666
rect 56490 59700 56686 59706
rect 56490 59666 56502 59700
rect 56674 59666 56686 59700
rect 56490 59660 56686 59666
rect 57184 59700 57380 59706
rect 57184 59666 57196 59700
rect 57368 59666 57380 59700
rect 57184 59660 57380 59666
rect 19364 59548 19534 59656
rect 20492 59548 20600 59656
rect 19364 59456 20600 59548
rect 19532 59352 19728 59358
rect 19532 59318 19544 59352
rect 19716 59318 19728 59352
rect 926 59302 1122 59308
rect 926 59268 938 59302
rect 1110 59268 1122 59302
rect 926 59262 1122 59268
rect 1620 59302 1816 59308
rect 1620 59268 1632 59302
rect 1804 59268 1816 59302
rect 1620 59262 1816 59268
rect 2314 59302 2510 59308
rect 6268 59304 6464 59310
rect 2314 59268 2326 59302
rect 2498 59268 2510 59302
rect 2314 59262 2510 59268
rect 3594 59298 3790 59304
rect 3594 59264 3606 59298
rect 3778 59264 3790 59298
rect 3594 59258 3790 59264
rect 4288 59298 4484 59304
rect 4288 59264 4300 59298
rect 4472 59264 4484 59298
rect 4288 59258 4484 59264
rect 4982 59298 5178 59304
rect 4982 59264 4994 59298
rect 5166 59264 5178 59298
rect 6268 59270 6280 59304
rect 6452 59270 6464 59304
rect 6268 59264 6464 59270
rect 6962 59304 7158 59310
rect 6962 59270 6974 59304
rect 7146 59270 7158 59304
rect 6962 59264 7158 59270
rect 7656 59304 7852 59310
rect 7656 59270 7668 59304
rect 7840 59270 7852 59304
rect 7656 59264 7852 59270
rect 8914 59304 9110 59310
rect 8914 59270 8926 59304
rect 9098 59270 9110 59304
rect 8914 59264 9110 59270
rect 9608 59304 9804 59310
rect 9608 59270 9620 59304
rect 9792 59270 9804 59304
rect 9608 59264 9804 59270
rect 10302 59304 10498 59310
rect 14222 59304 14418 59310
rect 10302 59270 10314 59304
rect 10486 59270 10498 59304
rect 10302 59264 10498 59270
rect 11568 59298 11764 59304
rect 11568 59264 11580 59298
rect 11752 59264 11764 59298
rect 4982 59258 5178 59264
rect 11568 59258 11764 59264
rect 12262 59298 12458 59304
rect 12262 59264 12274 59298
rect 12446 59264 12458 59298
rect 12262 59258 12458 59264
rect 12956 59298 13152 59304
rect 12956 59264 12968 59298
rect 13140 59264 13152 59298
rect 14222 59270 14234 59304
rect 14406 59270 14418 59304
rect 14222 59264 14418 59270
rect 14916 59304 15112 59310
rect 14916 59270 14928 59304
rect 15100 59270 15112 59304
rect 14916 59264 15112 59270
rect 15610 59304 15806 59310
rect 15610 59270 15622 59304
rect 15794 59270 15806 59304
rect 15610 59264 15806 59270
rect 16848 59308 17044 59314
rect 16848 59274 16860 59308
rect 17032 59274 17044 59308
rect 16848 59268 17044 59274
rect 17542 59308 17738 59314
rect 17542 59274 17554 59308
rect 17726 59274 17738 59308
rect 17542 59268 17738 59274
rect 18236 59308 18432 59314
rect 19532 59312 19728 59318
rect 20226 59352 20422 59358
rect 20226 59318 20238 59352
rect 20410 59318 20422 59352
rect 20226 59312 20422 59318
rect 18236 59274 18248 59308
rect 18420 59274 18432 59308
rect 18236 59268 18432 59274
rect 12956 59258 13152 59264
rect 42370 59042 42566 59048
rect 42370 59008 42382 59042
rect 42554 59008 42566 59042
rect 42370 59002 42566 59008
rect 43064 59042 43260 59048
rect 43064 59008 43076 59042
rect 43248 59008 43260 59042
rect 43064 59002 43260 59008
rect 43758 59042 43954 59048
rect 43758 59008 43770 59042
rect 43942 59008 43954 59042
rect 43758 59002 43954 59008
rect 44452 59042 44648 59048
rect 44452 59008 44464 59042
rect 44636 59008 44648 59042
rect 44452 59002 44648 59008
rect 45146 59042 45342 59048
rect 45146 59008 45158 59042
rect 45330 59008 45342 59042
rect 45146 59002 45342 59008
rect 46364 59042 46560 59048
rect 46364 59008 46376 59042
rect 46548 59008 46560 59042
rect 46364 59002 46560 59008
rect 47058 59042 47254 59048
rect 47058 59008 47070 59042
rect 47242 59008 47254 59042
rect 47058 59002 47254 59008
rect 47752 59042 47948 59048
rect 47752 59008 47764 59042
rect 47936 59008 47948 59042
rect 47752 59002 47948 59008
rect 48446 59042 48642 59048
rect 48446 59008 48458 59042
rect 48630 59008 48642 59042
rect 48446 59002 48642 59008
rect 49140 59042 49336 59048
rect 49140 59008 49152 59042
rect 49324 59008 49336 59042
rect 49140 59002 49336 59008
rect 50386 59042 50582 59048
rect 50386 59008 50398 59042
rect 50570 59008 50582 59042
rect 50386 59002 50582 59008
rect 51080 59042 51276 59048
rect 51080 59008 51092 59042
rect 51264 59008 51276 59042
rect 51080 59002 51276 59008
rect 51774 59042 51970 59048
rect 51774 59008 51786 59042
rect 51958 59008 51970 59042
rect 51774 59002 51970 59008
rect 52468 59042 52664 59048
rect 52468 59008 52480 59042
rect 52652 59008 52664 59042
rect 52468 59002 52664 59008
rect 53162 59042 53358 59048
rect 53162 59008 53174 59042
rect 53346 59008 53358 59042
rect 53162 59002 53358 59008
rect 54408 59042 54604 59048
rect 54408 59008 54420 59042
rect 54592 59008 54604 59042
rect 54408 59002 54604 59008
rect 55102 59042 55298 59048
rect 55102 59008 55114 59042
rect 55286 59008 55298 59042
rect 55102 59002 55298 59008
rect 55796 59042 55992 59048
rect 55796 59008 55808 59042
rect 55980 59008 55992 59042
rect 55796 59002 55992 59008
rect 56490 59042 56686 59048
rect 56490 59008 56502 59042
rect 56674 59008 56686 59042
rect 56490 59002 56686 59008
rect 57184 59042 57380 59048
rect 57184 59008 57196 59042
rect 57368 59008 57380 59042
rect 57184 59002 57380 59008
rect 19532 58694 19728 58700
rect 19532 58660 19544 58694
rect 19716 58660 19728 58694
rect 926 58644 1122 58650
rect 926 58610 938 58644
rect 1110 58610 1122 58644
rect 926 58604 1122 58610
rect 1620 58644 1816 58650
rect 1620 58610 1632 58644
rect 1804 58610 1816 58644
rect 1620 58604 1816 58610
rect 2314 58644 2510 58650
rect 6268 58646 6464 58652
rect 2314 58610 2326 58644
rect 2498 58610 2510 58644
rect 2314 58604 2510 58610
rect 3594 58640 3790 58646
rect 3594 58606 3606 58640
rect 3778 58606 3790 58640
rect 3594 58600 3790 58606
rect 4288 58640 4484 58646
rect 4288 58606 4300 58640
rect 4472 58606 4484 58640
rect 4288 58600 4484 58606
rect 4982 58640 5178 58646
rect 4982 58606 4994 58640
rect 5166 58606 5178 58640
rect 6268 58612 6280 58646
rect 6452 58612 6464 58646
rect 6268 58606 6464 58612
rect 6962 58646 7158 58652
rect 6962 58612 6974 58646
rect 7146 58612 7158 58646
rect 6962 58606 7158 58612
rect 7656 58646 7852 58652
rect 7656 58612 7668 58646
rect 7840 58612 7852 58646
rect 7656 58606 7852 58612
rect 8914 58646 9110 58652
rect 8914 58612 8926 58646
rect 9098 58612 9110 58646
rect 8914 58606 9110 58612
rect 9608 58646 9804 58652
rect 9608 58612 9620 58646
rect 9792 58612 9804 58646
rect 9608 58606 9804 58612
rect 10302 58646 10498 58652
rect 14222 58646 14418 58652
rect 10302 58612 10314 58646
rect 10486 58612 10498 58646
rect 10302 58606 10498 58612
rect 11568 58640 11764 58646
rect 11568 58606 11580 58640
rect 11752 58606 11764 58640
rect 4982 58600 5178 58606
rect 11568 58600 11764 58606
rect 12262 58640 12458 58646
rect 12262 58606 12274 58640
rect 12446 58606 12458 58640
rect 12262 58600 12458 58606
rect 12956 58640 13152 58646
rect 12956 58606 12968 58640
rect 13140 58606 13152 58640
rect 14222 58612 14234 58646
rect 14406 58612 14418 58646
rect 14222 58606 14418 58612
rect 14916 58646 15112 58652
rect 14916 58612 14928 58646
rect 15100 58612 15112 58646
rect 14916 58606 15112 58612
rect 15610 58646 15806 58652
rect 15610 58612 15622 58646
rect 15794 58612 15806 58646
rect 15610 58606 15806 58612
rect 16848 58650 17044 58656
rect 16848 58616 16860 58650
rect 17032 58616 17044 58650
rect 16848 58610 17044 58616
rect 17542 58650 17738 58656
rect 17542 58616 17554 58650
rect 17726 58616 17738 58650
rect 17542 58610 17738 58616
rect 18236 58650 18432 58656
rect 19532 58654 19728 58660
rect 20226 58694 20422 58700
rect 20226 58660 20238 58694
rect 20410 58660 20422 58694
rect 20226 58654 20422 58660
rect 18236 58616 18248 58650
rect 18420 58616 18432 58650
rect 18236 58610 18432 58616
rect 12956 58600 13152 58606
rect 42370 58384 42566 58390
rect 42370 58350 42382 58384
rect 42554 58350 42566 58384
rect 42370 58344 42566 58350
rect 43064 58384 43260 58390
rect 43064 58350 43076 58384
rect 43248 58350 43260 58384
rect 43064 58344 43260 58350
rect 43758 58384 43954 58390
rect 43758 58350 43770 58384
rect 43942 58350 43954 58384
rect 43758 58344 43954 58350
rect 44452 58384 44648 58390
rect 44452 58350 44464 58384
rect 44636 58350 44648 58384
rect 44452 58344 44648 58350
rect 45146 58384 45342 58390
rect 45146 58350 45158 58384
rect 45330 58350 45342 58384
rect 45146 58344 45342 58350
rect 46364 58384 46560 58390
rect 46364 58350 46376 58384
rect 46548 58350 46560 58384
rect 46364 58344 46560 58350
rect 47058 58384 47254 58390
rect 47058 58350 47070 58384
rect 47242 58350 47254 58384
rect 47058 58344 47254 58350
rect 47752 58384 47948 58390
rect 47752 58350 47764 58384
rect 47936 58350 47948 58384
rect 47752 58344 47948 58350
rect 48446 58384 48642 58390
rect 48446 58350 48458 58384
rect 48630 58350 48642 58384
rect 48446 58344 48642 58350
rect 49140 58384 49336 58390
rect 49140 58350 49152 58384
rect 49324 58350 49336 58384
rect 49140 58344 49336 58350
rect 50386 58384 50582 58390
rect 50386 58350 50398 58384
rect 50570 58350 50582 58384
rect 50386 58344 50582 58350
rect 51080 58384 51276 58390
rect 51080 58350 51092 58384
rect 51264 58350 51276 58384
rect 51080 58344 51276 58350
rect 51774 58384 51970 58390
rect 51774 58350 51786 58384
rect 51958 58350 51970 58384
rect 51774 58344 51970 58350
rect 52468 58384 52664 58390
rect 52468 58350 52480 58384
rect 52652 58350 52664 58384
rect 52468 58344 52664 58350
rect 53162 58384 53358 58390
rect 53162 58350 53174 58384
rect 53346 58350 53358 58384
rect 53162 58344 53358 58350
rect 54408 58384 54604 58390
rect 54408 58350 54420 58384
rect 54592 58350 54604 58384
rect 54408 58344 54604 58350
rect 55102 58384 55298 58390
rect 55102 58350 55114 58384
rect 55286 58350 55298 58384
rect 55102 58344 55298 58350
rect 55796 58384 55992 58390
rect 55796 58350 55808 58384
rect 55980 58350 55992 58384
rect 55796 58344 55992 58350
rect 56490 58384 56686 58390
rect 56490 58350 56502 58384
rect 56674 58350 56686 58384
rect 56490 58344 56686 58350
rect 57184 58384 57380 58390
rect 57184 58350 57196 58384
rect 57368 58350 57380 58384
rect 57184 58344 57380 58350
rect 19532 58036 19728 58042
rect 19532 58002 19544 58036
rect 19716 58002 19728 58036
rect 926 57986 1122 57992
rect 926 57952 938 57986
rect 1110 57952 1122 57986
rect 926 57946 1122 57952
rect 1620 57986 1816 57992
rect 1620 57952 1632 57986
rect 1804 57952 1816 57986
rect 1620 57946 1816 57952
rect 2314 57986 2510 57992
rect 6268 57988 6464 57994
rect 2314 57952 2326 57986
rect 2498 57952 2510 57986
rect 2314 57946 2510 57952
rect 3594 57982 3790 57988
rect 3594 57948 3606 57982
rect 3778 57948 3790 57982
rect 3594 57942 3790 57948
rect 4288 57982 4484 57988
rect 4288 57948 4300 57982
rect 4472 57948 4484 57982
rect 4288 57942 4484 57948
rect 4982 57982 5178 57988
rect 4982 57948 4994 57982
rect 5166 57948 5178 57982
rect 6268 57954 6280 57988
rect 6452 57954 6464 57988
rect 6268 57948 6464 57954
rect 6962 57988 7158 57994
rect 6962 57954 6974 57988
rect 7146 57954 7158 57988
rect 6962 57948 7158 57954
rect 7656 57988 7852 57994
rect 7656 57954 7668 57988
rect 7840 57954 7852 57988
rect 7656 57948 7852 57954
rect 8914 57988 9110 57994
rect 8914 57954 8926 57988
rect 9098 57954 9110 57988
rect 8914 57948 9110 57954
rect 9608 57988 9804 57994
rect 9608 57954 9620 57988
rect 9792 57954 9804 57988
rect 9608 57948 9804 57954
rect 10302 57988 10498 57994
rect 14222 57988 14418 57994
rect 10302 57954 10314 57988
rect 10486 57954 10498 57988
rect 10302 57948 10498 57954
rect 11568 57982 11764 57988
rect 11568 57948 11580 57982
rect 11752 57948 11764 57982
rect 4982 57942 5178 57948
rect 11568 57942 11764 57948
rect 12262 57982 12458 57988
rect 12262 57948 12274 57982
rect 12446 57948 12458 57982
rect 12262 57942 12458 57948
rect 12956 57982 13152 57988
rect 12956 57948 12968 57982
rect 13140 57948 13152 57982
rect 14222 57954 14234 57988
rect 14406 57954 14418 57988
rect 14222 57948 14418 57954
rect 14916 57988 15112 57994
rect 14916 57954 14928 57988
rect 15100 57954 15112 57988
rect 14916 57948 15112 57954
rect 15610 57988 15806 57994
rect 15610 57954 15622 57988
rect 15794 57954 15806 57988
rect 15610 57948 15806 57954
rect 16848 57992 17044 57998
rect 16848 57958 16860 57992
rect 17032 57958 17044 57992
rect 16848 57952 17044 57958
rect 17542 57992 17738 57998
rect 17542 57958 17554 57992
rect 17726 57958 17738 57992
rect 17542 57952 17738 57958
rect 18236 57992 18432 57998
rect 19532 57996 19728 58002
rect 20226 58036 20422 58042
rect 20226 58002 20238 58036
rect 20410 58002 20422 58036
rect 20226 57996 20422 58002
rect 18236 57958 18248 57992
rect 18420 57958 18432 57992
rect 18236 57952 18432 57958
rect 12956 57942 13152 57948
rect 222 57716 554 57874
rect 222 56766 338 57716
rect 438 56766 554 57716
rect 42370 57726 42566 57732
rect 42370 57692 42382 57726
rect 42554 57692 42566 57726
rect 42370 57686 42566 57692
rect 43064 57726 43260 57732
rect 43064 57692 43076 57726
rect 43248 57692 43260 57726
rect 43064 57686 43260 57692
rect 43758 57726 43954 57732
rect 43758 57692 43770 57726
rect 43942 57692 43954 57726
rect 43758 57686 43954 57692
rect 44452 57726 44648 57732
rect 44452 57692 44464 57726
rect 44636 57692 44648 57726
rect 44452 57686 44648 57692
rect 45146 57726 45342 57732
rect 45146 57692 45158 57726
rect 45330 57692 45342 57726
rect 45146 57686 45342 57692
rect 46364 57726 46560 57732
rect 46364 57692 46376 57726
rect 46548 57692 46560 57726
rect 46364 57686 46560 57692
rect 47058 57726 47254 57732
rect 47058 57692 47070 57726
rect 47242 57692 47254 57726
rect 47058 57686 47254 57692
rect 47752 57726 47948 57732
rect 47752 57692 47764 57726
rect 47936 57692 47948 57726
rect 47752 57686 47948 57692
rect 48446 57726 48642 57732
rect 48446 57692 48458 57726
rect 48630 57692 48642 57726
rect 48446 57686 48642 57692
rect 49140 57726 49336 57732
rect 49140 57692 49152 57726
rect 49324 57692 49336 57726
rect 49140 57686 49336 57692
rect 50386 57726 50582 57732
rect 50386 57692 50398 57726
rect 50570 57692 50582 57726
rect 50386 57686 50582 57692
rect 51080 57726 51276 57732
rect 51080 57692 51092 57726
rect 51264 57692 51276 57726
rect 51080 57686 51276 57692
rect 51774 57726 51970 57732
rect 51774 57692 51786 57726
rect 51958 57692 51970 57726
rect 51774 57686 51970 57692
rect 52468 57726 52664 57732
rect 52468 57692 52480 57726
rect 52652 57692 52664 57726
rect 52468 57686 52664 57692
rect 53162 57726 53358 57732
rect 53162 57692 53174 57726
rect 53346 57692 53358 57726
rect 53162 57686 53358 57692
rect 54408 57726 54604 57732
rect 54408 57692 54420 57726
rect 54592 57692 54604 57726
rect 54408 57686 54604 57692
rect 55102 57726 55298 57732
rect 55102 57692 55114 57726
rect 55286 57692 55298 57726
rect 55102 57686 55298 57692
rect 55796 57726 55992 57732
rect 55796 57692 55808 57726
rect 55980 57692 55992 57726
rect 55796 57686 55992 57692
rect 56490 57726 56686 57732
rect 56490 57692 56502 57726
rect 56674 57692 56686 57726
rect 56490 57686 56686 57692
rect 57184 57726 57380 57732
rect 57184 57692 57196 57726
rect 57368 57692 57380 57726
rect 57184 57686 57380 57692
rect 23622 57480 23818 57486
rect 23622 57446 23634 57480
rect 23806 57446 23818 57480
rect 23622 57440 23818 57446
rect 24316 57480 24512 57486
rect 24316 57446 24328 57480
rect 24500 57446 24512 57480
rect 24316 57440 24512 57446
rect 25010 57480 25206 57486
rect 25010 57446 25022 57480
rect 25194 57446 25206 57480
rect 25010 57440 25206 57446
rect 25704 57480 25900 57486
rect 25704 57446 25716 57480
rect 25888 57446 25900 57480
rect 25704 57440 25900 57446
rect 26398 57480 26594 57486
rect 26398 57446 26410 57480
rect 26582 57446 26594 57480
rect 26398 57440 26594 57446
rect 27092 57480 27288 57486
rect 27092 57446 27104 57480
rect 27276 57446 27288 57480
rect 27092 57440 27288 57446
rect 27786 57480 27982 57486
rect 27786 57446 27798 57480
rect 27970 57446 27982 57480
rect 27786 57440 27982 57446
rect 28480 57480 28676 57486
rect 28480 57446 28492 57480
rect 28664 57446 28676 57480
rect 28480 57440 28676 57446
rect 29174 57480 29370 57486
rect 29174 57446 29186 57480
rect 29358 57446 29370 57480
rect 29174 57440 29370 57446
rect 29868 57480 30064 57486
rect 29868 57446 29880 57480
rect 30052 57446 30064 57480
rect 29868 57440 30064 57446
rect 19532 57378 19728 57384
rect 19532 57344 19544 57378
rect 19716 57344 19728 57378
rect 926 57328 1122 57334
rect 926 57294 938 57328
rect 1110 57294 1122 57328
rect 926 57288 1122 57294
rect 1620 57328 1816 57334
rect 1620 57294 1632 57328
rect 1804 57294 1816 57328
rect 1620 57288 1816 57294
rect 2314 57328 2510 57334
rect 6268 57330 6464 57336
rect 2314 57294 2326 57328
rect 2498 57294 2510 57328
rect 2314 57288 2510 57294
rect 3594 57324 3790 57330
rect 3594 57290 3606 57324
rect 3778 57290 3790 57324
rect 3594 57284 3790 57290
rect 4288 57324 4484 57330
rect 4288 57290 4300 57324
rect 4472 57290 4484 57324
rect 4288 57284 4484 57290
rect 4982 57324 5178 57330
rect 4982 57290 4994 57324
rect 5166 57290 5178 57324
rect 6268 57296 6280 57330
rect 6452 57296 6464 57330
rect 6268 57290 6464 57296
rect 6962 57330 7158 57336
rect 6962 57296 6974 57330
rect 7146 57296 7158 57330
rect 6962 57290 7158 57296
rect 7656 57330 7852 57336
rect 7656 57296 7668 57330
rect 7840 57296 7852 57330
rect 7656 57290 7852 57296
rect 8914 57330 9110 57336
rect 8914 57296 8926 57330
rect 9098 57296 9110 57330
rect 8914 57290 9110 57296
rect 9608 57330 9804 57336
rect 9608 57296 9620 57330
rect 9792 57296 9804 57330
rect 9608 57290 9804 57296
rect 10302 57330 10498 57336
rect 14222 57330 14418 57336
rect 10302 57296 10314 57330
rect 10486 57296 10498 57330
rect 10302 57290 10498 57296
rect 11568 57324 11764 57330
rect 11568 57290 11580 57324
rect 11752 57290 11764 57324
rect 4982 57284 5178 57290
rect 11568 57284 11764 57290
rect 12262 57324 12458 57330
rect 12262 57290 12274 57324
rect 12446 57290 12458 57324
rect 12262 57284 12458 57290
rect 12956 57324 13152 57330
rect 12956 57290 12968 57324
rect 13140 57290 13152 57324
rect 14222 57296 14234 57330
rect 14406 57296 14418 57330
rect 14222 57290 14418 57296
rect 14916 57330 15112 57336
rect 14916 57296 14928 57330
rect 15100 57296 15112 57330
rect 14916 57290 15112 57296
rect 15610 57330 15806 57336
rect 15610 57296 15622 57330
rect 15794 57296 15806 57330
rect 15610 57290 15806 57296
rect 16848 57334 17044 57340
rect 16848 57300 16860 57334
rect 17032 57300 17044 57334
rect 16848 57294 17044 57300
rect 17542 57334 17738 57340
rect 17542 57300 17554 57334
rect 17726 57300 17738 57334
rect 17542 57294 17738 57300
rect 18236 57334 18432 57340
rect 19532 57338 19728 57344
rect 20226 57378 20422 57384
rect 20226 57344 20238 57378
rect 20410 57344 20422 57378
rect 20226 57338 20422 57344
rect 18236 57300 18248 57334
rect 18420 57300 18432 57334
rect 18236 57294 18432 57300
rect 12956 57284 13152 57290
rect 58862 57288 59190 57300
rect 42370 57068 42566 57074
rect 42370 57034 42382 57068
rect 42554 57034 42566 57068
rect 42370 57028 42566 57034
rect 43064 57068 43260 57074
rect 43064 57034 43076 57068
rect 43248 57034 43260 57068
rect 43064 57028 43260 57034
rect 43758 57068 43954 57074
rect 43758 57034 43770 57068
rect 43942 57034 43954 57068
rect 43758 57028 43954 57034
rect 44452 57068 44648 57074
rect 44452 57034 44464 57068
rect 44636 57034 44648 57068
rect 44452 57028 44648 57034
rect 45146 57068 45342 57074
rect 45146 57034 45158 57068
rect 45330 57034 45342 57068
rect 45146 57028 45342 57034
rect 46364 57068 46560 57074
rect 46364 57034 46376 57068
rect 46548 57034 46560 57068
rect 46364 57028 46560 57034
rect 47058 57068 47254 57074
rect 47058 57034 47070 57068
rect 47242 57034 47254 57068
rect 47058 57028 47254 57034
rect 47752 57068 47948 57074
rect 47752 57034 47764 57068
rect 47936 57034 47948 57068
rect 47752 57028 47948 57034
rect 48446 57068 48642 57074
rect 48446 57034 48458 57068
rect 48630 57034 48642 57068
rect 48446 57028 48642 57034
rect 49140 57068 49336 57074
rect 49140 57034 49152 57068
rect 49324 57034 49336 57068
rect 49140 57028 49336 57034
rect 50386 57068 50582 57074
rect 50386 57034 50398 57068
rect 50570 57034 50582 57068
rect 50386 57028 50582 57034
rect 51080 57068 51276 57074
rect 51080 57034 51092 57068
rect 51264 57034 51276 57068
rect 51080 57028 51276 57034
rect 51774 57068 51970 57074
rect 51774 57034 51786 57068
rect 51958 57034 51970 57068
rect 51774 57028 51970 57034
rect 52468 57068 52664 57074
rect 52468 57034 52480 57068
rect 52652 57034 52664 57068
rect 52468 57028 52664 57034
rect 53162 57068 53358 57074
rect 53162 57034 53174 57068
rect 53346 57034 53358 57068
rect 53162 57028 53358 57034
rect 54408 57068 54604 57074
rect 54408 57034 54420 57068
rect 54592 57034 54604 57068
rect 54408 57028 54604 57034
rect 55102 57068 55298 57074
rect 55102 57034 55114 57068
rect 55286 57034 55298 57068
rect 55102 57028 55298 57034
rect 55796 57068 55992 57074
rect 55796 57034 55808 57068
rect 55980 57034 55992 57068
rect 55796 57028 55992 57034
rect 56490 57068 56686 57074
rect 56490 57034 56502 57068
rect 56674 57034 56686 57068
rect 56490 57028 56686 57034
rect 57184 57068 57380 57074
rect 57184 57034 57196 57068
rect 57368 57034 57380 57068
rect 57184 57028 57380 57034
rect 30322 56840 30416 56870
rect 23622 56822 23818 56828
rect 23622 56788 23634 56822
rect 23806 56788 23818 56822
rect 23622 56782 23818 56788
rect 24316 56822 24512 56828
rect 24316 56788 24328 56822
rect 24500 56788 24512 56822
rect 24316 56782 24512 56788
rect 25010 56822 25206 56828
rect 25010 56788 25022 56822
rect 25194 56788 25206 56822
rect 25010 56782 25206 56788
rect 25704 56822 25900 56828
rect 25704 56788 25716 56822
rect 25888 56788 25900 56822
rect 25704 56782 25900 56788
rect 26398 56822 26594 56828
rect 26398 56788 26410 56822
rect 26582 56788 26594 56822
rect 26398 56782 26594 56788
rect 27092 56822 27288 56828
rect 27092 56788 27104 56822
rect 27276 56788 27288 56822
rect 27092 56782 27288 56788
rect 27786 56822 27982 56828
rect 27786 56788 27798 56822
rect 27970 56788 27982 56822
rect 27786 56782 27982 56788
rect 28480 56822 28676 56828
rect 28480 56788 28492 56822
rect 28664 56788 28676 56822
rect 28480 56782 28676 56788
rect 29174 56822 29370 56828
rect 29174 56788 29186 56822
rect 29358 56788 29370 56822
rect 29174 56782 29370 56788
rect 29868 56822 30064 56828
rect 29868 56788 29880 56822
rect 30052 56788 30064 56822
rect 29868 56782 30064 56788
rect 30322 56782 30348 56840
rect 30386 56782 30416 56840
rect 58862 56840 58868 57288
rect 59184 57078 59190 57288
rect 59226 57078 59236 57262
rect 59184 56938 59236 57078
rect 59184 56840 59190 56938
rect 59226 56850 59236 56938
rect 59510 56850 59520 57262
rect 58862 56828 59190 56840
rect 222 56552 554 56766
rect 30322 56750 30416 56782
rect 19532 56720 19728 56726
rect 19532 56686 19544 56720
rect 19716 56686 19728 56720
rect 926 56670 1122 56676
rect 926 56636 938 56670
rect 1110 56636 1122 56670
rect 926 56630 1122 56636
rect 1620 56670 1816 56676
rect 1620 56636 1632 56670
rect 1804 56636 1816 56670
rect 1620 56630 1816 56636
rect 2314 56670 2510 56676
rect 6268 56672 6464 56678
rect 2314 56636 2326 56670
rect 2498 56636 2510 56670
rect 2314 56630 2510 56636
rect 3594 56666 3790 56672
rect 3594 56632 3606 56666
rect 3778 56632 3790 56666
rect 3594 56626 3790 56632
rect 4288 56666 4484 56672
rect 4288 56632 4300 56666
rect 4472 56632 4484 56666
rect 4288 56626 4484 56632
rect 4982 56666 5178 56672
rect 4982 56632 4994 56666
rect 5166 56632 5178 56666
rect 6268 56638 6280 56672
rect 6452 56638 6464 56672
rect 6268 56632 6464 56638
rect 6962 56672 7158 56678
rect 6962 56638 6974 56672
rect 7146 56638 7158 56672
rect 6962 56632 7158 56638
rect 7656 56672 7852 56678
rect 7656 56638 7668 56672
rect 7840 56638 7852 56672
rect 7656 56632 7852 56638
rect 8914 56672 9110 56678
rect 8914 56638 8926 56672
rect 9098 56638 9110 56672
rect 8914 56632 9110 56638
rect 9608 56672 9804 56678
rect 9608 56638 9620 56672
rect 9792 56638 9804 56672
rect 9608 56632 9804 56638
rect 10302 56672 10498 56678
rect 14222 56672 14418 56678
rect 10302 56638 10314 56672
rect 10486 56638 10498 56672
rect 10302 56632 10498 56638
rect 11568 56666 11764 56672
rect 11568 56632 11580 56666
rect 11752 56632 11764 56666
rect 4982 56626 5178 56632
rect 11568 56626 11764 56632
rect 12262 56666 12458 56672
rect 12262 56632 12274 56666
rect 12446 56632 12458 56666
rect 12262 56626 12458 56632
rect 12956 56666 13152 56672
rect 12956 56632 12968 56666
rect 13140 56632 13152 56666
rect 14222 56638 14234 56672
rect 14406 56638 14418 56672
rect 14222 56632 14418 56638
rect 14916 56672 15112 56678
rect 14916 56638 14928 56672
rect 15100 56638 15112 56672
rect 14916 56632 15112 56638
rect 15610 56672 15806 56678
rect 15610 56638 15622 56672
rect 15794 56638 15806 56672
rect 15610 56632 15806 56638
rect 16848 56676 17044 56682
rect 16848 56642 16860 56676
rect 17032 56642 17044 56676
rect 16848 56636 17044 56642
rect 17542 56676 17738 56682
rect 17542 56642 17554 56676
rect 17726 56642 17738 56676
rect 17542 56636 17738 56642
rect 18236 56676 18432 56682
rect 19532 56680 19728 56686
rect 20226 56720 20422 56726
rect 20226 56686 20238 56720
rect 20410 56686 20422 56720
rect 20226 56680 20422 56686
rect 18236 56642 18248 56676
rect 18420 56642 18432 56676
rect 18236 56636 18432 56642
rect 12956 56626 13152 56632
rect 42678 56420 45324 56508
rect 42678 56218 42976 56420
rect 45150 56218 45324 56420
rect 23622 56164 23818 56170
rect 23622 56130 23634 56164
rect 23806 56130 23818 56164
rect 23622 56124 23818 56130
rect 24316 56164 24512 56170
rect 24316 56130 24328 56164
rect 24500 56130 24512 56164
rect 24316 56124 24512 56130
rect 25010 56164 25206 56170
rect 25010 56130 25022 56164
rect 25194 56130 25206 56164
rect 25010 56124 25206 56130
rect 25704 56164 25900 56170
rect 25704 56130 25716 56164
rect 25888 56130 25900 56164
rect 25704 56124 25900 56130
rect 26398 56164 26594 56170
rect 26398 56130 26410 56164
rect 26582 56130 26594 56164
rect 26398 56124 26594 56130
rect 27092 56164 27288 56170
rect 27092 56130 27104 56164
rect 27276 56130 27288 56164
rect 27092 56124 27288 56130
rect 27786 56164 27982 56170
rect 27786 56130 27798 56164
rect 27970 56130 27982 56164
rect 27786 56124 27982 56130
rect 28480 56164 28676 56170
rect 28480 56130 28492 56164
rect 28664 56130 28676 56164
rect 28480 56124 28676 56130
rect 29174 56164 29370 56170
rect 29174 56130 29186 56164
rect 29358 56130 29370 56164
rect 29174 56124 29370 56130
rect 29868 56164 30064 56170
rect 29868 56130 29880 56164
rect 30052 56130 30064 56164
rect 29868 56124 30064 56130
rect 42678 56106 45324 56218
rect 46686 56418 49332 56506
rect 46686 56216 46984 56418
rect 49158 56216 49332 56418
rect 46686 56104 49332 56216
rect 50698 56418 53344 56506
rect 50698 56216 50996 56418
rect 53170 56216 53344 56418
rect 50698 56104 53344 56216
rect 54708 56418 57354 56506
rect 54708 56216 55006 56418
rect 57180 56216 57354 56418
rect 54708 56104 57354 56216
rect 19532 56062 19728 56068
rect 19532 56028 19544 56062
rect 19716 56028 19728 56062
rect 926 56012 1122 56018
rect 926 55978 938 56012
rect 1110 55978 1122 56012
rect 926 55972 1122 55978
rect 1620 56012 1816 56018
rect 1620 55978 1632 56012
rect 1804 55978 1816 56012
rect 1620 55972 1816 55978
rect 2314 56012 2510 56018
rect 6268 56014 6464 56020
rect 2314 55978 2326 56012
rect 2498 55978 2510 56012
rect 2314 55972 2510 55978
rect 3594 56008 3790 56014
rect 3594 55974 3606 56008
rect 3778 55974 3790 56008
rect 3594 55968 3790 55974
rect 4288 56008 4484 56014
rect 4288 55974 4300 56008
rect 4472 55974 4484 56008
rect 4288 55968 4484 55974
rect 4982 56008 5178 56014
rect 4982 55974 4994 56008
rect 5166 55974 5178 56008
rect 6268 55980 6280 56014
rect 6452 55980 6464 56014
rect 6268 55974 6464 55980
rect 6962 56014 7158 56020
rect 6962 55980 6974 56014
rect 7146 55980 7158 56014
rect 6962 55974 7158 55980
rect 7656 56014 7852 56020
rect 7656 55980 7668 56014
rect 7840 55980 7852 56014
rect 7656 55974 7852 55980
rect 8914 56014 9110 56020
rect 8914 55980 8926 56014
rect 9098 55980 9110 56014
rect 8914 55974 9110 55980
rect 9608 56014 9804 56020
rect 9608 55980 9620 56014
rect 9792 55980 9804 56014
rect 9608 55974 9804 55980
rect 10302 56014 10498 56020
rect 14222 56014 14418 56020
rect 10302 55980 10314 56014
rect 10486 55980 10498 56014
rect 10302 55974 10498 55980
rect 11568 56008 11764 56014
rect 11568 55974 11580 56008
rect 11752 55974 11764 56008
rect 4982 55968 5178 55974
rect 11568 55968 11764 55974
rect 12262 56008 12458 56014
rect 12262 55974 12274 56008
rect 12446 55974 12458 56008
rect 12262 55968 12458 55974
rect 12956 56008 13152 56014
rect 12956 55974 12968 56008
rect 13140 55974 13152 56008
rect 14222 55980 14234 56014
rect 14406 55980 14418 56014
rect 14222 55974 14418 55980
rect 14916 56014 15112 56020
rect 14916 55980 14928 56014
rect 15100 55980 15112 56014
rect 14916 55974 15112 55980
rect 15610 56014 15806 56020
rect 15610 55980 15622 56014
rect 15794 55980 15806 56014
rect 15610 55974 15806 55980
rect 16848 56018 17044 56024
rect 16848 55984 16860 56018
rect 17032 55984 17044 56018
rect 16848 55978 17044 55984
rect 17542 56018 17738 56024
rect 17542 55984 17554 56018
rect 17726 55984 17738 56018
rect 17542 55978 17738 55984
rect 18236 56018 18432 56024
rect 19532 56022 19728 56028
rect 20226 56062 20422 56068
rect 20226 56028 20238 56062
rect 20410 56028 20422 56062
rect 20226 56022 20422 56028
rect 18236 55984 18248 56018
rect 18420 55984 18432 56018
rect 18236 55978 18432 55984
rect 12956 55968 13152 55974
rect 28686 55946 29576 55990
rect 24274 55844 25162 55908
rect 28686 55902 28824 55946
rect 29468 55902 29576 55946
rect 42322 55968 42518 55974
rect 42322 55934 42334 55968
rect 42506 55934 42518 55968
rect 42322 55928 42518 55934
rect 43016 55968 43212 55974
rect 43016 55934 43028 55968
rect 43200 55934 43212 55968
rect 43016 55928 43212 55934
rect 43710 55968 43906 55974
rect 43710 55934 43722 55968
rect 43894 55934 43906 55968
rect 43710 55928 43906 55934
rect 44404 55968 44600 55974
rect 44404 55934 44416 55968
rect 44588 55934 44600 55968
rect 44404 55928 44600 55934
rect 45098 55968 45294 55974
rect 45098 55934 45110 55968
rect 45282 55934 45294 55968
rect 45098 55928 45294 55934
rect 46330 55966 46526 55972
rect 46330 55932 46342 55966
rect 46514 55932 46526 55966
rect 46330 55926 46526 55932
rect 47024 55966 47220 55972
rect 47024 55932 47036 55966
rect 47208 55932 47220 55966
rect 47024 55926 47220 55932
rect 47718 55966 47914 55972
rect 47718 55932 47730 55966
rect 47902 55932 47914 55966
rect 47718 55926 47914 55932
rect 48412 55966 48608 55972
rect 48412 55932 48424 55966
rect 48596 55932 48608 55966
rect 48412 55926 48608 55932
rect 49106 55966 49302 55972
rect 49106 55932 49118 55966
rect 49290 55932 49302 55966
rect 49106 55926 49302 55932
rect 50342 55966 50538 55972
rect 50342 55932 50354 55966
rect 50526 55932 50538 55966
rect 50342 55926 50538 55932
rect 51036 55966 51232 55972
rect 51036 55932 51048 55966
rect 51220 55932 51232 55966
rect 51036 55926 51232 55932
rect 51730 55966 51926 55972
rect 51730 55932 51742 55966
rect 51914 55932 51926 55966
rect 51730 55926 51926 55932
rect 52424 55966 52620 55972
rect 52424 55932 52436 55966
rect 52608 55932 52620 55966
rect 52424 55926 52620 55932
rect 53118 55966 53314 55972
rect 53118 55932 53130 55966
rect 53302 55932 53314 55966
rect 53118 55926 53314 55932
rect 54352 55966 54548 55972
rect 54352 55932 54364 55966
rect 54536 55932 54548 55966
rect 54352 55926 54548 55932
rect 55046 55966 55242 55972
rect 55046 55932 55058 55966
rect 55230 55932 55242 55966
rect 55046 55926 55242 55932
rect 55740 55966 55936 55972
rect 55740 55932 55752 55966
rect 55924 55932 55936 55966
rect 55740 55926 55936 55932
rect 56434 55966 56630 55972
rect 56434 55932 56446 55966
rect 56618 55932 56630 55966
rect 56434 55926 56630 55932
rect 57128 55966 57324 55972
rect 57128 55932 57140 55966
rect 57312 55932 57324 55966
rect 57128 55926 57324 55932
rect 28686 55848 29576 55902
rect 24274 55788 24408 55844
rect 25052 55788 25162 55844
rect 24274 55732 25162 55788
rect 30970 55602 30980 55738
rect 29968 55596 30980 55602
rect 23628 55590 23824 55596
rect 23628 55556 23640 55590
rect 23812 55556 23824 55590
rect 23628 55550 23824 55556
rect 24322 55590 24518 55596
rect 24322 55556 24334 55590
rect 24506 55556 24518 55590
rect 24322 55550 24518 55556
rect 25016 55590 25212 55596
rect 25016 55556 25028 55590
rect 25200 55556 25212 55590
rect 25016 55550 25212 55556
rect 25710 55590 25906 55596
rect 25710 55556 25722 55590
rect 25894 55556 25906 55590
rect 25710 55550 25906 55556
rect 26404 55590 26600 55596
rect 26404 55556 26416 55590
rect 26588 55556 26600 55590
rect 26404 55550 26600 55556
rect 27098 55590 27294 55596
rect 27098 55556 27110 55590
rect 27282 55556 27294 55590
rect 27098 55550 27294 55556
rect 27792 55590 27988 55596
rect 27792 55556 27804 55590
rect 27976 55556 27988 55590
rect 27792 55550 27988 55556
rect 28486 55590 28682 55596
rect 28486 55556 28498 55590
rect 28670 55556 28682 55590
rect 28486 55550 28682 55556
rect 29180 55590 29376 55596
rect 29180 55556 29192 55590
rect 29364 55556 29376 55590
rect 29180 55550 29376 55556
rect 29874 55590 30980 55596
rect 29874 55556 29886 55590
rect 30058 55556 30980 55590
rect 29874 55550 30980 55556
rect 29968 55538 30980 55550
rect 30970 55430 30980 55538
rect 31268 55430 31278 55738
rect 19532 55404 19728 55410
rect 19532 55370 19544 55404
rect 19716 55370 19728 55404
rect 926 55354 1122 55360
rect 926 55320 938 55354
rect 1110 55320 1122 55354
rect 926 55314 1122 55320
rect 1620 55354 1816 55360
rect 1620 55320 1632 55354
rect 1804 55320 1816 55354
rect 1620 55314 1816 55320
rect 2314 55354 2510 55360
rect 6268 55356 6464 55362
rect 2314 55320 2326 55354
rect 2498 55320 2510 55354
rect 2314 55314 2510 55320
rect 3594 55350 3790 55356
rect 3594 55316 3606 55350
rect 3778 55316 3790 55350
rect 3594 55310 3790 55316
rect 4288 55350 4484 55356
rect 4288 55316 4300 55350
rect 4472 55316 4484 55350
rect 4288 55310 4484 55316
rect 4982 55350 5178 55356
rect 4982 55316 4994 55350
rect 5166 55316 5178 55350
rect 6268 55322 6280 55356
rect 6452 55322 6464 55356
rect 6268 55316 6464 55322
rect 6962 55356 7158 55362
rect 6962 55322 6974 55356
rect 7146 55322 7158 55356
rect 6962 55316 7158 55322
rect 7656 55356 7852 55362
rect 7656 55322 7668 55356
rect 7840 55322 7852 55356
rect 7656 55316 7852 55322
rect 8914 55356 9110 55362
rect 8914 55322 8926 55356
rect 9098 55322 9110 55356
rect 8914 55316 9110 55322
rect 9608 55356 9804 55362
rect 9608 55322 9620 55356
rect 9792 55322 9804 55356
rect 9608 55316 9804 55322
rect 10302 55356 10498 55362
rect 14222 55356 14418 55362
rect 10302 55322 10314 55356
rect 10486 55322 10498 55356
rect 10302 55316 10498 55322
rect 11568 55350 11764 55356
rect 11568 55316 11580 55350
rect 11752 55316 11764 55350
rect 4982 55310 5178 55316
rect 11568 55310 11764 55316
rect 12262 55350 12458 55356
rect 12262 55316 12274 55350
rect 12446 55316 12458 55350
rect 12262 55310 12458 55316
rect 12956 55350 13152 55356
rect 12956 55316 12968 55350
rect 13140 55316 13152 55350
rect 14222 55322 14234 55356
rect 14406 55322 14418 55356
rect 14222 55316 14418 55322
rect 14916 55356 15112 55362
rect 14916 55322 14928 55356
rect 15100 55322 15112 55356
rect 14916 55316 15112 55322
rect 15610 55356 15806 55362
rect 15610 55322 15622 55356
rect 15794 55322 15806 55356
rect 15610 55316 15806 55322
rect 16848 55360 17044 55366
rect 16848 55326 16860 55360
rect 17032 55326 17044 55360
rect 16848 55320 17044 55326
rect 17542 55360 17738 55366
rect 17542 55326 17554 55360
rect 17726 55326 17738 55360
rect 17542 55320 17738 55326
rect 18236 55360 18432 55366
rect 19532 55364 19728 55370
rect 20226 55404 20422 55410
rect 20226 55370 20238 55404
rect 20410 55370 20422 55404
rect 20226 55364 20422 55370
rect 18236 55326 18248 55360
rect 18420 55326 18432 55360
rect 18236 55320 18432 55326
rect 22916 55346 23202 55376
rect 12956 55310 13152 55316
rect 22916 55000 23006 55346
rect 23088 55000 23202 55346
rect 42322 55310 42518 55316
rect 42322 55276 42334 55310
rect 42506 55276 42518 55310
rect 42322 55270 42518 55276
rect 43016 55310 43212 55316
rect 43016 55276 43028 55310
rect 43200 55276 43212 55310
rect 43016 55270 43212 55276
rect 43710 55310 43906 55316
rect 43710 55276 43722 55310
rect 43894 55276 43906 55310
rect 43710 55270 43906 55276
rect 44404 55310 44600 55316
rect 44404 55276 44416 55310
rect 44588 55276 44600 55310
rect 44404 55270 44600 55276
rect 45098 55310 45294 55316
rect 45098 55276 45110 55310
rect 45282 55276 45294 55310
rect 45098 55270 45294 55276
rect 46330 55308 46526 55314
rect 46330 55274 46342 55308
rect 46514 55274 46526 55308
rect 46330 55268 46526 55274
rect 47024 55308 47220 55314
rect 47024 55274 47036 55308
rect 47208 55274 47220 55308
rect 47024 55268 47220 55274
rect 47718 55308 47914 55314
rect 47718 55274 47730 55308
rect 47902 55274 47914 55308
rect 47718 55268 47914 55274
rect 48412 55308 48608 55314
rect 48412 55274 48424 55308
rect 48596 55274 48608 55308
rect 48412 55268 48608 55274
rect 49106 55308 49302 55314
rect 49106 55274 49118 55308
rect 49290 55274 49302 55308
rect 49106 55268 49302 55274
rect 50342 55308 50538 55314
rect 50342 55274 50354 55308
rect 50526 55274 50538 55308
rect 50342 55268 50538 55274
rect 51036 55308 51232 55314
rect 51036 55274 51048 55308
rect 51220 55274 51232 55308
rect 51036 55268 51232 55274
rect 51730 55308 51926 55314
rect 51730 55274 51742 55308
rect 51914 55274 51926 55308
rect 51730 55268 51926 55274
rect 52424 55308 52620 55314
rect 52424 55274 52436 55308
rect 52608 55274 52620 55308
rect 52424 55268 52620 55274
rect 53118 55308 53314 55314
rect 53118 55274 53130 55308
rect 53302 55274 53314 55308
rect 53118 55268 53314 55274
rect 54352 55308 54548 55314
rect 54352 55274 54364 55308
rect 54536 55274 54548 55308
rect 54352 55268 54548 55274
rect 55046 55308 55242 55314
rect 55046 55274 55058 55308
rect 55230 55274 55242 55308
rect 55046 55268 55242 55274
rect 55740 55308 55936 55314
rect 55740 55274 55752 55308
rect 55924 55274 55936 55308
rect 55740 55268 55936 55274
rect 56434 55308 56630 55314
rect 56434 55274 56446 55308
rect 56618 55274 56630 55308
rect 56434 55268 56630 55274
rect 57128 55308 57324 55314
rect 57128 55274 57140 55308
rect 57312 55274 57324 55308
rect 57128 55268 57324 55274
rect 8346 54912 8560 54924
rect 5686 54836 5934 54848
rect 3052 54802 3282 54814
rect 3052 54752 3058 54802
rect 2368 54702 3058 54752
rect 926 54696 1122 54702
rect 926 54662 938 54696
rect 1110 54662 1122 54696
rect 926 54656 1122 54662
rect 1620 54696 1816 54702
rect 1620 54662 1632 54696
rect 1804 54662 1816 54696
rect 1620 54656 1816 54662
rect 2314 54696 3058 54702
rect 2314 54662 2326 54696
rect 2498 54662 3058 54696
rect 2314 54656 3058 54662
rect 2368 54592 3058 54656
rect 3052 54448 3058 54592
rect 3276 54448 3282 54802
rect 5686 54752 5692 54836
rect 5078 54698 5692 54752
rect 3594 54692 3790 54698
rect 3594 54658 3606 54692
rect 3778 54658 3790 54692
rect 3594 54652 3790 54658
rect 4288 54692 4484 54698
rect 4288 54658 4300 54692
rect 4472 54658 4484 54692
rect 4288 54652 4484 54658
rect 4982 54692 5692 54698
rect 4982 54658 4994 54692
rect 5166 54658 5692 54692
rect 4982 54652 5692 54658
rect 5078 54584 5692 54652
rect 5686 54474 5692 54584
rect 5928 54474 5934 54836
rect 8346 54794 8352 54912
rect 7720 54704 8352 54794
rect 6268 54698 6464 54704
rect 6268 54664 6280 54698
rect 6452 54664 6464 54698
rect 6268 54658 6464 54664
rect 6962 54698 7158 54704
rect 6962 54664 6974 54698
rect 7146 54664 7158 54698
rect 6962 54658 7158 54664
rect 7656 54698 8352 54704
rect 7656 54664 7668 54698
rect 7840 54664 8352 54698
rect 7656 54658 8352 54664
rect 7720 54558 8352 54658
rect 5686 54462 5934 54474
rect 3052 54436 3282 54448
rect 8346 54424 8352 54558
rect 8554 54424 8560 54912
rect 18838 54894 19060 54906
rect 13672 54860 13852 54872
rect 11022 54828 11252 54840
rect 11022 54742 11028 54828
rect 10380 54704 11028 54742
rect 8914 54698 9110 54704
rect 8914 54664 8926 54698
rect 9098 54664 9110 54698
rect 8914 54658 9110 54664
rect 9608 54698 9804 54704
rect 9608 54664 9620 54698
rect 9792 54664 9804 54698
rect 9608 54658 9804 54664
rect 10302 54698 11028 54704
rect 10302 54664 10314 54698
rect 10486 54664 11028 54698
rect 10302 54658 11028 54664
rect 10380 54550 11028 54658
rect 8346 54412 8560 54424
rect 11022 54390 11028 54550
rect 11246 54390 11252 54828
rect 13672 54734 13678 54860
rect 12988 54698 13678 54734
rect 11568 54692 11764 54698
rect 11568 54658 11580 54692
rect 11752 54658 11764 54692
rect 11568 54652 11764 54658
rect 12262 54692 12458 54698
rect 12262 54658 12274 54692
rect 12446 54658 12458 54692
rect 12262 54652 12458 54658
rect 12956 54692 13678 54698
rect 12956 54658 12968 54692
rect 13140 54658 13678 54692
rect 12956 54652 13678 54658
rect 12988 54616 13678 54652
rect 13672 54432 13678 54616
rect 13846 54432 13852 54860
rect 16288 54802 16554 54814
rect 16288 54760 16294 54802
rect 15664 54704 16294 54760
rect 14222 54698 14418 54704
rect 14222 54664 14234 54698
rect 14406 54664 14418 54698
rect 14222 54658 14418 54664
rect 14916 54698 15112 54704
rect 14916 54664 14928 54698
rect 15100 54664 15112 54698
rect 14916 54658 15112 54664
rect 15610 54698 16294 54704
rect 15610 54664 15622 54698
rect 15794 54664 16294 54698
rect 15610 54658 16294 54664
rect 15664 54642 16294 54658
rect 16288 54532 16294 54642
rect 16548 54532 16554 54802
rect 18838 54784 18844 54894
rect 18290 54708 18844 54784
rect 16848 54702 17044 54708
rect 16848 54668 16860 54702
rect 17032 54668 17044 54702
rect 16848 54662 17044 54668
rect 17542 54702 17738 54708
rect 17542 54668 17554 54702
rect 17726 54668 17738 54702
rect 17542 54662 17738 54668
rect 18236 54702 18844 54708
rect 18236 54668 18248 54702
rect 18420 54668 18844 54702
rect 18236 54662 18844 54668
rect 18290 54626 18844 54662
rect 16288 54520 16554 54532
rect 18716 54548 18844 54626
rect 19054 54548 19060 54894
rect 22916 54860 23202 55000
rect 23628 54932 23824 54938
rect 23628 54898 23640 54932
rect 23812 54898 23824 54932
rect 23628 54892 23824 54898
rect 24322 54932 24518 54938
rect 24322 54898 24334 54932
rect 24506 54898 24518 54932
rect 24322 54892 24518 54898
rect 25016 54932 25212 54938
rect 25016 54898 25028 54932
rect 25200 54898 25212 54932
rect 25016 54892 25212 54898
rect 25710 54932 25906 54938
rect 25710 54898 25722 54932
rect 25894 54898 25906 54932
rect 25710 54892 25906 54898
rect 26404 54932 26600 54938
rect 26404 54898 26416 54932
rect 26588 54898 26600 54932
rect 26404 54892 26600 54898
rect 27098 54932 27294 54938
rect 27098 54898 27110 54932
rect 27282 54898 27294 54932
rect 27098 54892 27294 54898
rect 27792 54932 27988 54938
rect 27792 54898 27804 54932
rect 27976 54898 27988 54932
rect 27792 54892 27988 54898
rect 28486 54932 28682 54938
rect 28486 54898 28498 54932
rect 28670 54898 28682 54932
rect 28486 54892 28682 54898
rect 29180 54932 29376 54938
rect 29180 54898 29192 54932
rect 29364 54898 29376 54932
rect 29180 54892 29376 54898
rect 29874 54932 30070 54938
rect 29874 54898 29886 54932
rect 30058 54898 30070 54932
rect 29874 54892 30070 54898
rect 19532 54746 19728 54752
rect 19532 54712 19544 54746
rect 19716 54712 19728 54746
rect 19532 54706 19728 54712
rect 20226 54746 20422 54752
rect 20226 54712 20238 54746
rect 20410 54712 20422 54746
rect 20226 54706 20422 54712
rect 23278 54720 23414 54780
rect 18716 54536 19060 54548
rect 20658 54628 20824 54672
rect 21354 54628 21608 54638
rect 23278 54628 23316 54720
rect 20658 54624 23316 54628
rect 13672 54420 13852 54432
rect 11022 54378 11252 54390
rect 926 54038 1122 54044
rect 926 54004 938 54038
rect 1110 54004 1122 54038
rect 926 53998 1122 54004
rect 1620 54038 1816 54044
rect 1620 54004 1632 54038
rect 1804 54004 1816 54038
rect 1620 53998 1816 54004
rect 2314 54038 2510 54044
rect 6268 54040 6464 54046
rect 2314 54004 2326 54038
rect 2498 54004 2510 54038
rect 2314 53998 2510 54004
rect 3594 54034 3790 54040
rect 3594 54000 3606 54034
rect 3778 54000 3790 54034
rect 3594 53994 3790 54000
rect 4288 54034 4484 54040
rect 4288 54000 4300 54034
rect 4472 54000 4484 54034
rect 4288 53994 4484 54000
rect 4982 54034 5178 54040
rect 4982 54000 4994 54034
rect 5166 54000 5178 54034
rect 6268 54006 6280 54040
rect 6452 54006 6464 54040
rect 6268 54000 6464 54006
rect 6962 54040 7158 54046
rect 6962 54006 6974 54040
rect 7146 54006 7158 54040
rect 6962 54000 7158 54006
rect 7656 54040 7852 54046
rect 7656 54006 7668 54040
rect 7840 54006 7852 54040
rect 7656 54000 7852 54006
rect 8914 54040 9110 54046
rect 8914 54006 8926 54040
rect 9098 54006 9110 54040
rect 8914 54000 9110 54006
rect 9608 54040 9804 54046
rect 9608 54006 9620 54040
rect 9792 54006 9804 54040
rect 9608 54000 9804 54006
rect 10302 54040 10498 54046
rect 14222 54040 14418 54046
rect 10302 54006 10314 54040
rect 10486 54006 10498 54040
rect 10302 54000 10498 54006
rect 11568 54034 11764 54040
rect 11568 54000 11580 54034
rect 11752 54000 11764 54034
rect 4982 53994 5178 54000
rect 11568 53994 11764 54000
rect 12262 54034 12458 54040
rect 12262 54000 12274 54034
rect 12446 54000 12458 54034
rect 12262 53994 12458 54000
rect 12956 54034 13152 54040
rect 12956 54000 12968 54034
rect 13140 54000 13152 54034
rect 14222 54006 14234 54040
rect 14406 54006 14418 54040
rect 14222 54000 14418 54006
rect 14916 54040 15112 54046
rect 14916 54006 14928 54040
rect 15100 54006 15112 54040
rect 14916 54000 15112 54006
rect 15610 54040 15806 54046
rect 15610 54006 15622 54040
rect 15794 54006 15806 54040
rect 15610 54000 15806 54006
rect 16848 54044 17044 54050
rect 16848 54010 16860 54044
rect 17032 54010 17044 54044
rect 16848 54004 17044 54010
rect 17542 54044 17738 54050
rect 17542 54010 17554 54044
rect 17726 54010 17738 54044
rect 17542 54004 17738 54010
rect 18236 54044 18432 54050
rect 18236 54010 18248 54044
rect 18420 54010 18432 54044
rect 18236 54004 18432 54010
rect 12956 53994 13152 54000
rect 18716 53726 18866 54536
rect 20658 54456 20690 54624
rect 20770 54504 23316 54624
rect 20770 54456 20824 54504
rect 20658 54392 20824 54456
rect 19532 54088 19728 54094
rect 19532 54054 19544 54088
rect 19716 54054 19728 54088
rect 19532 54048 19728 54054
rect 20226 54088 20422 54094
rect 20226 54054 20238 54088
rect 20410 54054 20422 54088
rect 20226 54048 20422 54054
rect 944 53270 2576 53328
rect 944 53200 1058 53270
rect 2462 53200 2576 53270
rect 944 53124 2576 53200
rect 3612 53266 5244 53324
rect 3612 53196 3726 53266
rect 5130 53196 5244 53266
rect 3612 53120 5244 53196
rect 6286 53272 7918 53330
rect 6286 53202 6400 53272
rect 7804 53202 7918 53272
rect 6286 53126 7918 53202
rect 8932 53272 10564 53330
rect 8932 53202 9046 53272
rect 10450 53202 10564 53272
rect 8932 53126 10564 53202
rect 11586 53266 13218 53324
rect 11586 53196 11700 53266
rect 13104 53196 13218 53266
rect 11586 53120 13218 53196
rect 14240 53272 15872 53330
rect 14240 53202 14354 53272
rect 15758 53202 15872 53272
rect 14240 53126 15872 53202
rect 16866 53276 18498 53334
rect 16866 53206 16980 53276
rect 18384 53206 18498 53276
rect 16866 53130 18498 53206
rect 19364 53290 20600 53360
rect 19364 53182 19534 53290
rect 20492 53182 20600 53290
rect 19364 53090 20600 53182
rect 19532 52986 19728 52992
rect 19532 52952 19544 52986
rect 19716 52952 19728 52986
rect 926 52936 1122 52942
rect 926 52902 938 52936
rect 1110 52902 1122 52936
rect 926 52896 1122 52902
rect 1620 52936 1816 52942
rect 1620 52902 1632 52936
rect 1804 52902 1816 52936
rect 1620 52896 1816 52902
rect 2314 52936 2510 52942
rect 6268 52938 6464 52944
rect 2314 52902 2326 52936
rect 2498 52902 2510 52936
rect 2314 52896 2510 52902
rect 3594 52932 3790 52938
rect 3594 52898 3606 52932
rect 3778 52898 3790 52932
rect 3594 52892 3790 52898
rect 4288 52932 4484 52938
rect 4288 52898 4300 52932
rect 4472 52898 4484 52932
rect 4288 52892 4484 52898
rect 4982 52932 5178 52938
rect 4982 52898 4994 52932
rect 5166 52898 5178 52932
rect 6268 52904 6280 52938
rect 6452 52904 6464 52938
rect 6268 52898 6464 52904
rect 6962 52938 7158 52944
rect 6962 52904 6974 52938
rect 7146 52904 7158 52938
rect 6962 52898 7158 52904
rect 7656 52938 7852 52944
rect 7656 52904 7668 52938
rect 7840 52904 7852 52938
rect 7656 52898 7852 52904
rect 8914 52938 9110 52944
rect 8914 52904 8926 52938
rect 9098 52904 9110 52938
rect 8914 52898 9110 52904
rect 9608 52938 9804 52944
rect 9608 52904 9620 52938
rect 9792 52904 9804 52938
rect 9608 52898 9804 52904
rect 10302 52938 10498 52944
rect 14222 52938 14418 52944
rect 10302 52904 10314 52938
rect 10486 52904 10498 52938
rect 10302 52898 10498 52904
rect 11568 52932 11764 52938
rect 11568 52898 11580 52932
rect 11752 52898 11764 52932
rect 4982 52892 5178 52898
rect 11568 52892 11764 52898
rect 12262 52932 12458 52938
rect 12262 52898 12274 52932
rect 12446 52898 12458 52932
rect 12262 52892 12458 52898
rect 12956 52932 13152 52938
rect 12956 52898 12968 52932
rect 13140 52898 13152 52932
rect 14222 52904 14234 52938
rect 14406 52904 14418 52938
rect 14222 52898 14418 52904
rect 14916 52938 15112 52944
rect 14916 52904 14928 52938
rect 15100 52904 15112 52938
rect 14916 52898 15112 52904
rect 15610 52938 15806 52944
rect 15610 52904 15622 52938
rect 15794 52904 15806 52938
rect 15610 52898 15806 52904
rect 16848 52942 17044 52948
rect 16848 52908 16860 52942
rect 17032 52908 17044 52942
rect 16848 52902 17044 52908
rect 17542 52942 17738 52948
rect 17542 52908 17554 52942
rect 17726 52908 17738 52942
rect 17542 52902 17738 52908
rect 18236 52942 18432 52948
rect 19532 52946 19728 52952
rect 20226 52986 20422 52992
rect 20226 52952 20238 52986
rect 20410 52952 20422 52986
rect 20226 52946 20422 52952
rect 18236 52908 18248 52942
rect 18420 52908 18432 52942
rect 18236 52902 18432 52908
rect 12956 52892 13152 52898
rect 19532 52328 19728 52334
rect 19532 52294 19544 52328
rect 19716 52294 19728 52328
rect 926 52278 1122 52284
rect 926 52244 938 52278
rect 1110 52244 1122 52278
rect 926 52238 1122 52244
rect 1620 52278 1816 52284
rect 1620 52244 1632 52278
rect 1804 52244 1816 52278
rect 1620 52238 1816 52244
rect 2314 52278 2510 52284
rect 6268 52280 6464 52286
rect 2314 52244 2326 52278
rect 2498 52244 2510 52278
rect 2314 52238 2510 52244
rect 3594 52274 3790 52280
rect 3594 52240 3606 52274
rect 3778 52240 3790 52274
rect 3594 52234 3790 52240
rect 4288 52274 4484 52280
rect 4288 52240 4300 52274
rect 4472 52240 4484 52274
rect 4288 52234 4484 52240
rect 4982 52274 5178 52280
rect 4982 52240 4994 52274
rect 5166 52240 5178 52274
rect 6268 52246 6280 52280
rect 6452 52246 6464 52280
rect 6268 52240 6464 52246
rect 6962 52280 7158 52286
rect 6962 52246 6974 52280
rect 7146 52246 7158 52280
rect 6962 52240 7158 52246
rect 7656 52280 7852 52286
rect 7656 52246 7668 52280
rect 7840 52246 7852 52280
rect 7656 52240 7852 52246
rect 8914 52280 9110 52286
rect 8914 52246 8926 52280
rect 9098 52246 9110 52280
rect 8914 52240 9110 52246
rect 9608 52280 9804 52286
rect 9608 52246 9620 52280
rect 9792 52246 9804 52280
rect 9608 52240 9804 52246
rect 10302 52280 10498 52286
rect 14222 52280 14418 52286
rect 10302 52246 10314 52280
rect 10486 52246 10498 52280
rect 10302 52240 10498 52246
rect 11568 52274 11764 52280
rect 11568 52240 11580 52274
rect 11752 52240 11764 52274
rect 4982 52234 5178 52240
rect 11568 52234 11764 52240
rect 12262 52274 12458 52280
rect 12262 52240 12274 52274
rect 12446 52240 12458 52274
rect 12262 52234 12458 52240
rect 12956 52274 13152 52280
rect 12956 52240 12968 52274
rect 13140 52240 13152 52274
rect 14222 52246 14234 52280
rect 14406 52246 14418 52280
rect 14222 52240 14418 52246
rect 14916 52280 15112 52286
rect 14916 52246 14928 52280
rect 15100 52246 15112 52280
rect 14916 52240 15112 52246
rect 15610 52280 15806 52286
rect 15610 52246 15622 52280
rect 15794 52246 15806 52280
rect 15610 52240 15806 52246
rect 16848 52284 17044 52290
rect 16848 52250 16860 52284
rect 17032 52250 17044 52284
rect 16848 52244 17044 52250
rect 17542 52284 17738 52290
rect 17542 52250 17554 52284
rect 17726 52250 17738 52284
rect 17542 52244 17738 52250
rect 18236 52284 18432 52290
rect 19532 52288 19728 52294
rect 20226 52328 20422 52334
rect 20226 52294 20238 52328
rect 20410 52294 20422 52328
rect 20226 52288 20422 52294
rect 18236 52250 18248 52284
rect 18420 52250 18432 52284
rect 18236 52244 18432 52250
rect 12956 52234 13152 52240
rect 19532 51670 19728 51676
rect 19532 51636 19544 51670
rect 19716 51636 19728 51670
rect 926 51620 1122 51626
rect 926 51586 938 51620
rect 1110 51586 1122 51620
rect 926 51580 1122 51586
rect 1620 51620 1816 51626
rect 1620 51586 1632 51620
rect 1804 51586 1816 51620
rect 1620 51580 1816 51586
rect 2314 51620 2510 51626
rect 6268 51622 6464 51628
rect 2314 51586 2326 51620
rect 2498 51586 2510 51620
rect 2314 51580 2510 51586
rect 3594 51616 3790 51622
rect 3594 51582 3606 51616
rect 3778 51582 3790 51616
rect 3594 51576 3790 51582
rect 4288 51616 4484 51622
rect 4288 51582 4300 51616
rect 4472 51582 4484 51616
rect 4288 51576 4484 51582
rect 4982 51616 5178 51622
rect 4982 51582 4994 51616
rect 5166 51582 5178 51616
rect 6268 51588 6280 51622
rect 6452 51588 6464 51622
rect 6268 51582 6464 51588
rect 6962 51622 7158 51628
rect 6962 51588 6974 51622
rect 7146 51588 7158 51622
rect 6962 51582 7158 51588
rect 7656 51622 7852 51628
rect 7656 51588 7668 51622
rect 7840 51588 7852 51622
rect 7656 51582 7852 51588
rect 8914 51622 9110 51628
rect 8914 51588 8926 51622
rect 9098 51588 9110 51622
rect 8914 51582 9110 51588
rect 9608 51622 9804 51628
rect 9608 51588 9620 51622
rect 9792 51588 9804 51622
rect 9608 51582 9804 51588
rect 10302 51622 10498 51628
rect 14222 51622 14418 51628
rect 10302 51588 10314 51622
rect 10486 51588 10498 51622
rect 10302 51582 10498 51588
rect 11568 51616 11764 51622
rect 11568 51582 11580 51616
rect 11752 51582 11764 51616
rect 4982 51576 5178 51582
rect 11568 51576 11764 51582
rect 12262 51616 12458 51622
rect 12262 51582 12274 51616
rect 12446 51582 12458 51616
rect 12262 51576 12458 51582
rect 12956 51616 13152 51622
rect 12956 51582 12968 51616
rect 13140 51582 13152 51616
rect 14222 51588 14234 51622
rect 14406 51588 14418 51622
rect 14222 51582 14418 51588
rect 14916 51622 15112 51628
rect 14916 51588 14928 51622
rect 15100 51588 15112 51622
rect 14916 51582 15112 51588
rect 15610 51622 15806 51628
rect 15610 51588 15622 51622
rect 15794 51588 15806 51622
rect 15610 51582 15806 51588
rect 16848 51626 17044 51632
rect 16848 51592 16860 51626
rect 17032 51592 17044 51626
rect 16848 51586 17044 51592
rect 17542 51626 17738 51632
rect 17542 51592 17554 51626
rect 17726 51592 17738 51626
rect 17542 51586 17738 51592
rect 18236 51626 18432 51632
rect 19532 51630 19728 51636
rect 20226 51670 20422 51676
rect 20226 51636 20238 51670
rect 20410 51636 20422 51670
rect 20226 51630 20422 51636
rect 18236 51592 18248 51626
rect 18420 51592 18432 51626
rect 18236 51586 18432 51592
rect 12956 51576 13152 51582
rect 19532 51012 19728 51018
rect 19532 50978 19544 51012
rect 19716 50978 19728 51012
rect 926 50962 1122 50968
rect 926 50928 938 50962
rect 1110 50928 1122 50962
rect 926 50922 1122 50928
rect 1620 50962 1816 50968
rect 1620 50928 1632 50962
rect 1804 50928 1816 50962
rect 1620 50922 1816 50928
rect 2314 50962 2510 50968
rect 6268 50964 6464 50970
rect 2314 50928 2326 50962
rect 2498 50928 2510 50962
rect 2314 50922 2510 50928
rect 3594 50958 3790 50964
rect 3594 50924 3606 50958
rect 3778 50924 3790 50958
rect 3594 50918 3790 50924
rect 4288 50958 4484 50964
rect 4288 50924 4300 50958
rect 4472 50924 4484 50958
rect 4288 50918 4484 50924
rect 4982 50958 5178 50964
rect 4982 50924 4994 50958
rect 5166 50924 5178 50958
rect 6268 50930 6280 50964
rect 6452 50930 6464 50964
rect 6268 50924 6464 50930
rect 6962 50964 7158 50970
rect 6962 50930 6974 50964
rect 7146 50930 7158 50964
rect 6962 50924 7158 50930
rect 7656 50964 7852 50970
rect 7656 50930 7668 50964
rect 7840 50930 7852 50964
rect 7656 50924 7852 50930
rect 8914 50964 9110 50970
rect 8914 50930 8926 50964
rect 9098 50930 9110 50964
rect 8914 50924 9110 50930
rect 9608 50964 9804 50970
rect 9608 50930 9620 50964
rect 9792 50930 9804 50964
rect 9608 50924 9804 50930
rect 10302 50964 10498 50970
rect 14222 50964 14418 50970
rect 10302 50930 10314 50964
rect 10486 50930 10498 50964
rect 10302 50924 10498 50930
rect 11568 50958 11764 50964
rect 11568 50924 11580 50958
rect 11752 50924 11764 50958
rect 4982 50918 5178 50924
rect 11568 50918 11764 50924
rect 12262 50958 12458 50964
rect 12262 50924 12274 50958
rect 12446 50924 12458 50958
rect 12262 50918 12458 50924
rect 12956 50958 13152 50964
rect 12956 50924 12968 50958
rect 13140 50924 13152 50958
rect 14222 50930 14234 50964
rect 14406 50930 14418 50964
rect 14222 50924 14418 50930
rect 14916 50964 15112 50970
rect 14916 50930 14928 50964
rect 15100 50930 15112 50964
rect 14916 50924 15112 50930
rect 15610 50964 15806 50970
rect 15610 50930 15622 50964
rect 15794 50930 15806 50964
rect 15610 50924 15806 50930
rect 16848 50968 17044 50974
rect 16848 50934 16860 50968
rect 17032 50934 17044 50968
rect 16848 50928 17044 50934
rect 17542 50968 17738 50974
rect 17542 50934 17554 50968
rect 17726 50934 17738 50968
rect 17542 50928 17738 50934
rect 18236 50968 18432 50974
rect 19532 50972 19728 50978
rect 20226 51012 20422 51018
rect 20226 50978 20238 51012
rect 20410 50978 20422 51012
rect 20226 50972 20422 50978
rect 18236 50934 18248 50968
rect 18420 50934 18432 50968
rect 18236 50928 18432 50934
rect 12956 50918 13152 50924
rect 19532 50354 19728 50360
rect 19532 50320 19544 50354
rect 19716 50320 19728 50354
rect 926 50304 1122 50310
rect 926 50270 938 50304
rect 1110 50270 1122 50304
rect 926 50264 1122 50270
rect 1620 50304 1816 50310
rect 1620 50270 1632 50304
rect 1804 50270 1816 50304
rect 1620 50264 1816 50270
rect 2314 50304 2510 50310
rect 6268 50306 6464 50312
rect 2314 50270 2326 50304
rect 2498 50270 2510 50304
rect 2314 50264 2510 50270
rect 3594 50300 3790 50306
rect 3594 50266 3606 50300
rect 3778 50266 3790 50300
rect 3594 50260 3790 50266
rect 4288 50300 4484 50306
rect 4288 50266 4300 50300
rect 4472 50266 4484 50300
rect 4288 50260 4484 50266
rect 4982 50300 5178 50306
rect 4982 50266 4994 50300
rect 5166 50266 5178 50300
rect 6268 50272 6280 50306
rect 6452 50272 6464 50306
rect 6268 50266 6464 50272
rect 6962 50306 7158 50312
rect 6962 50272 6974 50306
rect 7146 50272 7158 50306
rect 6962 50266 7158 50272
rect 7656 50306 7852 50312
rect 7656 50272 7668 50306
rect 7840 50272 7852 50306
rect 7656 50266 7852 50272
rect 8914 50306 9110 50312
rect 8914 50272 8926 50306
rect 9098 50272 9110 50306
rect 8914 50266 9110 50272
rect 9608 50306 9804 50312
rect 9608 50272 9620 50306
rect 9792 50272 9804 50306
rect 9608 50266 9804 50272
rect 10302 50306 10498 50312
rect 14222 50306 14418 50312
rect 10302 50272 10314 50306
rect 10486 50272 10498 50306
rect 10302 50266 10498 50272
rect 11568 50300 11764 50306
rect 11568 50266 11580 50300
rect 11752 50266 11764 50300
rect 4982 50260 5178 50266
rect 11568 50260 11764 50266
rect 12262 50300 12458 50306
rect 12262 50266 12274 50300
rect 12446 50266 12458 50300
rect 12262 50260 12458 50266
rect 12956 50300 13152 50306
rect 12956 50266 12968 50300
rect 13140 50266 13152 50300
rect 14222 50272 14234 50306
rect 14406 50272 14418 50306
rect 14222 50266 14418 50272
rect 14916 50306 15112 50312
rect 14916 50272 14928 50306
rect 15100 50272 15112 50306
rect 14916 50266 15112 50272
rect 15610 50306 15806 50312
rect 15610 50272 15622 50306
rect 15794 50272 15806 50306
rect 15610 50266 15806 50272
rect 16848 50310 17044 50316
rect 16848 50276 16860 50310
rect 17032 50276 17044 50310
rect 16848 50270 17044 50276
rect 17542 50310 17738 50316
rect 17542 50276 17554 50310
rect 17726 50276 17738 50310
rect 17542 50270 17738 50276
rect 18236 50310 18432 50316
rect 19532 50314 19728 50320
rect 20226 50354 20422 50360
rect 20226 50320 20238 50354
rect 20410 50320 20422 50354
rect 20226 50314 20422 50320
rect 18236 50276 18248 50310
rect 18420 50276 18432 50310
rect 18236 50270 18432 50276
rect 12956 50260 13152 50266
rect 19532 49696 19728 49702
rect 19532 49662 19544 49696
rect 19716 49662 19728 49696
rect 926 49646 1122 49652
rect 926 49612 938 49646
rect 1110 49612 1122 49646
rect 926 49606 1122 49612
rect 1620 49646 1816 49652
rect 1620 49612 1632 49646
rect 1804 49612 1816 49646
rect 1620 49606 1816 49612
rect 2314 49646 2510 49652
rect 6268 49648 6464 49654
rect 2314 49612 2326 49646
rect 2498 49612 2510 49646
rect 2314 49606 2510 49612
rect 3594 49642 3790 49648
rect 3594 49608 3606 49642
rect 3778 49608 3790 49642
rect 3594 49602 3790 49608
rect 4288 49642 4484 49648
rect 4288 49608 4300 49642
rect 4472 49608 4484 49642
rect 4288 49602 4484 49608
rect 4982 49642 5178 49648
rect 4982 49608 4994 49642
rect 5166 49608 5178 49642
rect 6268 49614 6280 49648
rect 6452 49614 6464 49648
rect 6268 49608 6464 49614
rect 6962 49648 7158 49654
rect 6962 49614 6974 49648
rect 7146 49614 7158 49648
rect 6962 49608 7158 49614
rect 7656 49648 7852 49654
rect 7656 49614 7668 49648
rect 7840 49614 7852 49648
rect 7656 49608 7852 49614
rect 8914 49648 9110 49654
rect 8914 49614 8926 49648
rect 9098 49614 9110 49648
rect 8914 49608 9110 49614
rect 9608 49648 9804 49654
rect 9608 49614 9620 49648
rect 9792 49614 9804 49648
rect 9608 49608 9804 49614
rect 10302 49648 10498 49654
rect 14222 49648 14418 49654
rect 10302 49614 10314 49648
rect 10486 49614 10498 49648
rect 10302 49608 10498 49614
rect 11568 49642 11764 49648
rect 11568 49608 11580 49642
rect 11752 49608 11764 49642
rect 4982 49602 5178 49608
rect 11568 49602 11764 49608
rect 12262 49642 12458 49648
rect 12262 49608 12274 49642
rect 12446 49608 12458 49642
rect 12262 49602 12458 49608
rect 12956 49642 13152 49648
rect 12956 49608 12968 49642
rect 13140 49608 13152 49642
rect 14222 49614 14234 49648
rect 14406 49614 14418 49648
rect 14222 49608 14418 49614
rect 14916 49648 15112 49654
rect 14916 49614 14928 49648
rect 15100 49614 15112 49648
rect 14916 49608 15112 49614
rect 15610 49648 15806 49654
rect 15610 49614 15622 49648
rect 15794 49614 15806 49648
rect 15610 49608 15806 49614
rect 16848 49652 17044 49658
rect 16848 49618 16860 49652
rect 17032 49618 17044 49652
rect 16848 49612 17044 49618
rect 17542 49652 17738 49658
rect 17542 49618 17554 49652
rect 17726 49618 17738 49652
rect 17542 49612 17738 49618
rect 18236 49652 18432 49658
rect 19532 49656 19728 49662
rect 20226 49696 20422 49702
rect 20226 49662 20238 49696
rect 20410 49662 20422 49696
rect 20226 49656 20422 49662
rect 18236 49618 18248 49652
rect 18420 49618 18432 49652
rect 18236 49612 18432 49618
rect 12956 49602 13152 49608
rect 21354 49318 21608 54504
rect 23278 54452 23316 54504
rect 23374 54452 23414 54720
rect 42322 54652 42518 54658
rect 42322 54618 42334 54652
rect 42506 54618 42518 54652
rect 42322 54612 42518 54618
rect 43016 54652 43212 54658
rect 43016 54618 43028 54652
rect 43200 54618 43212 54652
rect 43016 54612 43212 54618
rect 43710 54652 43906 54658
rect 43710 54618 43722 54652
rect 43894 54618 43906 54652
rect 43710 54612 43906 54618
rect 44404 54652 44600 54658
rect 44404 54618 44416 54652
rect 44588 54618 44600 54652
rect 44404 54612 44600 54618
rect 45098 54652 45294 54658
rect 45098 54618 45110 54652
rect 45282 54618 45294 54652
rect 45098 54612 45294 54618
rect 46330 54650 46526 54656
rect 46330 54616 46342 54650
rect 46514 54616 46526 54650
rect 46330 54610 46526 54616
rect 47024 54650 47220 54656
rect 47024 54616 47036 54650
rect 47208 54616 47220 54650
rect 47024 54610 47220 54616
rect 47718 54650 47914 54656
rect 47718 54616 47730 54650
rect 47902 54616 47914 54650
rect 47718 54610 47914 54616
rect 48412 54650 48608 54656
rect 48412 54616 48424 54650
rect 48596 54616 48608 54650
rect 48412 54610 48608 54616
rect 49106 54650 49302 54656
rect 49106 54616 49118 54650
rect 49290 54616 49302 54650
rect 49106 54610 49302 54616
rect 50342 54650 50538 54656
rect 50342 54616 50354 54650
rect 50526 54616 50538 54650
rect 50342 54610 50538 54616
rect 51036 54650 51232 54656
rect 51036 54616 51048 54650
rect 51220 54616 51232 54650
rect 51036 54610 51232 54616
rect 51730 54650 51926 54656
rect 51730 54616 51742 54650
rect 51914 54616 51926 54650
rect 51730 54610 51926 54616
rect 52424 54650 52620 54656
rect 52424 54616 52436 54650
rect 52608 54616 52620 54650
rect 52424 54610 52620 54616
rect 53118 54650 53314 54656
rect 53118 54616 53130 54650
rect 53302 54616 53314 54650
rect 53118 54610 53314 54616
rect 54352 54650 54548 54656
rect 54352 54616 54364 54650
rect 54536 54616 54548 54650
rect 54352 54610 54548 54616
rect 55046 54650 55242 54656
rect 55046 54616 55058 54650
rect 55230 54616 55242 54650
rect 55046 54610 55242 54616
rect 55740 54650 55936 54656
rect 55740 54616 55752 54650
rect 55924 54616 55936 54650
rect 55740 54610 55936 54616
rect 56434 54650 56630 54656
rect 56434 54616 56446 54650
rect 56618 54616 56630 54650
rect 56434 54610 56630 54616
rect 57128 54650 57324 54656
rect 57128 54616 57140 54650
rect 57312 54616 57324 54650
rect 57128 54610 57324 54616
rect 23278 54366 23414 54452
rect 23628 54274 23824 54280
rect 23628 54240 23640 54274
rect 23812 54240 23824 54274
rect 23628 54234 23824 54240
rect 24322 54274 24518 54280
rect 24322 54240 24334 54274
rect 24506 54240 24518 54274
rect 24322 54234 24518 54240
rect 25016 54274 25212 54280
rect 25016 54240 25028 54274
rect 25200 54240 25212 54274
rect 25016 54234 25212 54240
rect 25710 54274 25906 54280
rect 25710 54240 25722 54274
rect 25894 54240 25906 54274
rect 25710 54234 25906 54240
rect 26404 54274 26600 54280
rect 26404 54240 26416 54274
rect 26588 54240 26600 54274
rect 26404 54234 26600 54240
rect 27098 54274 27294 54280
rect 27098 54240 27110 54274
rect 27282 54240 27294 54274
rect 27098 54234 27294 54240
rect 27792 54274 27988 54280
rect 27792 54240 27804 54274
rect 27976 54240 27988 54274
rect 27792 54234 27988 54240
rect 28486 54274 28682 54280
rect 28486 54240 28498 54274
rect 28670 54240 28682 54274
rect 28486 54234 28682 54240
rect 29180 54274 29376 54280
rect 29180 54240 29192 54274
rect 29364 54240 29376 54274
rect 29180 54234 29376 54240
rect 29874 54274 30070 54280
rect 29874 54240 29886 54274
rect 30058 54240 30070 54274
rect 29874 54234 30070 54240
rect 28692 54056 29582 54100
rect 24280 53954 25168 54018
rect 28692 54012 28830 54056
rect 29474 54012 29582 54056
rect 28692 53958 29582 54012
rect 42322 53994 42518 54000
rect 42322 53960 42334 53994
rect 42506 53960 42518 53994
rect 42322 53954 42518 53960
rect 43016 53994 43212 54000
rect 43016 53960 43028 53994
rect 43200 53960 43212 53994
rect 43016 53954 43212 53960
rect 43710 53994 43906 54000
rect 43710 53960 43722 53994
rect 43894 53960 43906 53994
rect 43710 53954 43906 53960
rect 44404 53994 44600 54000
rect 44404 53960 44416 53994
rect 44588 53960 44600 53994
rect 44404 53954 44600 53960
rect 45098 53994 45294 54000
rect 45098 53960 45110 53994
rect 45282 53960 45294 53994
rect 45098 53954 45294 53960
rect 46330 53992 46526 53998
rect 46330 53958 46342 53992
rect 46514 53958 46526 53992
rect 24280 53898 24414 53954
rect 25058 53898 25168 53954
rect 46330 53952 46526 53958
rect 47024 53992 47220 53998
rect 47024 53958 47036 53992
rect 47208 53958 47220 53992
rect 47024 53952 47220 53958
rect 47718 53992 47914 53998
rect 47718 53958 47730 53992
rect 47902 53958 47914 53992
rect 47718 53952 47914 53958
rect 48412 53992 48608 53998
rect 48412 53958 48424 53992
rect 48596 53958 48608 53992
rect 48412 53952 48608 53958
rect 49106 53992 49302 53998
rect 49106 53958 49118 53992
rect 49290 53958 49302 53992
rect 49106 53952 49302 53958
rect 50342 53992 50538 53998
rect 50342 53958 50354 53992
rect 50526 53958 50538 53992
rect 50342 53952 50538 53958
rect 51036 53992 51232 53998
rect 51036 53958 51048 53992
rect 51220 53958 51232 53992
rect 51036 53952 51232 53958
rect 51730 53992 51926 53998
rect 51730 53958 51742 53992
rect 51914 53958 51926 53992
rect 51730 53952 51926 53958
rect 52424 53992 52620 53998
rect 52424 53958 52436 53992
rect 52608 53958 52620 53992
rect 52424 53952 52620 53958
rect 53118 53992 53314 53998
rect 53118 53958 53130 53992
rect 53302 53958 53314 53992
rect 53118 53952 53314 53958
rect 54352 53992 54548 53998
rect 54352 53958 54364 53992
rect 54536 53958 54548 53992
rect 54352 53952 54548 53958
rect 55046 53992 55242 53998
rect 55046 53958 55058 53992
rect 55230 53958 55242 53992
rect 55046 53952 55242 53958
rect 55740 53992 55936 53998
rect 55740 53958 55752 53992
rect 55924 53958 55936 53992
rect 55740 53952 55936 53958
rect 56434 53992 56630 53998
rect 56434 53958 56446 53992
rect 56618 53958 56630 53992
rect 56434 53952 56630 53958
rect 57128 53992 57324 53998
rect 57128 53958 57140 53992
rect 57312 53958 57324 53992
rect 57128 53952 57324 53958
rect 24280 53842 25168 53898
rect 23644 53648 23840 53654
rect 23644 53614 23656 53648
rect 23828 53614 23840 53648
rect 23644 53608 23840 53614
rect 24338 53648 24534 53654
rect 24338 53614 24350 53648
rect 24522 53614 24534 53648
rect 24338 53608 24534 53614
rect 25032 53648 25228 53654
rect 25032 53614 25044 53648
rect 25216 53614 25228 53648
rect 25032 53608 25228 53614
rect 25726 53648 25922 53654
rect 25726 53614 25738 53648
rect 25910 53614 25922 53648
rect 25726 53608 25922 53614
rect 26420 53648 26616 53654
rect 26420 53614 26432 53648
rect 26604 53614 26616 53648
rect 26420 53608 26616 53614
rect 27114 53648 27310 53654
rect 27114 53614 27126 53648
rect 27298 53614 27310 53648
rect 27114 53608 27310 53614
rect 27808 53648 28004 53654
rect 27808 53614 27820 53648
rect 27992 53614 28004 53648
rect 27808 53608 28004 53614
rect 28502 53648 28698 53654
rect 28502 53614 28514 53648
rect 28686 53614 28698 53648
rect 28502 53608 28698 53614
rect 29196 53648 29392 53654
rect 29196 53614 29208 53648
rect 29380 53614 29392 53648
rect 29196 53608 29392 53614
rect 29890 53648 30086 53654
rect 29890 53614 29902 53648
rect 30074 53614 30086 53648
rect 29890 53608 30086 53614
rect 42322 53336 42518 53342
rect 42322 53302 42334 53336
rect 42506 53302 42518 53336
rect 42322 53296 42518 53302
rect 43016 53336 43212 53342
rect 43016 53302 43028 53336
rect 43200 53302 43212 53336
rect 43016 53296 43212 53302
rect 43710 53336 43906 53342
rect 43710 53302 43722 53336
rect 43894 53302 43906 53336
rect 43710 53296 43906 53302
rect 44404 53336 44600 53342
rect 44404 53302 44416 53336
rect 44588 53302 44600 53336
rect 44404 53296 44600 53302
rect 45098 53336 45294 53342
rect 45098 53302 45110 53336
rect 45282 53302 45294 53336
rect 45098 53296 45294 53302
rect 46330 53334 46526 53340
rect 46330 53300 46342 53334
rect 46514 53300 46526 53334
rect 46330 53294 46526 53300
rect 47024 53334 47220 53340
rect 47024 53300 47036 53334
rect 47208 53300 47220 53334
rect 47024 53294 47220 53300
rect 47718 53334 47914 53340
rect 47718 53300 47730 53334
rect 47902 53300 47914 53334
rect 47718 53294 47914 53300
rect 48412 53334 48608 53340
rect 48412 53300 48424 53334
rect 48596 53300 48608 53334
rect 48412 53294 48608 53300
rect 49106 53334 49302 53340
rect 49106 53300 49118 53334
rect 49290 53300 49302 53334
rect 49106 53294 49302 53300
rect 50342 53334 50538 53340
rect 50342 53300 50354 53334
rect 50526 53300 50538 53334
rect 50342 53294 50538 53300
rect 51036 53334 51232 53340
rect 51036 53300 51048 53334
rect 51220 53300 51232 53334
rect 51036 53294 51232 53300
rect 51730 53334 51926 53340
rect 51730 53300 51742 53334
rect 51914 53300 51926 53334
rect 51730 53294 51926 53300
rect 52424 53334 52620 53340
rect 52424 53300 52436 53334
rect 52608 53300 52620 53334
rect 52424 53294 52620 53300
rect 53118 53334 53314 53340
rect 53118 53300 53130 53334
rect 53302 53300 53314 53334
rect 53118 53294 53314 53300
rect 54352 53334 54548 53340
rect 54352 53300 54364 53334
rect 54536 53300 54548 53334
rect 54352 53294 54548 53300
rect 55046 53334 55242 53340
rect 55046 53300 55058 53334
rect 55230 53300 55242 53334
rect 55046 53294 55242 53300
rect 55740 53334 55936 53340
rect 55740 53300 55752 53334
rect 55924 53300 55936 53334
rect 55740 53294 55936 53300
rect 56434 53334 56630 53340
rect 56434 53300 56446 53334
rect 56618 53300 56630 53334
rect 56434 53294 56630 53300
rect 57128 53334 57324 53340
rect 57128 53300 57140 53334
rect 57312 53300 57324 53334
rect 57128 53294 57324 53300
rect 30360 53048 30510 53106
rect 23644 52990 23840 52996
rect 23644 52956 23656 52990
rect 23828 52956 23840 52990
rect 23644 52950 23840 52956
rect 24338 52990 24534 52996
rect 24338 52956 24350 52990
rect 24522 52956 24534 52990
rect 24338 52950 24534 52956
rect 25032 52990 25228 52996
rect 25032 52956 25044 52990
rect 25216 52956 25228 52990
rect 25032 52950 25228 52956
rect 25726 52990 25922 52996
rect 25726 52956 25738 52990
rect 25910 52956 25922 52990
rect 25726 52950 25922 52956
rect 26420 52990 26616 52996
rect 26420 52956 26432 52990
rect 26604 52956 26616 52990
rect 26420 52950 26616 52956
rect 27114 52990 27310 52996
rect 27114 52956 27126 52990
rect 27298 52956 27310 52990
rect 27114 52950 27310 52956
rect 27808 52990 28004 52996
rect 27808 52956 27820 52990
rect 27992 52956 28004 52990
rect 27808 52950 28004 52956
rect 28502 52990 28698 52996
rect 28502 52956 28514 52990
rect 28686 52956 28698 52990
rect 28502 52950 28698 52956
rect 29196 52990 29392 52996
rect 29196 52956 29208 52990
rect 29380 52956 29392 52990
rect 29196 52950 29392 52956
rect 29890 52990 30086 52996
rect 29890 52956 29902 52990
rect 30074 52956 30086 52990
rect 29890 52950 30086 52956
rect 30360 52964 30390 53048
rect 30444 52964 30510 53048
rect 30360 52892 30510 52964
rect 42322 52678 42518 52684
rect 42322 52644 42334 52678
rect 42506 52644 42518 52678
rect 42322 52638 42518 52644
rect 43016 52678 43212 52684
rect 43016 52644 43028 52678
rect 43200 52644 43212 52678
rect 43016 52638 43212 52644
rect 43710 52678 43906 52684
rect 43710 52644 43722 52678
rect 43894 52644 43906 52678
rect 43710 52638 43906 52644
rect 44404 52678 44600 52684
rect 44404 52644 44416 52678
rect 44588 52644 44600 52678
rect 44404 52638 44600 52644
rect 45098 52678 45294 52684
rect 45098 52644 45110 52678
rect 45282 52644 45294 52678
rect 45098 52638 45294 52644
rect 46330 52676 46526 52682
rect 46330 52642 46342 52676
rect 46514 52642 46526 52676
rect 46330 52636 46526 52642
rect 47024 52676 47220 52682
rect 47024 52642 47036 52676
rect 47208 52642 47220 52676
rect 47024 52636 47220 52642
rect 47718 52676 47914 52682
rect 47718 52642 47730 52676
rect 47902 52642 47914 52676
rect 47718 52636 47914 52642
rect 48412 52676 48608 52682
rect 48412 52642 48424 52676
rect 48596 52642 48608 52676
rect 48412 52636 48608 52642
rect 49106 52676 49302 52682
rect 49106 52642 49118 52676
rect 49290 52642 49302 52676
rect 49106 52636 49302 52642
rect 50342 52676 50538 52682
rect 50342 52642 50354 52676
rect 50526 52642 50538 52676
rect 50342 52636 50538 52642
rect 51036 52676 51232 52682
rect 51036 52642 51048 52676
rect 51220 52642 51232 52676
rect 51036 52636 51232 52642
rect 51730 52676 51926 52682
rect 51730 52642 51742 52676
rect 51914 52642 51926 52676
rect 51730 52636 51926 52642
rect 52424 52676 52620 52682
rect 52424 52642 52436 52676
rect 52608 52642 52620 52676
rect 52424 52636 52620 52642
rect 53118 52676 53314 52682
rect 53118 52642 53130 52676
rect 53302 52642 53314 52676
rect 53118 52636 53314 52642
rect 54352 52676 54548 52682
rect 54352 52642 54364 52676
rect 54536 52642 54548 52676
rect 54352 52636 54548 52642
rect 55046 52676 55242 52682
rect 55046 52642 55058 52676
rect 55230 52642 55242 52676
rect 55046 52636 55242 52642
rect 55740 52676 55936 52682
rect 55740 52642 55752 52676
rect 55924 52642 55936 52676
rect 55740 52636 55936 52642
rect 56434 52676 56630 52682
rect 56434 52642 56446 52676
rect 56618 52642 56630 52676
rect 56434 52636 56630 52642
rect 57128 52676 57324 52682
rect 57128 52642 57140 52676
rect 57312 52642 57324 52676
rect 57128 52636 57324 52642
rect 23644 52332 23840 52338
rect 23644 52298 23656 52332
rect 23828 52298 23840 52332
rect 23644 52292 23840 52298
rect 24338 52332 24534 52338
rect 24338 52298 24350 52332
rect 24522 52298 24534 52332
rect 24338 52292 24534 52298
rect 25032 52332 25228 52338
rect 25032 52298 25044 52332
rect 25216 52298 25228 52332
rect 25032 52292 25228 52298
rect 25726 52332 25922 52338
rect 25726 52298 25738 52332
rect 25910 52298 25922 52332
rect 25726 52292 25922 52298
rect 26420 52332 26616 52338
rect 26420 52298 26432 52332
rect 26604 52298 26616 52332
rect 26420 52292 26616 52298
rect 27114 52332 27310 52338
rect 27114 52298 27126 52332
rect 27298 52298 27310 52332
rect 27114 52292 27310 52298
rect 27808 52332 28004 52338
rect 27808 52298 27820 52332
rect 27992 52298 28004 52332
rect 27808 52292 28004 52298
rect 28502 52332 28698 52338
rect 28502 52298 28514 52332
rect 28686 52298 28698 52332
rect 28502 52292 28698 52298
rect 29196 52332 29392 52338
rect 29196 52298 29208 52332
rect 29380 52298 29392 52332
rect 29196 52292 29392 52298
rect 29890 52332 30086 52338
rect 29890 52298 29902 52332
rect 30074 52298 30086 52332
rect 57610 52328 57800 52450
rect 29890 52292 30086 52298
rect 42670 52222 45316 52310
rect 28708 52114 29598 52158
rect 24296 52012 25184 52076
rect 28708 52070 28846 52114
rect 29490 52070 29598 52114
rect 28708 52016 29598 52070
rect 42670 52020 42968 52222
rect 45142 52020 45316 52222
rect 24296 51956 24430 52012
rect 25074 51956 25184 52012
rect 24296 51900 25184 51956
rect 42670 51908 45316 52020
rect 46664 52222 49310 52310
rect 46664 52020 46962 52222
rect 49136 52020 49310 52222
rect 46664 51908 49310 52020
rect 50686 52222 53332 52310
rect 50686 52020 50984 52222
rect 53158 52020 53332 52222
rect 50686 51908 53332 52020
rect 54708 52222 57354 52310
rect 54708 52020 55006 52222
rect 57180 52020 57354 52222
rect 54708 51908 57354 52020
rect 57610 52026 57636 52328
rect 57760 52026 57800 52328
rect 57610 51908 57800 52026
rect 42314 51770 42510 51776
rect 42314 51736 42326 51770
rect 42498 51736 42510 51770
rect 42314 51730 42510 51736
rect 43008 51770 43204 51776
rect 43008 51736 43020 51770
rect 43192 51736 43204 51770
rect 43008 51730 43204 51736
rect 43702 51770 43898 51776
rect 43702 51736 43714 51770
rect 43886 51736 43898 51770
rect 43702 51730 43898 51736
rect 44396 51770 44592 51776
rect 44396 51736 44408 51770
rect 44580 51736 44592 51770
rect 44396 51730 44592 51736
rect 45090 51770 45286 51776
rect 45090 51736 45102 51770
rect 45274 51736 45286 51770
rect 45090 51730 45286 51736
rect 46308 51770 46504 51776
rect 46308 51736 46320 51770
rect 46492 51736 46504 51770
rect 46308 51730 46504 51736
rect 47002 51770 47198 51776
rect 47002 51736 47014 51770
rect 47186 51736 47198 51770
rect 47002 51730 47198 51736
rect 47696 51770 47892 51776
rect 47696 51736 47708 51770
rect 47880 51736 47892 51770
rect 47696 51730 47892 51736
rect 48390 51770 48586 51776
rect 48390 51736 48402 51770
rect 48574 51736 48586 51770
rect 48390 51730 48586 51736
rect 49084 51770 49280 51776
rect 49084 51736 49096 51770
rect 49268 51736 49280 51770
rect 49084 51730 49280 51736
rect 50330 51770 50526 51776
rect 50330 51736 50342 51770
rect 50514 51736 50526 51770
rect 50330 51730 50526 51736
rect 51024 51770 51220 51776
rect 51024 51736 51036 51770
rect 51208 51736 51220 51770
rect 51024 51730 51220 51736
rect 51718 51770 51914 51776
rect 51718 51736 51730 51770
rect 51902 51736 51914 51770
rect 51718 51730 51914 51736
rect 52412 51770 52608 51776
rect 52412 51736 52424 51770
rect 52596 51736 52608 51770
rect 52412 51730 52608 51736
rect 53106 51770 53302 51776
rect 53106 51736 53118 51770
rect 53290 51736 53302 51770
rect 53106 51730 53302 51736
rect 54352 51770 54548 51776
rect 54352 51736 54364 51770
rect 54536 51736 54548 51770
rect 54352 51730 54548 51736
rect 55046 51770 55242 51776
rect 55046 51736 55058 51770
rect 55230 51736 55242 51770
rect 55046 51730 55242 51736
rect 55740 51770 55936 51776
rect 55740 51736 55752 51770
rect 55924 51736 55936 51770
rect 55740 51730 55936 51736
rect 56434 51770 56630 51776
rect 56434 51736 56446 51770
rect 56618 51736 56630 51770
rect 56434 51730 56630 51736
rect 57128 51770 57324 51776
rect 57128 51736 57140 51770
rect 57312 51736 57324 51770
rect 57128 51730 57324 51736
rect 42314 51112 42510 51118
rect 42314 51078 42326 51112
rect 42498 51078 42510 51112
rect 42314 51072 42510 51078
rect 43008 51112 43204 51118
rect 43008 51078 43020 51112
rect 43192 51078 43204 51112
rect 43008 51072 43204 51078
rect 43702 51112 43898 51118
rect 43702 51078 43714 51112
rect 43886 51078 43898 51112
rect 43702 51072 43898 51078
rect 44396 51112 44592 51118
rect 44396 51078 44408 51112
rect 44580 51078 44592 51112
rect 44396 51072 44592 51078
rect 45090 51112 45286 51118
rect 45090 51078 45102 51112
rect 45274 51078 45286 51112
rect 45090 51072 45286 51078
rect 46308 51112 46504 51118
rect 46308 51078 46320 51112
rect 46492 51078 46504 51112
rect 46308 51072 46504 51078
rect 47002 51112 47198 51118
rect 47002 51078 47014 51112
rect 47186 51078 47198 51112
rect 47002 51072 47198 51078
rect 47696 51112 47892 51118
rect 47696 51078 47708 51112
rect 47880 51078 47892 51112
rect 47696 51072 47892 51078
rect 48390 51112 48586 51118
rect 48390 51078 48402 51112
rect 48574 51078 48586 51112
rect 48390 51072 48586 51078
rect 49084 51112 49280 51118
rect 49084 51078 49096 51112
rect 49268 51078 49280 51112
rect 49084 51072 49280 51078
rect 50330 51112 50526 51118
rect 50330 51078 50342 51112
rect 50514 51078 50526 51112
rect 50330 51072 50526 51078
rect 51024 51112 51220 51118
rect 51024 51078 51036 51112
rect 51208 51078 51220 51112
rect 51024 51072 51220 51078
rect 51718 51112 51914 51118
rect 51718 51078 51730 51112
rect 51902 51078 51914 51112
rect 51718 51072 51914 51078
rect 52412 51112 52608 51118
rect 52412 51078 52424 51112
rect 52596 51078 52608 51112
rect 52412 51072 52608 51078
rect 53106 51112 53302 51118
rect 53106 51078 53118 51112
rect 53290 51078 53302 51112
rect 53106 51072 53302 51078
rect 54352 51112 54548 51118
rect 54352 51078 54364 51112
rect 54536 51078 54548 51112
rect 54352 51072 54548 51078
rect 55046 51112 55242 51118
rect 55046 51078 55058 51112
rect 55230 51078 55242 51112
rect 55046 51072 55242 51078
rect 55740 51112 55936 51118
rect 55740 51078 55752 51112
rect 55924 51078 55936 51112
rect 55740 51072 55936 51078
rect 56434 51112 56630 51118
rect 56434 51078 56446 51112
rect 56618 51078 56630 51112
rect 56434 51072 56630 51078
rect 57128 51112 57324 51118
rect 57128 51078 57140 51112
rect 57312 51078 57324 51112
rect 57128 51072 57324 51078
rect 42314 50454 42510 50460
rect 42314 50420 42326 50454
rect 42498 50420 42510 50454
rect 42314 50414 42510 50420
rect 43008 50454 43204 50460
rect 43008 50420 43020 50454
rect 43192 50420 43204 50454
rect 43008 50414 43204 50420
rect 43702 50454 43898 50460
rect 43702 50420 43714 50454
rect 43886 50420 43898 50454
rect 43702 50414 43898 50420
rect 44396 50454 44592 50460
rect 44396 50420 44408 50454
rect 44580 50420 44592 50454
rect 44396 50414 44592 50420
rect 45090 50454 45286 50460
rect 45090 50420 45102 50454
rect 45274 50420 45286 50454
rect 45090 50414 45286 50420
rect 46308 50454 46504 50460
rect 46308 50420 46320 50454
rect 46492 50420 46504 50454
rect 46308 50414 46504 50420
rect 47002 50454 47198 50460
rect 47002 50420 47014 50454
rect 47186 50420 47198 50454
rect 47002 50414 47198 50420
rect 47696 50454 47892 50460
rect 47696 50420 47708 50454
rect 47880 50420 47892 50454
rect 47696 50414 47892 50420
rect 48390 50454 48586 50460
rect 48390 50420 48402 50454
rect 48574 50420 48586 50454
rect 48390 50414 48586 50420
rect 49084 50454 49280 50460
rect 49084 50420 49096 50454
rect 49268 50420 49280 50454
rect 49084 50414 49280 50420
rect 50330 50454 50526 50460
rect 50330 50420 50342 50454
rect 50514 50420 50526 50454
rect 50330 50414 50526 50420
rect 51024 50454 51220 50460
rect 51024 50420 51036 50454
rect 51208 50420 51220 50454
rect 51024 50414 51220 50420
rect 51718 50454 51914 50460
rect 51718 50420 51730 50454
rect 51902 50420 51914 50454
rect 51718 50414 51914 50420
rect 52412 50454 52608 50460
rect 52412 50420 52424 50454
rect 52596 50420 52608 50454
rect 52412 50414 52608 50420
rect 53106 50454 53302 50460
rect 53106 50420 53118 50454
rect 53290 50420 53302 50454
rect 53106 50414 53302 50420
rect 54352 50454 54548 50460
rect 54352 50420 54364 50454
rect 54536 50420 54548 50454
rect 54352 50414 54548 50420
rect 55046 50454 55242 50460
rect 55046 50420 55058 50454
rect 55230 50420 55242 50454
rect 55046 50414 55242 50420
rect 55740 50454 55936 50460
rect 55740 50420 55752 50454
rect 55924 50420 55936 50454
rect 55740 50414 55936 50420
rect 56434 50454 56630 50460
rect 56434 50420 56446 50454
rect 56618 50420 56630 50454
rect 56434 50414 56630 50420
rect 57128 50454 57324 50460
rect 57128 50420 57140 50454
rect 57312 50420 57324 50454
rect 59906 50432 60318 60764
rect 71008 59102 71062 61670
rect 71146 59102 71224 61670
rect 71300 61644 71306 61816
rect 71340 61644 71346 61816
rect 71300 61632 71346 61644
rect 71958 61816 72004 61828
rect 71958 61644 71964 61816
rect 71998 61644 72004 61816
rect 71958 61632 72004 61644
rect 72616 61816 72662 61828
rect 72616 61644 72622 61816
rect 72656 61644 72662 61816
rect 73260 61816 73336 62632
rect 73932 62632 73938 62804
rect 73972 62632 73978 62804
rect 74872 62700 75088 62846
rect 78722 62860 78776 65428
rect 78860 62860 78938 65428
rect 79014 65402 79020 65574
rect 79054 65402 79060 65574
rect 79014 65390 79060 65402
rect 79672 65574 79718 65586
rect 79672 65402 79678 65574
rect 79712 65402 79718 65574
rect 79672 65390 79718 65402
rect 80330 65574 80376 65586
rect 80330 65402 80336 65574
rect 80370 65402 80376 65574
rect 80952 65574 81076 66396
rect 81646 66396 81652 66568
rect 81686 66396 81692 66568
rect 81646 66384 81692 66396
rect 80952 65472 80994 65574
rect 80330 65390 80376 65402
rect 80988 65402 80994 65472
rect 81028 65472 81076 65574
rect 81646 65574 81692 65586
rect 81028 65402 81034 65472
rect 80988 65390 81034 65402
rect 81646 65402 81652 65574
rect 81686 65402 81692 65574
rect 81646 65390 81692 65402
rect 79014 64880 79060 64892
rect 79014 64708 79020 64880
rect 79054 64708 79060 64880
rect 79014 64696 79060 64708
rect 79672 64880 79718 64892
rect 79672 64708 79678 64880
rect 79712 64708 79718 64880
rect 79672 64696 79718 64708
rect 80330 64880 80376 64892
rect 80330 64708 80336 64880
rect 80370 64708 80376 64880
rect 80330 64696 80376 64708
rect 80988 64880 81034 64892
rect 80988 64708 80994 64880
rect 81028 64708 81034 64880
rect 80988 64696 81034 64708
rect 81646 64880 81692 64892
rect 81646 64708 81652 64880
rect 81686 64708 81692 64880
rect 81646 64696 81692 64708
rect 79014 64186 79060 64198
rect 79014 64014 79020 64186
rect 79054 64014 79060 64186
rect 79014 64002 79060 64014
rect 79672 64186 79718 64198
rect 79672 64014 79678 64186
rect 79712 64014 79718 64186
rect 79672 64002 79718 64014
rect 80330 64186 80376 64198
rect 80330 64014 80336 64186
rect 80370 64014 80376 64186
rect 80330 64002 80376 64014
rect 80988 64186 81034 64198
rect 80988 64014 80994 64186
rect 81028 64014 81034 64186
rect 80988 64002 81034 64014
rect 81646 64186 81692 64198
rect 81646 64014 81652 64186
rect 81686 64014 81692 64186
rect 81646 64002 81692 64014
rect 79014 63492 79060 63504
rect 79014 63320 79020 63492
rect 79054 63320 79060 63492
rect 79014 63308 79060 63320
rect 79672 63492 79718 63504
rect 79672 63320 79678 63492
rect 79712 63320 79718 63492
rect 79672 63308 79718 63320
rect 80330 63492 80376 63504
rect 80330 63320 80336 63492
rect 80370 63320 80376 63492
rect 80330 63308 80376 63320
rect 80988 63492 81034 63504
rect 80988 63320 80994 63492
rect 81028 63320 81034 63492
rect 80988 63308 81034 63320
rect 81646 63492 81692 63504
rect 81646 63320 81652 63492
rect 81686 63320 81692 63492
rect 81646 63308 81692 63320
rect 75164 62784 75210 62796
rect 73932 62620 73978 62632
rect 75164 62612 75170 62784
rect 75204 62612 75210 62784
rect 75164 62600 75210 62612
rect 75822 62784 75868 62796
rect 75822 62612 75828 62784
rect 75862 62612 75868 62784
rect 75822 62600 75868 62612
rect 76480 62784 76526 62796
rect 76480 62612 76486 62784
rect 76520 62612 76526 62784
rect 77138 62784 77184 62796
rect 77138 62756 77144 62784
rect 76480 62600 76526 62612
rect 77124 62612 77144 62756
rect 77178 62756 77184 62784
rect 77796 62784 77842 62796
rect 77178 62612 77200 62756
rect 73260 61708 73280 61816
rect 72616 61632 72662 61644
rect 73274 61644 73280 61708
rect 73314 61708 73336 61816
rect 73932 61816 73978 61828
rect 73314 61644 73320 61708
rect 73274 61632 73320 61644
rect 73932 61644 73938 61816
rect 73972 61644 73978 61816
rect 75164 61796 75210 61808
rect 73932 61632 73978 61644
rect 74872 61650 75088 61796
rect 71300 61122 71346 61134
rect 71300 60950 71306 61122
rect 71340 60950 71346 61122
rect 71300 60938 71346 60950
rect 71958 61122 72004 61134
rect 71958 60950 71964 61122
rect 71998 60950 72004 61122
rect 71958 60938 72004 60950
rect 72616 61122 72662 61134
rect 72616 60950 72622 61122
rect 72656 60950 72662 61122
rect 72616 60938 72662 60950
rect 73274 61122 73320 61134
rect 73274 60950 73280 61122
rect 73314 60950 73320 61122
rect 73274 60938 73320 60950
rect 73932 61122 73978 61134
rect 73932 60950 73938 61122
rect 73972 60950 73978 61122
rect 73932 60938 73978 60950
rect 71300 60428 71346 60440
rect 71300 60256 71306 60428
rect 71340 60256 71346 60428
rect 71300 60244 71346 60256
rect 71958 60428 72004 60440
rect 71958 60256 71964 60428
rect 71998 60256 72004 60428
rect 71958 60244 72004 60256
rect 72616 60428 72662 60440
rect 72616 60256 72622 60428
rect 72656 60256 72662 60428
rect 72616 60244 72662 60256
rect 73274 60428 73320 60440
rect 73274 60256 73280 60428
rect 73314 60256 73320 60428
rect 73274 60244 73320 60256
rect 73932 60428 73978 60440
rect 73932 60256 73938 60428
rect 73972 60256 73978 60428
rect 73932 60244 73978 60256
rect 71300 59734 71346 59746
rect 71300 59562 71306 59734
rect 71340 59562 71346 59734
rect 71300 59550 71346 59562
rect 71958 59734 72004 59746
rect 71958 59562 71964 59734
rect 71998 59562 72004 59734
rect 71958 59550 72004 59562
rect 72616 59734 72662 59746
rect 72616 59562 72622 59734
rect 72656 59562 72662 59734
rect 72616 59550 72662 59562
rect 73274 59734 73320 59746
rect 73274 59562 73280 59734
rect 73314 59562 73320 59734
rect 73274 59550 73320 59562
rect 73932 59734 73978 59746
rect 73932 59562 73938 59734
rect 73972 59562 73978 59734
rect 73932 59550 73978 59562
rect 71008 58956 71224 59102
rect 74872 59082 74926 61650
rect 75010 59082 75088 61650
rect 75164 61624 75170 61796
rect 75204 61624 75210 61796
rect 75164 61612 75210 61624
rect 75822 61796 75868 61808
rect 75822 61624 75828 61796
rect 75862 61624 75868 61796
rect 75822 61612 75868 61624
rect 76480 61796 76526 61808
rect 76480 61624 76486 61796
rect 76520 61624 76526 61796
rect 77124 61796 77200 62612
rect 77796 62612 77802 62784
rect 77836 62612 77842 62784
rect 78722 62714 78938 62860
rect 79014 62798 79060 62810
rect 79014 62626 79020 62798
rect 79054 62626 79060 62798
rect 79014 62614 79060 62626
rect 79672 62798 79718 62810
rect 79672 62626 79678 62798
rect 79712 62626 79718 62798
rect 79672 62614 79718 62626
rect 80330 62798 80376 62810
rect 80330 62626 80336 62798
rect 80370 62626 80376 62798
rect 80988 62798 81034 62810
rect 80988 62770 80994 62798
rect 80330 62614 80376 62626
rect 80974 62626 80994 62770
rect 81028 62770 81034 62798
rect 81646 62798 81692 62810
rect 81028 62626 81050 62770
rect 77796 62600 77842 62612
rect 79014 61810 79060 61822
rect 77124 61688 77144 61796
rect 76480 61612 76526 61624
rect 77138 61624 77144 61688
rect 77178 61688 77200 61796
rect 77796 61796 77842 61808
rect 77178 61624 77184 61688
rect 77138 61612 77184 61624
rect 77796 61624 77802 61796
rect 77836 61624 77842 61796
rect 77796 61612 77842 61624
rect 78722 61664 78938 61810
rect 75164 61102 75210 61114
rect 75164 60930 75170 61102
rect 75204 60930 75210 61102
rect 75164 60918 75210 60930
rect 75822 61102 75868 61114
rect 75822 60930 75828 61102
rect 75862 60930 75868 61102
rect 75822 60918 75868 60930
rect 76480 61102 76526 61114
rect 76480 60930 76486 61102
rect 76520 60930 76526 61102
rect 76480 60918 76526 60930
rect 77138 61102 77184 61114
rect 77138 60930 77144 61102
rect 77178 60930 77184 61102
rect 77138 60918 77184 60930
rect 77796 61102 77842 61114
rect 77796 60930 77802 61102
rect 77836 60930 77842 61102
rect 77796 60918 77842 60930
rect 75164 60408 75210 60420
rect 75164 60236 75170 60408
rect 75204 60236 75210 60408
rect 75164 60224 75210 60236
rect 75822 60408 75868 60420
rect 75822 60236 75828 60408
rect 75862 60236 75868 60408
rect 75822 60224 75868 60236
rect 76480 60408 76526 60420
rect 76480 60236 76486 60408
rect 76520 60236 76526 60408
rect 76480 60224 76526 60236
rect 77138 60408 77184 60420
rect 77138 60236 77144 60408
rect 77178 60236 77184 60408
rect 77138 60224 77184 60236
rect 77796 60408 77842 60420
rect 77796 60236 77802 60408
rect 77836 60236 77842 60408
rect 77796 60224 77842 60236
rect 75164 59714 75210 59726
rect 75164 59542 75170 59714
rect 75204 59542 75210 59714
rect 75164 59530 75210 59542
rect 75822 59714 75868 59726
rect 75822 59542 75828 59714
rect 75862 59542 75868 59714
rect 75822 59530 75868 59542
rect 76480 59714 76526 59726
rect 76480 59542 76486 59714
rect 76520 59542 76526 59714
rect 76480 59530 76526 59542
rect 77138 59714 77184 59726
rect 77138 59542 77144 59714
rect 77178 59542 77184 59714
rect 77138 59530 77184 59542
rect 77796 59714 77842 59726
rect 77796 59542 77802 59714
rect 77836 59542 77842 59714
rect 77796 59530 77842 59542
rect 71300 59040 71346 59052
rect 71300 58868 71306 59040
rect 71340 58868 71346 59040
rect 71300 58856 71346 58868
rect 71958 59040 72004 59052
rect 71958 58868 71964 59040
rect 71998 58868 72004 59040
rect 71958 58856 72004 58868
rect 72616 59040 72662 59052
rect 72616 58868 72622 59040
rect 72656 58868 72662 59040
rect 73274 59040 73320 59052
rect 73274 59006 73280 59040
rect 72616 58856 72662 58868
rect 73260 58868 73280 59006
rect 73314 59006 73320 59040
rect 73932 59040 73978 59052
rect 73314 58868 73336 59006
rect 71300 58040 71346 58052
rect 71008 57894 71224 58040
rect 71008 55326 71062 57894
rect 71146 55326 71224 57894
rect 71300 57868 71306 58040
rect 71340 57868 71346 58040
rect 71300 57856 71346 57868
rect 71958 58040 72004 58052
rect 71958 57868 71964 58040
rect 71998 57868 72004 58040
rect 71958 57856 72004 57868
rect 72616 58040 72662 58052
rect 72616 57868 72622 58040
rect 72656 57868 72662 58040
rect 73260 58040 73336 58868
rect 73932 58868 73938 59040
rect 73972 58868 73978 59040
rect 74872 58936 75088 59082
rect 78722 59096 78776 61664
rect 78860 59096 78938 61664
rect 79014 61638 79020 61810
rect 79054 61638 79060 61810
rect 79014 61626 79060 61638
rect 79672 61810 79718 61822
rect 79672 61638 79678 61810
rect 79712 61638 79718 61810
rect 79672 61626 79718 61638
rect 80330 61810 80376 61822
rect 80330 61638 80336 61810
rect 80370 61638 80376 61810
rect 80974 61810 81050 62626
rect 81646 62626 81652 62798
rect 81686 62626 81692 62798
rect 81646 62614 81692 62626
rect 80974 61702 80994 61810
rect 80330 61626 80376 61638
rect 80988 61638 80994 61702
rect 81028 61702 81050 61810
rect 81646 61810 81692 61822
rect 81028 61638 81034 61702
rect 80988 61626 81034 61638
rect 81646 61638 81652 61810
rect 81686 61638 81692 61810
rect 81646 61626 81692 61638
rect 79014 61116 79060 61128
rect 79014 60944 79020 61116
rect 79054 60944 79060 61116
rect 79014 60932 79060 60944
rect 79672 61116 79718 61128
rect 79672 60944 79678 61116
rect 79712 60944 79718 61116
rect 79672 60932 79718 60944
rect 80330 61116 80376 61128
rect 80330 60944 80336 61116
rect 80370 60944 80376 61116
rect 80330 60932 80376 60944
rect 80988 61116 81034 61128
rect 80988 60944 80994 61116
rect 81028 60944 81034 61116
rect 80988 60932 81034 60944
rect 81646 61116 81692 61128
rect 81646 60944 81652 61116
rect 81686 60944 81692 61116
rect 81646 60932 81692 60944
rect 79014 60422 79060 60434
rect 79014 60250 79020 60422
rect 79054 60250 79060 60422
rect 79014 60238 79060 60250
rect 79672 60422 79718 60434
rect 79672 60250 79678 60422
rect 79712 60250 79718 60422
rect 79672 60238 79718 60250
rect 80330 60422 80376 60434
rect 80330 60250 80336 60422
rect 80370 60250 80376 60422
rect 80330 60238 80376 60250
rect 80988 60422 81034 60434
rect 80988 60250 80994 60422
rect 81028 60250 81034 60422
rect 80988 60238 81034 60250
rect 81646 60422 81692 60434
rect 81646 60250 81652 60422
rect 81686 60250 81692 60422
rect 81646 60238 81692 60250
rect 79014 59728 79060 59740
rect 79014 59556 79020 59728
rect 79054 59556 79060 59728
rect 79014 59544 79060 59556
rect 79672 59728 79718 59740
rect 79672 59556 79678 59728
rect 79712 59556 79718 59728
rect 79672 59544 79718 59556
rect 80330 59728 80376 59740
rect 80330 59556 80336 59728
rect 80370 59556 80376 59728
rect 80330 59544 80376 59556
rect 80988 59728 81034 59740
rect 80988 59556 80994 59728
rect 81028 59556 81034 59728
rect 80988 59544 81034 59556
rect 81646 59728 81692 59740
rect 81646 59556 81652 59728
rect 81686 59556 81692 59728
rect 81646 59544 81692 59556
rect 75164 59020 75210 59032
rect 73932 58856 73978 58868
rect 75164 58848 75170 59020
rect 75204 58848 75210 59020
rect 75164 58836 75210 58848
rect 75822 59020 75868 59032
rect 75822 58848 75828 59020
rect 75862 58848 75868 59020
rect 75822 58836 75868 58848
rect 76480 59020 76526 59032
rect 76480 58848 76486 59020
rect 76520 58848 76526 59020
rect 77138 59020 77184 59032
rect 77138 58986 77144 59020
rect 76480 58836 76526 58848
rect 77124 58848 77144 58986
rect 77178 58986 77184 59020
rect 77796 59020 77842 59032
rect 77178 58848 77200 58986
rect 73260 57938 73280 58040
rect 72616 57856 72662 57868
rect 73274 57868 73280 57938
rect 73314 57938 73336 58040
rect 73932 58040 73978 58052
rect 73314 57868 73320 57938
rect 73274 57856 73320 57868
rect 73932 57868 73938 58040
rect 73972 57868 73978 58040
rect 75164 58020 75210 58032
rect 73932 57856 73978 57868
rect 74872 57874 75088 58020
rect 71300 57346 71346 57358
rect 71300 57174 71306 57346
rect 71340 57174 71346 57346
rect 71300 57162 71346 57174
rect 71958 57346 72004 57358
rect 71958 57174 71964 57346
rect 71998 57174 72004 57346
rect 71958 57162 72004 57174
rect 72616 57346 72662 57358
rect 72616 57174 72622 57346
rect 72656 57174 72662 57346
rect 72616 57162 72662 57174
rect 73274 57346 73320 57358
rect 73274 57174 73280 57346
rect 73314 57174 73320 57346
rect 73274 57162 73320 57174
rect 73932 57346 73978 57358
rect 73932 57174 73938 57346
rect 73972 57174 73978 57346
rect 73932 57162 73978 57174
rect 71300 56652 71346 56664
rect 71300 56480 71306 56652
rect 71340 56480 71346 56652
rect 71300 56468 71346 56480
rect 71958 56652 72004 56664
rect 71958 56480 71964 56652
rect 71998 56480 72004 56652
rect 71958 56468 72004 56480
rect 72616 56652 72662 56664
rect 72616 56480 72622 56652
rect 72656 56480 72662 56652
rect 72616 56468 72662 56480
rect 73274 56652 73320 56664
rect 73274 56480 73280 56652
rect 73314 56480 73320 56652
rect 73274 56468 73320 56480
rect 73932 56652 73978 56664
rect 73932 56480 73938 56652
rect 73972 56480 73978 56652
rect 73932 56468 73978 56480
rect 71300 55958 71346 55970
rect 71300 55786 71306 55958
rect 71340 55786 71346 55958
rect 71300 55774 71346 55786
rect 71958 55958 72004 55970
rect 71958 55786 71964 55958
rect 71998 55786 72004 55958
rect 71958 55774 72004 55786
rect 72616 55958 72662 55970
rect 72616 55786 72622 55958
rect 72656 55786 72662 55958
rect 72616 55774 72662 55786
rect 73274 55958 73320 55970
rect 73274 55786 73280 55958
rect 73314 55786 73320 55958
rect 73274 55774 73320 55786
rect 73932 55958 73978 55970
rect 73932 55786 73938 55958
rect 73972 55786 73978 55958
rect 73932 55774 73978 55786
rect 71008 55180 71224 55326
rect 74872 55306 74926 57874
rect 75010 55306 75088 57874
rect 75164 57848 75170 58020
rect 75204 57848 75210 58020
rect 75164 57836 75210 57848
rect 75822 58020 75868 58032
rect 75822 57848 75828 58020
rect 75862 57848 75868 58020
rect 75822 57836 75868 57848
rect 76480 58020 76526 58032
rect 76480 57848 76486 58020
rect 76520 57848 76526 58020
rect 77124 58020 77200 58848
rect 77796 58848 77802 59020
rect 77836 58848 77842 59020
rect 78722 58950 78938 59096
rect 79014 59034 79060 59046
rect 79014 58862 79020 59034
rect 79054 58862 79060 59034
rect 79014 58850 79060 58862
rect 79672 59034 79718 59046
rect 79672 58862 79678 59034
rect 79712 58862 79718 59034
rect 79672 58850 79718 58862
rect 80330 59034 80376 59046
rect 80330 58862 80336 59034
rect 80370 58862 80376 59034
rect 80988 59034 81034 59046
rect 80988 59000 80994 59034
rect 80330 58850 80376 58862
rect 80974 58862 80994 59000
rect 81028 59000 81034 59034
rect 81646 59034 81692 59046
rect 81028 58862 81050 59000
rect 77796 58836 77842 58848
rect 79014 58034 79060 58046
rect 77124 57918 77144 58020
rect 76480 57836 76526 57848
rect 77138 57848 77144 57918
rect 77178 57918 77200 58020
rect 77796 58020 77842 58032
rect 77178 57848 77184 57918
rect 77138 57836 77184 57848
rect 77796 57848 77802 58020
rect 77836 57848 77842 58020
rect 77796 57836 77842 57848
rect 78722 57888 78938 58034
rect 75164 57326 75210 57338
rect 75164 57154 75170 57326
rect 75204 57154 75210 57326
rect 75164 57142 75210 57154
rect 75822 57326 75868 57338
rect 75822 57154 75828 57326
rect 75862 57154 75868 57326
rect 75822 57142 75868 57154
rect 76480 57326 76526 57338
rect 76480 57154 76486 57326
rect 76520 57154 76526 57326
rect 76480 57142 76526 57154
rect 77138 57326 77184 57338
rect 77138 57154 77144 57326
rect 77178 57154 77184 57326
rect 77138 57142 77184 57154
rect 77796 57326 77842 57338
rect 77796 57154 77802 57326
rect 77836 57154 77842 57326
rect 77796 57142 77842 57154
rect 75164 56632 75210 56644
rect 75164 56460 75170 56632
rect 75204 56460 75210 56632
rect 75164 56448 75210 56460
rect 75822 56632 75868 56644
rect 75822 56460 75828 56632
rect 75862 56460 75868 56632
rect 75822 56448 75868 56460
rect 76480 56632 76526 56644
rect 76480 56460 76486 56632
rect 76520 56460 76526 56632
rect 76480 56448 76526 56460
rect 77138 56632 77184 56644
rect 77138 56460 77144 56632
rect 77178 56460 77184 56632
rect 77138 56448 77184 56460
rect 77796 56632 77842 56644
rect 77796 56460 77802 56632
rect 77836 56460 77842 56632
rect 77796 56448 77842 56460
rect 75164 55938 75210 55950
rect 75164 55766 75170 55938
rect 75204 55766 75210 55938
rect 75164 55754 75210 55766
rect 75822 55938 75868 55950
rect 75822 55766 75828 55938
rect 75862 55766 75868 55938
rect 75822 55754 75868 55766
rect 76480 55938 76526 55950
rect 76480 55766 76486 55938
rect 76520 55766 76526 55938
rect 76480 55754 76526 55766
rect 77138 55938 77184 55950
rect 77138 55766 77144 55938
rect 77178 55766 77184 55938
rect 77138 55754 77184 55766
rect 77796 55938 77842 55950
rect 77796 55766 77802 55938
rect 77836 55766 77842 55938
rect 77796 55754 77842 55766
rect 71300 55264 71346 55276
rect 71300 55092 71306 55264
rect 71340 55092 71346 55264
rect 71300 55080 71346 55092
rect 71958 55264 72004 55276
rect 71958 55092 71964 55264
rect 71998 55092 72004 55264
rect 71958 55080 72004 55092
rect 72616 55264 72662 55276
rect 72616 55092 72622 55264
rect 72656 55092 72662 55264
rect 73274 55264 73320 55276
rect 73274 55226 73280 55264
rect 72616 55080 72662 55092
rect 73260 55092 73280 55226
rect 73314 55226 73320 55264
rect 73932 55264 73978 55276
rect 73314 55092 73336 55226
rect 71304 54268 71350 54280
rect 71012 54122 71228 54268
rect 71012 51554 71066 54122
rect 71150 51554 71228 54122
rect 71304 54096 71310 54268
rect 71344 54096 71350 54268
rect 71304 54084 71350 54096
rect 71962 54268 72008 54280
rect 71962 54096 71968 54268
rect 72002 54096 72008 54268
rect 71962 54084 72008 54096
rect 72620 54268 72666 54280
rect 72620 54096 72626 54268
rect 72660 54096 72666 54268
rect 73260 54268 73336 55092
rect 73932 55092 73938 55264
rect 73972 55092 73978 55264
rect 74872 55160 75088 55306
rect 78722 55320 78776 57888
rect 78860 55320 78938 57888
rect 79014 57862 79020 58034
rect 79054 57862 79060 58034
rect 79014 57850 79060 57862
rect 79672 58034 79718 58046
rect 79672 57862 79678 58034
rect 79712 57862 79718 58034
rect 79672 57850 79718 57862
rect 80330 58034 80376 58046
rect 80330 57862 80336 58034
rect 80370 57862 80376 58034
rect 80974 58034 81050 58862
rect 81646 58862 81652 59034
rect 81686 58862 81692 59034
rect 81646 58850 81692 58862
rect 80974 57932 80994 58034
rect 80330 57850 80376 57862
rect 80988 57862 80994 57932
rect 81028 57932 81050 58034
rect 81646 58034 81692 58046
rect 81028 57862 81034 57932
rect 80988 57850 81034 57862
rect 81646 57862 81652 58034
rect 81686 57862 81692 58034
rect 81646 57850 81692 57862
rect 79014 57340 79060 57352
rect 79014 57168 79020 57340
rect 79054 57168 79060 57340
rect 79014 57156 79060 57168
rect 79672 57340 79718 57352
rect 79672 57168 79678 57340
rect 79712 57168 79718 57340
rect 79672 57156 79718 57168
rect 80330 57340 80376 57352
rect 80330 57168 80336 57340
rect 80370 57168 80376 57340
rect 80330 57156 80376 57168
rect 80988 57340 81034 57352
rect 80988 57168 80994 57340
rect 81028 57168 81034 57340
rect 80988 57156 81034 57168
rect 81646 57340 81692 57352
rect 81646 57168 81652 57340
rect 81686 57168 81692 57340
rect 81646 57156 81692 57168
rect 79014 56646 79060 56658
rect 79014 56474 79020 56646
rect 79054 56474 79060 56646
rect 79014 56462 79060 56474
rect 79672 56646 79718 56658
rect 79672 56474 79678 56646
rect 79712 56474 79718 56646
rect 79672 56462 79718 56474
rect 80330 56646 80376 56658
rect 80330 56474 80336 56646
rect 80370 56474 80376 56646
rect 80330 56462 80376 56474
rect 80988 56646 81034 56658
rect 80988 56474 80994 56646
rect 81028 56474 81034 56646
rect 80988 56462 81034 56474
rect 81646 56646 81692 56658
rect 81646 56474 81652 56646
rect 81686 56474 81692 56646
rect 81646 56462 81692 56474
rect 79014 55952 79060 55964
rect 79014 55780 79020 55952
rect 79054 55780 79060 55952
rect 79014 55768 79060 55780
rect 79672 55952 79718 55964
rect 79672 55780 79678 55952
rect 79712 55780 79718 55952
rect 79672 55768 79718 55780
rect 80330 55952 80376 55964
rect 80330 55780 80336 55952
rect 80370 55780 80376 55952
rect 80330 55768 80376 55780
rect 80988 55952 81034 55964
rect 80988 55780 80994 55952
rect 81028 55780 81034 55952
rect 80988 55768 81034 55780
rect 81646 55952 81692 55964
rect 81646 55780 81652 55952
rect 81686 55780 81692 55952
rect 81646 55768 81692 55780
rect 75164 55244 75210 55256
rect 73932 55080 73978 55092
rect 75164 55072 75170 55244
rect 75204 55072 75210 55244
rect 75164 55060 75210 55072
rect 75822 55244 75868 55256
rect 75822 55072 75828 55244
rect 75862 55072 75868 55244
rect 75822 55060 75868 55072
rect 76480 55244 76526 55256
rect 76480 55072 76486 55244
rect 76520 55072 76526 55244
rect 77138 55244 77184 55256
rect 77138 55206 77144 55244
rect 76480 55060 76526 55072
rect 77124 55072 77144 55206
rect 77178 55206 77184 55244
rect 77796 55244 77842 55256
rect 77178 55072 77200 55206
rect 73260 54158 73284 54268
rect 72620 54084 72666 54096
rect 73278 54096 73284 54158
rect 73318 54158 73336 54268
rect 73936 54268 73982 54280
rect 73318 54096 73324 54158
rect 73278 54084 73324 54096
rect 73936 54096 73942 54268
rect 73976 54096 73982 54268
rect 75168 54248 75214 54260
rect 73936 54084 73982 54096
rect 74876 54102 75092 54248
rect 71304 53574 71350 53586
rect 71304 53402 71310 53574
rect 71344 53402 71350 53574
rect 71304 53390 71350 53402
rect 71962 53574 72008 53586
rect 71962 53402 71968 53574
rect 72002 53402 72008 53574
rect 71962 53390 72008 53402
rect 72620 53574 72666 53586
rect 72620 53402 72626 53574
rect 72660 53402 72666 53574
rect 72620 53390 72666 53402
rect 73278 53574 73324 53586
rect 73278 53402 73284 53574
rect 73318 53402 73324 53574
rect 73278 53390 73324 53402
rect 73936 53574 73982 53586
rect 73936 53402 73942 53574
rect 73976 53402 73982 53574
rect 73936 53390 73982 53402
rect 71304 52880 71350 52892
rect 71304 52708 71310 52880
rect 71344 52708 71350 52880
rect 71304 52696 71350 52708
rect 71962 52880 72008 52892
rect 71962 52708 71968 52880
rect 72002 52708 72008 52880
rect 71962 52696 72008 52708
rect 72620 52880 72666 52892
rect 72620 52708 72626 52880
rect 72660 52708 72666 52880
rect 72620 52696 72666 52708
rect 73278 52880 73324 52892
rect 73278 52708 73284 52880
rect 73318 52708 73324 52880
rect 73278 52696 73324 52708
rect 73936 52880 73982 52892
rect 73936 52708 73942 52880
rect 73976 52708 73982 52880
rect 73936 52696 73982 52708
rect 71304 52186 71350 52198
rect 71304 52014 71310 52186
rect 71344 52014 71350 52186
rect 71304 52002 71350 52014
rect 71962 52186 72008 52198
rect 71962 52014 71968 52186
rect 72002 52014 72008 52186
rect 71962 52002 72008 52014
rect 72620 52186 72666 52198
rect 72620 52014 72626 52186
rect 72660 52014 72666 52186
rect 72620 52002 72666 52014
rect 73278 52186 73324 52198
rect 73278 52014 73284 52186
rect 73318 52014 73324 52186
rect 73278 52002 73324 52014
rect 73936 52186 73982 52198
rect 73936 52014 73942 52186
rect 73976 52014 73982 52186
rect 73936 52002 73982 52014
rect 71012 51408 71228 51554
rect 74876 51534 74930 54102
rect 75014 51534 75092 54102
rect 75168 54076 75174 54248
rect 75208 54076 75214 54248
rect 75168 54064 75214 54076
rect 75826 54248 75872 54260
rect 75826 54076 75832 54248
rect 75866 54076 75872 54248
rect 75826 54064 75872 54076
rect 76484 54248 76530 54260
rect 76484 54076 76490 54248
rect 76524 54076 76530 54248
rect 77124 54248 77200 55072
rect 77796 55072 77802 55244
rect 77836 55072 77842 55244
rect 78722 55174 78938 55320
rect 79014 55258 79060 55270
rect 79014 55086 79020 55258
rect 79054 55086 79060 55258
rect 79014 55074 79060 55086
rect 79672 55258 79718 55270
rect 79672 55086 79678 55258
rect 79712 55086 79718 55258
rect 79672 55074 79718 55086
rect 80330 55258 80376 55270
rect 80330 55086 80336 55258
rect 80370 55086 80376 55258
rect 80988 55258 81034 55270
rect 80988 55220 80994 55258
rect 80330 55074 80376 55086
rect 80974 55086 80994 55220
rect 81028 55220 81034 55258
rect 81646 55258 81692 55270
rect 81028 55086 81050 55220
rect 77796 55060 77842 55072
rect 79018 54262 79064 54274
rect 77124 54138 77148 54248
rect 76484 54064 76530 54076
rect 77142 54076 77148 54138
rect 77182 54138 77200 54248
rect 77800 54248 77846 54260
rect 77182 54076 77188 54138
rect 77142 54064 77188 54076
rect 77800 54076 77806 54248
rect 77840 54076 77846 54248
rect 77800 54064 77846 54076
rect 78726 54116 78942 54262
rect 75168 53554 75214 53566
rect 75168 53382 75174 53554
rect 75208 53382 75214 53554
rect 75168 53370 75214 53382
rect 75826 53554 75872 53566
rect 75826 53382 75832 53554
rect 75866 53382 75872 53554
rect 75826 53370 75872 53382
rect 76484 53554 76530 53566
rect 76484 53382 76490 53554
rect 76524 53382 76530 53554
rect 76484 53370 76530 53382
rect 77142 53554 77188 53566
rect 77142 53382 77148 53554
rect 77182 53382 77188 53554
rect 77142 53370 77188 53382
rect 77800 53554 77846 53566
rect 77800 53382 77806 53554
rect 77840 53382 77846 53554
rect 77800 53370 77846 53382
rect 75168 52860 75214 52872
rect 75168 52688 75174 52860
rect 75208 52688 75214 52860
rect 75168 52676 75214 52688
rect 75826 52860 75872 52872
rect 75826 52688 75832 52860
rect 75866 52688 75872 52860
rect 75826 52676 75872 52688
rect 76484 52860 76530 52872
rect 76484 52688 76490 52860
rect 76524 52688 76530 52860
rect 76484 52676 76530 52688
rect 77142 52860 77188 52872
rect 77142 52688 77148 52860
rect 77182 52688 77188 52860
rect 77142 52676 77188 52688
rect 77800 52860 77846 52872
rect 77800 52688 77806 52860
rect 77840 52688 77846 52860
rect 77800 52676 77846 52688
rect 75168 52166 75214 52178
rect 75168 51994 75174 52166
rect 75208 51994 75214 52166
rect 75168 51982 75214 51994
rect 75826 52166 75872 52178
rect 75826 51994 75832 52166
rect 75866 51994 75872 52166
rect 75826 51982 75872 51994
rect 76484 52166 76530 52178
rect 76484 51994 76490 52166
rect 76524 51994 76530 52166
rect 76484 51982 76530 51994
rect 77142 52166 77188 52178
rect 77142 51994 77148 52166
rect 77182 51994 77188 52166
rect 77142 51982 77188 51994
rect 77800 52166 77846 52178
rect 77800 51994 77806 52166
rect 77840 51994 77846 52166
rect 77800 51982 77846 51994
rect 71304 51492 71350 51504
rect 71304 51320 71310 51492
rect 71344 51320 71350 51492
rect 71304 51308 71350 51320
rect 71962 51492 72008 51504
rect 71962 51320 71968 51492
rect 72002 51320 72008 51492
rect 71962 51308 72008 51320
rect 72620 51492 72666 51504
rect 72620 51320 72626 51492
rect 72660 51320 72666 51492
rect 72620 51308 72666 51320
rect 73278 51492 73324 51504
rect 73278 51320 73284 51492
rect 73318 51320 73324 51492
rect 73278 51308 73324 51320
rect 73936 51492 73982 51504
rect 73936 51320 73942 51492
rect 73976 51320 73982 51492
rect 74876 51388 75092 51534
rect 78726 51548 78780 54116
rect 78864 51548 78942 54116
rect 79018 54090 79024 54262
rect 79058 54090 79064 54262
rect 79018 54078 79064 54090
rect 79676 54262 79722 54274
rect 79676 54090 79682 54262
rect 79716 54090 79722 54262
rect 79676 54078 79722 54090
rect 80334 54262 80380 54274
rect 80334 54090 80340 54262
rect 80374 54090 80380 54262
rect 80974 54262 81050 55086
rect 81646 55086 81652 55258
rect 81686 55086 81692 55258
rect 81646 55074 81692 55086
rect 81894 54946 81928 54954
rect 81894 54918 82128 54946
rect 81896 54890 82128 54918
rect 80974 54152 80998 54262
rect 80334 54078 80380 54090
rect 80992 54090 80998 54152
rect 81032 54152 81050 54262
rect 81650 54262 81696 54274
rect 81032 54090 81038 54152
rect 80992 54078 81038 54090
rect 81650 54090 81656 54262
rect 81690 54090 81696 54262
rect 81896 54218 81924 54890
rect 82048 54294 82128 54890
rect 83280 54294 83328 54300
rect 82048 54218 83332 54294
rect 81896 54146 83332 54218
rect 81896 54108 82128 54146
rect 81650 54078 81696 54090
rect 83004 54070 83090 54146
rect 83280 54105 83328 54146
rect 83272 54099 86344 54105
rect 82966 53912 82976 54070
rect 83164 53912 83174 54070
rect 83272 54065 83303 54099
rect 83337 54065 83399 54099
rect 83433 54065 83495 54099
rect 83529 54065 83591 54099
rect 83625 54065 83687 54099
rect 83721 54065 83783 54099
rect 83817 54065 83879 54099
rect 83913 54065 83975 54099
rect 84009 54065 84071 54099
rect 84105 54065 84167 54099
rect 84201 54065 84263 54099
rect 84297 54065 84359 54099
rect 84393 54065 84455 54099
rect 84489 54065 84551 54099
rect 84585 54065 84647 54099
rect 84681 54065 84743 54099
rect 84777 54065 84839 54099
rect 84873 54065 84935 54099
rect 84969 54065 85031 54099
rect 85065 54065 85127 54099
rect 85161 54065 85223 54099
rect 85257 54065 85319 54099
rect 85353 54065 85415 54099
rect 85449 54065 85511 54099
rect 85545 54065 85607 54099
rect 85641 54065 85703 54099
rect 85737 54065 85799 54099
rect 85833 54065 85895 54099
rect 85929 54065 85991 54099
rect 86025 54065 86087 54099
rect 86121 54065 86183 54099
rect 86217 54065 86279 54099
rect 86313 54065 86344 54099
rect 83272 54059 86344 54065
rect 83280 54031 83328 54059
rect 83272 54003 86344 54031
rect 83272 53969 83404 54003
rect 83438 53969 83476 54003
rect 83510 53969 83882 54003
rect 83916 53969 84368 54003
rect 84402 53969 84440 54003
rect 84474 53969 84512 54003
rect 84546 53969 84836 54003
rect 84870 53969 84908 54003
rect 84942 53969 84980 54003
rect 85014 53969 85375 54003
rect 85409 53969 85447 54003
rect 85481 53969 85519 54003
rect 85553 53969 85726 54003
rect 85760 53969 85798 54003
rect 85832 53969 85870 54003
rect 85904 53969 86032 54003
rect 86066 53969 86104 54003
rect 86138 53969 86176 54003
rect 86210 53969 86344 54003
rect 83272 53957 86344 53969
rect 83370 53700 83460 53706
rect 83370 53682 83382 53700
rect 79018 53568 79064 53580
rect 79018 53396 79024 53568
rect 79058 53396 79064 53568
rect 79018 53384 79064 53396
rect 79676 53568 79722 53580
rect 79676 53396 79682 53568
rect 79716 53396 79722 53568
rect 79676 53384 79722 53396
rect 80334 53568 80380 53580
rect 80334 53396 80340 53568
rect 80374 53396 80380 53568
rect 80334 53384 80380 53396
rect 80992 53568 81038 53580
rect 80992 53396 80998 53568
rect 81032 53396 81038 53568
rect 80992 53384 81038 53396
rect 81650 53568 81696 53580
rect 81650 53396 81656 53568
rect 81690 53396 81696 53568
rect 82548 53468 82558 53658
rect 82674 53584 82684 53658
rect 83236 53652 83382 53682
rect 83370 53640 83382 53652
rect 83448 53640 83460 53700
rect 83675 53692 83733 53698
rect 83675 53658 83687 53692
rect 83721 53689 83733 53692
rect 84155 53692 84213 53698
rect 84155 53689 84167 53692
rect 83721 53661 84167 53689
rect 83721 53658 83733 53661
rect 83675 53652 83733 53658
rect 84155 53658 84167 53661
rect 84201 53689 84213 53692
rect 85211 53692 85269 53698
rect 85211 53689 85223 53692
rect 84201 53661 85223 53689
rect 84201 53658 84213 53661
rect 84155 53652 84213 53658
rect 85211 53658 85223 53661
rect 85257 53658 85269 53692
rect 85211 53652 85269 53658
rect 83370 53634 83460 53640
rect 86258 53630 86328 53636
rect 83964 53606 84026 53618
rect 83964 53584 83970 53606
rect 82674 53550 83970 53584
rect 84020 53550 84026 53606
rect 86258 53586 86270 53630
rect 86316 53590 86440 53630
rect 86316 53586 86328 53590
rect 86258 53580 86328 53586
rect 82674 53538 84026 53550
rect 82674 53528 83248 53538
rect 82674 53468 82684 53528
rect 83858 53498 83932 53504
rect 82998 53424 83008 53498
rect 83100 53492 83110 53498
rect 83100 53490 83758 53492
rect 83858 53490 83870 53498
rect 83100 53460 83870 53490
rect 83920 53460 83932 53498
rect 83100 53454 83932 53460
rect 83100 53452 83880 53454
rect 83100 53450 83758 53452
rect 83100 53424 83110 53450
rect 81650 53384 81696 53396
rect 83272 53381 86344 53393
rect 83272 53347 83390 53381
rect 83424 53347 83462 53381
rect 83496 53347 83534 53381
rect 83568 53347 83718 53381
rect 83752 53347 83790 53381
rect 83824 53347 84710 53381
rect 84744 53347 84782 53381
rect 84816 53347 84854 53381
rect 84888 53347 85504 53381
rect 85538 53347 85576 53381
rect 85610 53347 85648 53381
rect 85682 53347 86025 53381
rect 86059 53347 86097 53381
rect 86131 53347 86169 53381
rect 86203 53347 86344 53381
rect 83272 53319 86344 53347
rect 86140 53291 86212 53319
rect 83272 53285 86344 53291
rect 83272 53251 83303 53285
rect 83337 53251 83399 53285
rect 83433 53251 83495 53285
rect 83529 53251 83591 53285
rect 83625 53251 83687 53285
rect 83721 53251 83783 53285
rect 83817 53251 83879 53285
rect 83913 53251 83975 53285
rect 84009 53251 84071 53285
rect 84105 53251 84167 53285
rect 84201 53251 84263 53285
rect 84297 53251 84359 53285
rect 84393 53251 84455 53285
rect 84489 53251 84551 53285
rect 84585 53251 84647 53285
rect 84681 53251 84743 53285
rect 84777 53251 84839 53285
rect 84873 53251 84935 53285
rect 84969 53251 85031 53285
rect 85065 53251 85127 53285
rect 85161 53251 85223 53285
rect 85257 53251 85319 53285
rect 85353 53251 85415 53285
rect 85449 53251 85511 53285
rect 85545 53251 85607 53285
rect 85641 53251 85703 53285
rect 85737 53251 85799 53285
rect 85833 53251 85895 53285
rect 85929 53251 85991 53285
rect 86025 53251 86087 53285
rect 86121 53251 86183 53285
rect 86217 53251 86279 53285
rect 86313 53251 86344 53285
rect 83272 53245 86344 53251
rect 79018 52874 79064 52886
rect 79018 52702 79024 52874
rect 79058 52702 79064 52874
rect 79018 52690 79064 52702
rect 79676 52874 79722 52886
rect 79676 52702 79682 52874
rect 79716 52702 79722 52874
rect 79676 52690 79722 52702
rect 80334 52874 80380 52886
rect 80334 52702 80340 52874
rect 80374 52702 80380 52874
rect 80334 52690 80380 52702
rect 80992 52874 81038 52886
rect 80992 52702 80998 52874
rect 81032 52702 81038 52874
rect 80992 52690 81038 52702
rect 81650 52874 81696 52886
rect 81650 52702 81656 52874
rect 81690 52702 81696 52874
rect 81650 52690 81696 52702
rect 79018 52180 79064 52192
rect 79018 52008 79024 52180
rect 79058 52008 79064 52180
rect 79018 51996 79064 52008
rect 79676 52180 79722 52192
rect 79676 52008 79682 52180
rect 79716 52008 79722 52180
rect 79676 51996 79722 52008
rect 80334 52180 80380 52192
rect 80334 52008 80340 52180
rect 80374 52008 80380 52180
rect 80334 51996 80380 52008
rect 80992 52180 81038 52192
rect 80992 52008 80998 52180
rect 81032 52008 81038 52180
rect 80992 51996 81038 52008
rect 81650 52180 81696 52192
rect 81650 52008 81656 52180
rect 81690 52008 81696 52180
rect 81650 51996 81696 52008
rect 86140 51866 86212 53245
rect 88266 51866 88276 51918
rect 86140 51792 88276 51866
rect 86140 51778 86212 51792
rect 88266 51730 88276 51792
rect 88474 51730 88484 51918
rect 75168 51472 75214 51484
rect 73936 51308 73982 51320
rect 75168 51300 75174 51472
rect 75208 51300 75214 51472
rect 75168 51288 75214 51300
rect 75826 51472 75872 51484
rect 75826 51300 75832 51472
rect 75866 51300 75872 51472
rect 75826 51288 75872 51300
rect 76484 51472 76530 51484
rect 76484 51300 76490 51472
rect 76524 51300 76530 51472
rect 76484 51288 76530 51300
rect 77142 51472 77188 51484
rect 77142 51300 77148 51472
rect 77182 51300 77188 51472
rect 77142 51288 77188 51300
rect 77800 51472 77846 51484
rect 77800 51300 77806 51472
rect 77840 51300 77846 51472
rect 78726 51402 78942 51548
rect 79018 51486 79064 51498
rect 79018 51314 79024 51486
rect 79058 51314 79064 51486
rect 79018 51302 79064 51314
rect 79676 51486 79722 51498
rect 79676 51314 79682 51486
rect 79716 51314 79722 51486
rect 79676 51302 79722 51314
rect 80334 51486 80380 51498
rect 80334 51314 80340 51486
rect 80374 51314 80380 51486
rect 80334 51302 80380 51314
rect 80992 51486 81038 51498
rect 80992 51314 80998 51486
rect 81032 51314 81038 51486
rect 80992 51302 81038 51314
rect 81650 51486 81696 51498
rect 81650 51314 81656 51486
rect 81690 51314 81696 51486
rect 81650 51302 81696 51314
rect 77800 51288 77846 51300
rect 77322 51022 77690 51054
rect 77294 51008 77690 51022
rect 77294 50850 77384 51008
rect 77634 50850 77690 51008
rect 77294 50798 77690 50850
rect 57128 50414 57324 50420
rect 59872 49850 68038 50432
rect 59906 49814 60318 49850
rect 42314 49796 42510 49802
rect 42314 49762 42326 49796
rect 42498 49762 42510 49796
rect 42314 49756 42510 49762
rect 43008 49796 43204 49802
rect 43008 49762 43020 49796
rect 43192 49762 43204 49796
rect 43008 49756 43204 49762
rect 43702 49796 43898 49802
rect 43702 49762 43714 49796
rect 43886 49762 43898 49796
rect 43702 49756 43898 49762
rect 44396 49796 44592 49802
rect 44396 49762 44408 49796
rect 44580 49762 44592 49796
rect 44396 49756 44592 49762
rect 45090 49796 45286 49802
rect 45090 49762 45102 49796
rect 45274 49762 45286 49796
rect 45090 49756 45286 49762
rect 46308 49796 46504 49802
rect 46308 49762 46320 49796
rect 46492 49762 46504 49796
rect 46308 49756 46504 49762
rect 47002 49796 47198 49802
rect 47002 49762 47014 49796
rect 47186 49762 47198 49796
rect 47002 49756 47198 49762
rect 47696 49796 47892 49802
rect 47696 49762 47708 49796
rect 47880 49762 47892 49796
rect 47696 49756 47892 49762
rect 48390 49796 48586 49802
rect 48390 49762 48402 49796
rect 48574 49762 48586 49796
rect 48390 49756 48586 49762
rect 49084 49796 49280 49802
rect 49084 49762 49096 49796
rect 49268 49762 49280 49796
rect 49084 49756 49280 49762
rect 50330 49796 50526 49802
rect 50330 49762 50342 49796
rect 50514 49762 50526 49796
rect 50330 49756 50526 49762
rect 51024 49796 51220 49802
rect 51024 49762 51036 49796
rect 51208 49762 51220 49796
rect 51024 49756 51220 49762
rect 51718 49796 51914 49802
rect 51718 49762 51730 49796
rect 51902 49762 51914 49796
rect 51718 49756 51914 49762
rect 52412 49796 52608 49802
rect 52412 49762 52424 49796
rect 52596 49762 52608 49796
rect 52412 49756 52608 49762
rect 53106 49796 53302 49802
rect 53106 49762 53118 49796
rect 53290 49762 53302 49796
rect 53106 49756 53302 49762
rect 54352 49796 54548 49802
rect 54352 49762 54364 49796
rect 54536 49762 54548 49796
rect 54352 49756 54548 49762
rect 55046 49796 55242 49802
rect 55046 49762 55058 49796
rect 55230 49762 55242 49796
rect 55046 49756 55242 49762
rect 55740 49796 55936 49802
rect 55740 49762 55752 49796
rect 55924 49762 55936 49796
rect 55740 49756 55936 49762
rect 56434 49796 56630 49802
rect 56434 49762 56446 49796
rect 56618 49762 56630 49796
rect 56434 49756 56630 49762
rect 57128 49796 57324 49802
rect 57128 49762 57140 49796
rect 57312 49762 57324 49796
rect 57128 49756 57324 49762
rect 19532 49038 19728 49044
rect 19532 49004 19544 49038
rect 19716 49004 19728 49038
rect 926 48988 1122 48994
rect 926 48954 938 48988
rect 1110 48954 1122 48988
rect 926 48948 1122 48954
rect 1620 48988 1816 48994
rect 1620 48954 1632 48988
rect 1804 48954 1816 48988
rect 1620 48948 1816 48954
rect 2314 48988 2510 48994
rect 6268 48990 6464 48996
rect 2314 48954 2326 48988
rect 2498 48954 2510 48988
rect 2314 48948 2510 48954
rect 3594 48984 3790 48990
rect 3594 48950 3606 48984
rect 3778 48950 3790 48984
rect 3594 48944 3790 48950
rect 4288 48984 4484 48990
rect 4288 48950 4300 48984
rect 4472 48950 4484 48984
rect 4288 48944 4484 48950
rect 4982 48984 5178 48990
rect 4982 48950 4994 48984
rect 5166 48950 5178 48984
rect 6268 48956 6280 48990
rect 6452 48956 6464 48990
rect 6268 48950 6464 48956
rect 6962 48990 7158 48996
rect 6962 48956 6974 48990
rect 7146 48956 7158 48990
rect 6962 48950 7158 48956
rect 7656 48990 7852 48996
rect 7656 48956 7668 48990
rect 7840 48956 7852 48990
rect 7656 48950 7852 48956
rect 8914 48990 9110 48996
rect 8914 48956 8926 48990
rect 9098 48956 9110 48990
rect 8914 48950 9110 48956
rect 9608 48990 9804 48996
rect 9608 48956 9620 48990
rect 9792 48956 9804 48990
rect 9608 48950 9804 48956
rect 10302 48990 10498 48996
rect 14222 48990 14418 48996
rect 10302 48956 10314 48990
rect 10486 48956 10498 48990
rect 10302 48950 10498 48956
rect 11568 48984 11764 48990
rect 11568 48950 11580 48984
rect 11752 48950 11764 48984
rect 4982 48944 5178 48950
rect 11568 48944 11764 48950
rect 12262 48984 12458 48990
rect 12262 48950 12274 48984
rect 12446 48950 12458 48984
rect 12262 48944 12458 48950
rect 12956 48984 13152 48990
rect 12956 48950 12968 48984
rect 13140 48950 13152 48984
rect 14222 48956 14234 48990
rect 14406 48956 14418 48990
rect 14222 48950 14418 48956
rect 14916 48990 15112 48996
rect 14916 48956 14928 48990
rect 15100 48956 15112 48990
rect 14916 48950 15112 48956
rect 15610 48990 15806 48996
rect 15610 48956 15622 48990
rect 15794 48956 15806 48990
rect 15610 48950 15806 48956
rect 16848 48994 17044 49000
rect 16848 48960 16860 48994
rect 17032 48960 17044 48994
rect 16848 48954 17044 48960
rect 17542 48994 17738 49000
rect 17542 48960 17554 48994
rect 17726 48960 17738 48994
rect 17542 48954 17738 48960
rect 18236 48994 18432 49000
rect 19532 48998 19728 49004
rect 20226 49038 20422 49044
rect 20226 49004 20238 49038
rect 20410 49004 20422 49038
rect 20226 48998 20422 49004
rect 18236 48960 18248 48994
rect 18420 48960 18432 48994
rect 18236 48954 18432 48960
rect 12956 48944 13152 48950
rect 20654 48728 20766 48758
rect 20654 48694 20690 48728
rect 20742 48694 20766 48728
rect 20654 48666 20766 48694
rect 8346 48546 8560 48558
rect 5686 48470 5934 48482
rect 3052 48436 3282 48448
rect 3052 48386 3058 48436
rect 2368 48336 3058 48386
rect 926 48330 1122 48336
rect 926 48296 938 48330
rect 1110 48296 1122 48330
rect 926 48290 1122 48296
rect 1620 48330 1816 48336
rect 1620 48296 1632 48330
rect 1804 48296 1816 48330
rect 1620 48290 1816 48296
rect 2314 48330 3058 48336
rect 2314 48296 2326 48330
rect 2498 48296 3058 48330
rect 2314 48290 3058 48296
rect 2368 48226 3058 48290
rect 3052 48082 3058 48226
rect 3276 48082 3282 48436
rect 5686 48386 5692 48470
rect 5078 48332 5692 48386
rect 3594 48326 3790 48332
rect 3594 48292 3606 48326
rect 3778 48292 3790 48326
rect 3594 48286 3790 48292
rect 4288 48326 4484 48332
rect 4288 48292 4300 48326
rect 4472 48292 4484 48326
rect 4288 48286 4484 48292
rect 4982 48326 5692 48332
rect 4982 48292 4994 48326
rect 5166 48292 5692 48326
rect 4982 48286 5692 48292
rect 5078 48218 5692 48286
rect 5686 48108 5692 48218
rect 5928 48108 5934 48470
rect 8346 48428 8352 48546
rect 7720 48338 8352 48428
rect 6268 48332 6464 48338
rect 6268 48298 6280 48332
rect 6452 48298 6464 48332
rect 6268 48292 6464 48298
rect 6962 48332 7158 48338
rect 6962 48298 6974 48332
rect 7146 48298 7158 48332
rect 6962 48292 7158 48298
rect 7656 48332 8352 48338
rect 7656 48298 7668 48332
rect 7840 48298 8352 48332
rect 7656 48292 8352 48298
rect 7720 48192 8352 48292
rect 5686 48096 5934 48108
rect 3052 48070 3282 48082
rect 8346 48058 8352 48192
rect 8554 48058 8560 48546
rect 18838 48528 19060 48540
rect 13672 48494 13852 48506
rect 11022 48462 11252 48474
rect 11022 48376 11028 48462
rect 10380 48338 11028 48376
rect 8914 48332 9110 48338
rect 8914 48298 8926 48332
rect 9098 48298 9110 48332
rect 8914 48292 9110 48298
rect 9608 48332 9804 48338
rect 9608 48298 9620 48332
rect 9792 48298 9804 48332
rect 9608 48292 9804 48298
rect 10302 48332 11028 48338
rect 10302 48298 10314 48332
rect 10486 48298 11028 48332
rect 10302 48292 11028 48298
rect 10380 48184 11028 48292
rect 8346 48046 8560 48058
rect 11022 48024 11028 48184
rect 11246 48024 11252 48462
rect 13672 48368 13678 48494
rect 12988 48332 13678 48368
rect 11568 48326 11764 48332
rect 11568 48292 11580 48326
rect 11752 48292 11764 48326
rect 11568 48286 11764 48292
rect 12262 48326 12458 48332
rect 12262 48292 12274 48326
rect 12446 48292 12458 48326
rect 12262 48286 12458 48292
rect 12956 48326 13678 48332
rect 12956 48292 12968 48326
rect 13140 48292 13678 48326
rect 12956 48286 13678 48292
rect 12988 48250 13678 48286
rect 13672 48066 13678 48250
rect 13846 48066 13852 48494
rect 16288 48436 16554 48448
rect 16288 48394 16294 48436
rect 15664 48338 16294 48394
rect 14222 48332 14418 48338
rect 14222 48298 14234 48332
rect 14406 48298 14418 48332
rect 14222 48292 14418 48298
rect 14916 48332 15112 48338
rect 14916 48298 14928 48332
rect 15100 48298 15112 48332
rect 14916 48292 15112 48298
rect 15610 48332 16294 48338
rect 15610 48298 15622 48332
rect 15794 48298 16294 48332
rect 15610 48292 16294 48298
rect 15664 48276 16294 48292
rect 16288 48166 16294 48276
rect 16548 48166 16554 48436
rect 18838 48418 18844 48528
rect 18290 48342 18844 48418
rect 16848 48336 17044 48342
rect 16848 48302 16860 48336
rect 17032 48302 17044 48336
rect 16848 48296 17044 48302
rect 17542 48336 17738 48342
rect 17542 48302 17554 48336
rect 17726 48302 17738 48336
rect 17542 48296 17738 48302
rect 18236 48336 18844 48342
rect 18236 48302 18248 48336
rect 18420 48302 18844 48336
rect 18236 48296 18844 48302
rect 18290 48260 18844 48296
rect 18838 48182 18844 48260
rect 19054 48182 19060 48528
rect 19532 48380 19728 48386
rect 19532 48346 19544 48380
rect 19716 48346 19728 48380
rect 19532 48340 19728 48346
rect 20226 48380 20422 48386
rect 20226 48346 20238 48380
rect 20410 48346 20422 48380
rect 20226 48340 20422 48346
rect 18838 48170 19060 48182
rect 16288 48154 16554 48166
rect 13672 48054 13852 48066
rect 11022 48012 11252 48024
rect 19532 47722 19728 47728
rect 19532 47688 19544 47722
rect 19716 47688 19728 47722
rect 926 47672 1122 47678
rect 926 47638 938 47672
rect 1110 47638 1122 47672
rect 926 47632 1122 47638
rect 1620 47672 1816 47678
rect 1620 47638 1632 47672
rect 1804 47638 1816 47672
rect 1620 47632 1816 47638
rect 2314 47672 2510 47678
rect 6268 47674 6464 47680
rect 2314 47638 2326 47672
rect 2498 47638 2510 47672
rect 2314 47632 2510 47638
rect 3594 47668 3790 47674
rect 3594 47634 3606 47668
rect 3778 47634 3790 47668
rect 3594 47628 3790 47634
rect 4288 47668 4484 47674
rect 4288 47634 4300 47668
rect 4472 47634 4484 47668
rect 4288 47628 4484 47634
rect 4982 47668 5178 47674
rect 4982 47634 4994 47668
rect 5166 47634 5178 47668
rect 6268 47640 6280 47674
rect 6452 47640 6464 47674
rect 6268 47634 6464 47640
rect 6962 47674 7158 47680
rect 6962 47640 6974 47674
rect 7146 47640 7158 47674
rect 6962 47634 7158 47640
rect 7656 47674 7852 47680
rect 7656 47640 7668 47674
rect 7840 47640 7852 47674
rect 7656 47634 7852 47640
rect 8914 47674 9110 47680
rect 8914 47640 8926 47674
rect 9098 47640 9110 47674
rect 8914 47634 9110 47640
rect 9608 47674 9804 47680
rect 9608 47640 9620 47674
rect 9792 47640 9804 47674
rect 9608 47634 9804 47640
rect 10302 47674 10498 47680
rect 14222 47674 14418 47680
rect 10302 47640 10314 47674
rect 10486 47640 10498 47674
rect 10302 47634 10498 47640
rect 11568 47668 11764 47674
rect 11568 47634 11580 47668
rect 11752 47634 11764 47668
rect 4982 47628 5178 47634
rect 11568 47628 11764 47634
rect 12262 47668 12458 47674
rect 12262 47634 12274 47668
rect 12446 47634 12458 47668
rect 12262 47628 12458 47634
rect 12956 47668 13152 47674
rect 12956 47634 12968 47668
rect 13140 47634 13152 47668
rect 14222 47640 14234 47674
rect 14406 47640 14418 47674
rect 14222 47634 14418 47640
rect 14916 47674 15112 47680
rect 14916 47640 14928 47674
rect 15100 47640 15112 47674
rect 14916 47634 15112 47640
rect 15610 47674 15806 47680
rect 15610 47640 15622 47674
rect 15794 47640 15806 47674
rect 15610 47634 15806 47640
rect 16848 47678 17044 47684
rect 16848 47644 16860 47678
rect 17032 47644 17044 47678
rect 16848 47638 17044 47644
rect 17542 47678 17738 47684
rect 17542 47644 17554 47678
rect 17726 47644 17738 47678
rect 17542 47638 17738 47644
rect 18236 47678 18432 47684
rect 19532 47682 19728 47688
rect 20226 47722 20422 47728
rect 20226 47688 20238 47722
rect 20410 47688 20422 47722
rect 20226 47682 20422 47688
rect 18236 47644 18248 47678
rect 18420 47644 18432 47678
rect 18236 47638 18432 47644
rect 12956 47628 13152 47634
rect 2460 47334 4416 47400
rect 2460 47258 2730 47334
rect 4298 47258 4416 47334
rect 2460 47210 4416 47258
rect 9038 47394 10634 47430
rect 9038 47266 9218 47394
rect 10514 47266 10634 47394
rect 9038 47202 10634 47266
rect 14164 47360 15696 47416
rect 14164 47244 14392 47360
rect 15472 47244 15696 47360
rect 14164 47188 15696 47244
rect 16962 47394 18414 47434
rect 16962 47292 17118 47394
rect 18328 47292 18414 47394
rect 16962 47206 18414 47292
rect 19406 47364 20524 47412
rect 19406 47256 19582 47364
rect 20426 47256 20524 47364
rect 19406 47190 20524 47256
rect 21354 46432 21634 49318
rect 42314 49138 42510 49144
rect 42314 49104 42326 49138
rect 42498 49104 42510 49138
rect 42314 49098 42510 49104
rect 43008 49138 43204 49144
rect 43008 49104 43020 49138
rect 43192 49104 43204 49138
rect 43008 49098 43204 49104
rect 43702 49138 43898 49144
rect 43702 49104 43714 49138
rect 43886 49104 43898 49138
rect 43702 49098 43898 49104
rect 44396 49138 44592 49144
rect 44396 49104 44408 49138
rect 44580 49104 44592 49138
rect 44396 49098 44592 49104
rect 45090 49138 45286 49144
rect 45090 49104 45102 49138
rect 45274 49104 45286 49138
rect 45090 49098 45286 49104
rect 46308 49138 46504 49144
rect 46308 49104 46320 49138
rect 46492 49104 46504 49138
rect 46308 49098 46504 49104
rect 47002 49138 47198 49144
rect 47002 49104 47014 49138
rect 47186 49104 47198 49138
rect 47002 49098 47198 49104
rect 47696 49138 47892 49144
rect 47696 49104 47708 49138
rect 47880 49104 47892 49138
rect 47696 49098 47892 49104
rect 48390 49138 48586 49144
rect 48390 49104 48402 49138
rect 48574 49104 48586 49138
rect 48390 49098 48586 49104
rect 49084 49138 49280 49144
rect 49084 49104 49096 49138
rect 49268 49104 49280 49138
rect 49084 49098 49280 49104
rect 50330 49138 50526 49144
rect 50330 49104 50342 49138
rect 50514 49104 50526 49138
rect 50330 49098 50526 49104
rect 51024 49138 51220 49144
rect 51024 49104 51036 49138
rect 51208 49104 51220 49138
rect 51024 49098 51220 49104
rect 51718 49138 51914 49144
rect 51718 49104 51730 49138
rect 51902 49104 51914 49138
rect 51718 49098 51914 49104
rect 52412 49138 52608 49144
rect 52412 49104 52424 49138
rect 52596 49104 52608 49138
rect 52412 49098 52608 49104
rect 53106 49138 53302 49144
rect 53106 49104 53118 49138
rect 53290 49104 53302 49138
rect 53106 49098 53302 49104
rect 54352 49138 54548 49144
rect 54352 49104 54364 49138
rect 54536 49104 54548 49138
rect 54352 49098 54548 49104
rect 55046 49138 55242 49144
rect 55046 49104 55058 49138
rect 55230 49104 55242 49138
rect 55046 49098 55242 49104
rect 55740 49138 55936 49144
rect 55740 49104 55752 49138
rect 55924 49104 55936 49138
rect 55740 49098 55936 49104
rect 56434 49138 56630 49144
rect 56434 49104 56446 49138
rect 56618 49104 56630 49138
rect 56434 49098 56630 49104
rect 57128 49138 57324 49144
rect 57128 49104 57140 49138
rect 57312 49104 57324 49138
rect 57128 49098 57324 49104
rect 38414 47838 38424 48764
rect 39756 47838 39766 48764
rect 42314 48480 42510 48486
rect 42314 48446 42326 48480
rect 42498 48446 42510 48480
rect 42314 48440 42510 48446
rect 43008 48480 43204 48486
rect 43008 48446 43020 48480
rect 43192 48446 43204 48480
rect 43008 48440 43204 48446
rect 43702 48480 43898 48486
rect 43702 48446 43714 48480
rect 43886 48446 43898 48480
rect 43702 48440 43898 48446
rect 44396 48480 44592 48486
rect 44396 48446 44408 48480
rect 44580 48446 44592 48480
rect 44396 48440 44592 48446
rect 45090 48480 45286 48486
rect 45090 48446 45102 48480
rect 45274 48446 45286 48480
rect 45090 48440 45286 48446
rect 46308 48480 46504 48486
rect 46308 48446 46320 48480
rect 46492 48446 46504 48480
rect 46308 48440 46504 48446
rect 47002 48480 47198 48486
rect 47002 48446 47014 48480
rect 47186 48446 47198 48480
rect 47002 48440 47198 48446
rect 47696 48480 47892 48486
rect 47696 48446 47708 48480
rect 47880 48446 47892 48480
rect 47696 48440 47892 48446
rect 48390 48480 48586 48486
rect 48390 48446 48402 48480
rect 48574 48446 48586 48480
rect 48390 48440 48586 48446
rect 49084 48480 49280 48486
rect 49084 48446 49096 48480
rect 49268 48446 49280 48480
rect 49084 48440 49280 48446
rect 50330 48480 50526 48486
rect 50330 48446 50342 48480
rect 50514 48446 50526 48480
rect 50330 48440 50526 48446
rect 51024 48480 51220 48486
rect 51024 48446 51036 48480
rect 51208 48446 51220 48480
rect 51024 48440 51220 48446
rect 51718 48480 51914 48486
rect 51718 48446 51730 48480
rect 51902 48446 51914 48480
rect 51718 48440 51914 48446
rect 52412 48480 52608 48486
rect 52412 48446 52424 48480
rect 52596 48446 52608 48480
rect 52412 48440 52608 48446
rect 53106 48480 53302 48486
rect 53106 48446 53118 48480
rect 53290 48446 53302 48480
rect 53106 48440 53302 48446
rect 54352 48480 54548 48486
rect 54352 48446 54364 48480
rect 54536 48446 54548 48480
rect 54352 48440 54548 48446
rect 55046 48480 55242 48486
rect 55046 48446 55058 48480
rect 55230 48446 55242 48480
rect 55046 48440 55242 48446
rect 55740 48480 55936 48486
rect 55740 48446 55752 48480
rect 55924 48446 55936 48480
rect 55740 48440 55936 48446
rect 56434 48480 56630 48486
rect 56434 48446 56446 48480
rect 56618 48446 56630 48480
rect 56434 48440 56630 48446
rect 57128 48480 57324 48486
rect 57128 48446 57140 48480
rect 57312 48446 57324 48480
rect 57128 48440 57324 48446
rect 42620 48112 44984 48258
rect 42620 47994 42872 48112
rect 44786 47994 44984 48112
rect 21354 46256 21640 46432
rect 11016 43708 11290 43774
rect 11016 43646 11074 43708
rect 11216 43646 11290 43708
rect 11016 43566 11290 43646
rect 1952 43052 1998 43064
rect 1952 42760 1958 43052
rect 1992 42760 1998 43052
rect 1952 42748 1998 42760
rect 3010 43052 3056 43064
rect 3010 42760 3016 43052
rect 3050 42760 3056 43052
rect 3010 42748 3056 42760
rect 4068 43052 4114 43064
rect 4068 42760 4074 43052
rect 4108 42760 4114 43052
rect 4068 42748 4114 42760
rect 5126 43052 5172 43064
rect 5126 42760 5132 43052
rect 5166 42760 5172 43052
rect 5126 42748 5172 42760
rect 6184 43052 6230 43064
rect 6184 42760 6190 43052
rect 6224 42760 6230 43052
rect 6184 42748 6230 42760
rect 7242 43052 7288 43064
rect 7242 42760 7248 43052
rect 7282 42760 7288 43052
rect 7242 42748 7288 42760
rect 8466 43060 8512 43072
rect 8466 42768 8472 43060
rect 8506 42768 8512 43060
rect 8466 42756 8512 42768
rect 9524 43060 9570 43072
rect 9524 42768 9530 43060
rect 9564 42768 9570 43060
rect 9524 42756 9570 42768
rect 10582 43060 10628 43072
rect 10582 42768 10588 43060
rect 10622 42768 10628 43060
rect 10582 42756 10628 42768
rect 11640 43060 11686 43072
rect 11640 42768 11646 43060
rect 11680 42768 11686 43060
rect 11640 42756 11686 42768
rect 12698 43060 12744 43072
rect 12698 42768 12704 43060
rect 12738 42768 12744 43060
rect 12698 42756 12744 42768
rect 13756 43060 13802 43072
rect 13756 42768 13762 43060
rect 13796 42768 13802 43060
rect 13756 42756 13802 42768
rect 14972 43068 15018 43080
rect 14972 42776 14978 43068
rect 15012 42776 15018 43068
rect 14972 42764 15018 42776
rect 16030 43068 16076 43080
rect 16030 42776 16036 43068
rect 16070 42776 16076 43068
rect 16030 42764 16076 42776
rect 17088 43068 17134 43080
rect 17088 42776 17094 43068
rect 17128 42776 17134 43068
rect 17088 42764 17134 42776
rect 18146 43068 18192 43080
rect 18146 42776 18152 43068
rect 18186 42776 18192 43068
rect 18146 42764 18192 42776
rect 19204 43068 19250 43080
rect 19204 42776 19210 43068
rect 19244 42776 19250 43068
rect 19204 42764 19250 42776
rect 20262 43068 20308 43080
rect 20262 42776 20268 43068
rect 20302 42776 20308 43068
rect 21384 43052 21640 46256
rect 39090 45178 39496 47838
rect 42620 47836 44984 47994
rect 46528 48126 49418 48218
rect 46528 47968 46870 48126
rect 49234 47968 49418 48126
rect 46528 47862 49418 47968
rect 50606 48086 53444 48206
rect 50606 47954 50844 48086
rect 53232 47954 53444 48086
rect 50606 47848 53444 47954
rect 54354 48140 57272 48218
rect 54354 47954 54540 48140
rect 57088 47954 57272 48140
rect 54354 47862 57272 47954
rect 66814 46560 66824 46688
rect 66550 46530 66824 46560
rect 66172 46524 66824 46530
rect 66172 46248 66184 46524
rect 66696 46248 66824 46524
rect 66172 46242 66824 46248
rect 66550 46158 66824 46242
rect 66814 45974 66824 46158
rect 67244 45974 67254 46688
rect 24024 44984 25442 45070
rect 24024 44696 24382 44984
rect 25184 44696 25442 44984
rect 24024 44582 25442 44696
rect 38714 45004 42794 45178
rect 38714 44424 39408 45004
rect 41694 44424 42794 45004
rect 38714 44308 42794 44424
rect 49454 43888 50070 44004
rect 49454 43720 49622 43888
rect 49866 43720 50070 43888
rect 49454 43614 50070 43720
rect 63792 43614 64238 43652
rect 67818 43628 68038 49850
rect 75722 48690 76408 48696
rect 75722 48226 75734 48690
rect 76396 48226 76408 48690
rect 75722 48220 76408 48226
rect 68188 47424 68198 47812
rect 68884 47424 68894 47812
rect 75960 47790 76198 48220
rect 77294 48002 77620 50798
rect 68408 43984 68610 47424
rect 75714 47308 75724 47790
rect 76368 47308 76378 47790
rect 73050 46020 73060 46882
rect 73674 46672 73684 46882
rect 77264 46672 77620 48002
rect 73674 46636 77620 46672
rect 80598 46636 80954 46672
rect 73674 46204 80954 46636
rect 73674 46020 73684 46204
rect 68276 43922 69060 43984
rect 68276 43844 68426 43922
rect 68848 43844 69060 43922
rect 68276 43782 69060 43844
rect 63792 43492 63846 43614
rect 64132 43492 64238 43614
rect 63792 43444 64238 43492
rect 67732 43614 68038 43628
rect 67732 43584 68228 43614
rect 67732 43482 67844 43584
rect 68066 43482 68228 43584
rect 67732 43396 68228 43482
rect 71570 43584 71878 43638
rect 71570 43472 71644 43584
rect 71790 43472 71878 43584
rect 71570 43426 71878 43472
rect 70104 43124 70150 43136
rect 54086 43110 54132 43122
rect 47572 43096 47618 43108
rect 27984 43068 28030 43080
rect 21384 42946 21468 43052
rect 20262 42764 20308 42776
rect 21462 42760 21468 42946
rect 21502 42946 21640 43052
rect 22520 43052 22566 43064
rect 21502 42760 21508 42946
rect 21462 42748 21508 42760
rect 22520 42760 22526 43052
rect 22560 42760 22566 43052
rect 22520 42748 22566 42760
rect 23578 43052 23624 43064
rect 23578 42760 23584 43052
rect 23618 42760 23624 43052
rect 23578 42748 23624 42760
rect 24636 43052 24682 43064
rect 24636 42760 24642 43052
rect 24676 42760 24682 43052
rect 24636 42748 24682 42760
rect 25694 43052 25740 43064
rect 25694 42760 25700 43052
rect 25734 42760 25740 43052
rect 25694 42748 25740 42760
rect 26752 43052 26798 43064
rect 26752 42760 26758 43052
rect 26792 42760 26798 43052
rect 27984 42776 27990 43068
rect 28024 42776 28030 43068
rect 27984 42764 28030 42776
rect 29042 43068 29088 43080
rect 29042 42776 29048 43068
rect 29082 42776 29088 43068
rect 29042 42764 29088 42776
rect 30100 43068 30146 43080
rect 30100 42776 30106 43068
rect 30140 42776 30146 43068
rect 30100 42764 30146 42776
rect 31158 43068 31204 43080
rect 31158 42776 31164 43068
rect 31198 42776 31204 43068
rect 31158 42764 31204 42776
rect 32216 43068 32262 43080
rect 32216 42776 32222 43068
rect 32256 42776 32262 43068
rect 32216 42764 32262 42776
rect 33274 43068 33320 43080
rect 33274 42776 33280 43068
rect 33314 42776 33320 43068
rect 33274 42764 33320 42776
rect 34494 43074 34540 43086
rect 34494 42782 34500 43074
rect 34534 42782 34540 43074
rect 34494 42770 34540 42782
rect 35552 43074 35598 43086
rect 35552 42782 35558 43074
rect 35592 42782 35598 43074
rect 35552 42770 35598 42782
rect 36610 43074 36656 43086
rect 36610 42782 36616 43074
rect 36650 42782 36656 43074
rect 36610 42770 36656 42782
rect 37668 43074 37714 43086
rect 37668 42782 37674 43074
rect 37708 42782 37714 43074
rect 37668 42770 37714 42782
rect 38726 43074 38772 43086
rect 38726 42782 38732 43074
rect 38766 42782 38772 43074
rect 38726 42770 38772 42782
rect 39784 43074 39830 43086
rect 39784 42782 39790 43074
rect 39824 42782 39830 43074
rect 39784 42770 39830 42782
rect 40984 43074 41030 43086
rect 40984 42782 40990 43074
rect 41024 42782 41030 43074
rect 40984 42770 41030 42782
rect 42042 43074 42088 43086
rect 42042 42782 42048 43074
rect 42082 42782 42088 43074
rect 42042 42770 42088 42782
rect 43100 43074 43146 43086
rect 43100 42782 43106 43074
rect 43140 42782 43146 43074
rect 43100 42770 43146 42782
rect 44158 43074 44204 43086
rect 44158 42782 44164 43074
rect 44198 42782 44204 43074
rect 44158 42770 44204 42782
rect 45216 43074 45262 43086
rect 45216 42782 45222 43074
rect 45256 42782 45262 43074
rect 45216 42770 45262 42782
rect 46274 43074 46320 43086
rect 46274 42782 46280 43074
rect 46314 42782 46320 43074
rect 47572 42804 47578 43096
rect 47612 42804 47618 43096
rect 47572 42792 47618 42804
rect 48630 43096 48676 43108
rect 48630 42804 48636 43096
rect 48670 42804 48676 43096
rect 48630 42792 48676 42804
rect 49688 43096 49734 43108
rect 49688 42804 49694 43096
rect 49728 42804 49734 43096
rect 49688 42792 49734 42804
rect 50746 43096 50792 43108
rect 50746 42804 50752 43096
rect 50786 42804 50792 43096
rect 50746 42792 50792 42804
rect 51804 43096 51850 43108
rect 51804 42804 51810 43096
rect 51844 42804 51850 43096
rect 51804 42792 51850 42804
rect 52862 43096 52908 43108
rect 52862 42804 52868 43096
rect 52902 42804 52908 43096
rect 54086 42818 54092 43110
rect 54126 42818 54132 43110
rect 54086 42806 54132 42818
rect 55144 43110 55190 43122
rect 55144 42818 55150 43110
rect 55184 42818 55190 43110
rect 55144 42806 55190 42818
rect 56202 43110 56248 43122
rect 56202 42818 56208 43110
rect 56242 42818 56248 43110
rect 56202 42806 56248 42818
rect 57260 43110 57306 43122
rect 57260 42818 57266 43110
rect 57300 42818 57306 43110
rect 57260 42806 57306 42818
rect 58318 43110 58364 43122
rect 58318 42818 58324 43110
rect 58358 42818 58364 43110
rect 58318 42806 58364 42818
rect 59376 43110 59422 43122
rect 59376 42818 59382 43110
rect 59416 42818 59422 43110
rect 62502 43108 62548 43120
rect 62502 42936 62508 43108
rect 62542 42936 62548 43108
rect 62502 42924 62548 42936
rect 63160 43108 63206 43120
rect 63160 42936 63166 43108
rect 63200 42936 63206 43108
rect 63160 42924 63206 42936
rect 63818 43108 63864 43120
rect 63818 42936 63824 43108
rect 63858 42936 63864 43108
rect 63818 42924 63864 42936
rect 64476 43108 64522 43120
rect 64476 42936 64482 43108
rect 64516 42936 64522 43108
rect 64476 42924 64522 42936
rect 65134 43108 65180 43120
rect 65134 42936 65140 43108
rect 65174 42936 65180 43108
rect 65134 42924 65180 42936
rect 65792 43108 65838 43120
rect 65792 42936 65798 43108
rect 65832 42936 65838 43108
rect 65792 42924 65838 42936
rect 66296 43110 66342 43122
rect 66296 42938 66302 43110
rect 66336 42938 66342 43110
rect 66296 42926 66342 42938
rect 66954 43110 67000 43122
rect 66954 42938 66960 43110
rect 66994 42938 67000 43110
rect 66954 42926 67000 42938
rect 67612 43110 67658 43122
rect 67612 42938 67618 43110
rect 67652 42938 67658 43110
rect 67612 42926 67658 42938
rect 68270 43110 68316 43122
rect 68270 42938 68276 43110
rect 68310 42938 68316 43110
rect 68270 42926 68316 42938
rect 68928 43110 68974 43122
rect 68928 42938 68934 43110
rect 68968 42938 68974 43110
rect 68928 42926 68974 42938
rect 69586 43110 69632 43122
rect 69586 42938 69592 43110
rect 69626 42938 69632 43110
rect 70104 42952 70110 43124
rect 70144 42952 70150 43124
rect 70104 42940 70150 42952
rect 70762 43124 70808 43136
rect 70762 42952 70768 43124
rect 70802 42952 70808 43124
rect 70762 42940 70808 42952
rect 71420 43124 71466 43136
rect 71420 42952 71426 43124
rect 71460 42952 71466 43124
rect 71420 42940 71466 42952
rect 72078 43124 72124 43136
rect 72078 42952 72084 43124
rect 72118 42952 72124 43124
rect 72078 42940 72124 42952
rect 72736 43124 72782 43136
rect 72736 42952 72742 43124
rect 72776 42952 72782 43124
rect 72736 42940 72782 42952
rect 73394 43124 73440 43136
rect 73394 42952 73400 43124
rect 73434 42952 73440 43124
rect 79160 43104 79170 43578
rect 79870 43104 79880 43578
rect 79424 43100 79728 43104
rect 79424 43084 79608 43100
rect 73394 42940 73440 42952
rect 69586 42926 69632 42938
rect 59376 42806 59422 42818
rect 73610 42876 73950 43002
rect 52862 42792 52908 42804
rect 46274 42770 46320 42782
rect 26752 42748 26798 42760
rect 62148 42532 62360 42700
rect 54086 42016 54132 42028
rect 47572 42002 47618 42014
rect 1952 41958 1998 41970
rect 1952 41666 1958 41958
rect 1992 41666 1998 41958
rect 1952 41654 1998 41666
rect 3010 41958 3056 41970
rect 3010 41666 3016 41958
rect 3050 41666 3056 41958
rect 3010 41654 3056 41666
rect 4068 41958 4114 41970
rect 4068 41666 4074 41958
rect 4108 41666 4114 41958
rect 4068 41654 4114 41666
rect 5126 41958 5172 41970
rect 5126 41666 5132 41958
rect 5166 41666 5172 41958
rect 5126 41654 5172 41666
rect 6184 41958 6230 41970
rect 6184 41666 6190 41958
rect 6224 41666 6230 41958
rect 6184 41654 6230 41666
rect 7242 41958 7288 41970
rect 7242 41666 7248 41958
rect 7282 41666 7288 41958
rect 8466 41966 8512 41978
rect 7242 41654 7288 41666
rect 1304 41518 1454 41644
rect 1304 41416 1326 41518
rect 1264 40322 1326 41416
rect 1420 41416 1454 41518
rect 7722 41526 8018 41824
rect 8466 41674 8472 41966
rect 8506 41674 8512 41966
rect 8466 41662 8512 41674
rect 9524 41966 9570 41978
rect 9524 41674 9530 41966
rect 9564 41674 9570 41966
rect 9524 41662 9570 41674
rect 10582 41966 10628 41978
rect 10582 41674 10588 41966
rect 10622 41674 10628 41966
rect 10582 41662 10628 41674
rect 11640 41966 11686 41978
rect 11640 41674 11646 41966
rect 11680 41674 11686 41966
rect 11640 41662 11686 41674
rect 12698 41966 12744 41978
rect 12698 41674 12704 41966
rect 12738 41674 12744 41966
rect 12698 41662 12744 41674
rect 13756 41966 13802 41978
rect 13756 41674 13762 41966
rect 13796 41674 13802 41966
rect 13756 41662 13802 41674
rect 14972 41974 15018 41986
rect 14972 41682 14978 41974
rect 15012 41682 15018 41974
rect 14972 41670 15018 41682
rect 16030 41974 16076 41986
rect 16030 41682 16036 41974
rect 16070 41682 16076 41974
rect 16030 41670 16076 41682
rect 17088 41974 17134 41986
rect 17088 41682 17094 41974
rect 17128 41682 17134 41974
rect 17088 41670 17134 41682
rect 18146 41974 18192 41986
rect 18146 41682 18152 41974
rect 18186 41682 18192 41974
rect 18146 41670 18192 41682
rect 19204 41974 19250 41986
rect 19204 41682 19210 41974
rect 19244 41682 19250 41974
rect 19204 41670 19250 41682
rect 20262 41974 20308 41986
rect 20262 41682 20268 41974
rect 20302 41682 20308 41974
rect 27984 41974 28030 41986
rect 21462 41958 21508 41970
rect 20262 41670 20308 41682
rect 14324 41602 14474 41660
rect 1420 40322 1560 41416
rect 1952 40864 1998 40876
rect 1952 40572 1958 40864
rect 1992 40572 1998 40864
rect 1952 40560 1998 40572
rect 3010 40864 3056 40876
rect 3010 40572 3016 40864
rect 3050 40572 3056 40864
rect 3010 40560 3056 40572
rect 4068 40864 4114 40876
rect 4068 40572 4074 40864
rect 4108 40572 4114 40864
rect 4068 40560 4114 40572
rect 5126 40864 5172 40876
rect 5126 40572 5132 40864
rect 5166 40572 5172 40864
rect 5126 40560 5172 40572
rect 6184 40864 6230 40876
rect 6184 40572 6190 40864
rect 6224 40572 6230 40864
rect 6184 40560 6230 40572
rect 7242 40864 7288 40876
rect 7242 40572 7248 40864
rect 7282 40572 7288 40864
rect 7242 40560 7288 40572
rect 1264 35702 1560 40322
rect 7722 40330 7840 41526
rect 7934 40838 8018 41526
rect 14216 41534 14512 41602
rect 8466 40872 8512 40884
rect 8466 40838 8472 40872
rect 7934 40580 8472 40838
rect 8506 40580 8512 40872
rect 7934 40568 8512 40580
rect 9524 40872 9570 40884
rect 9524 40580 9530 40872
rect 9564 40580 9570 40872
rect 9524 40568 9570 40580
rect 10582 40872 10628 40884
rect 10582 40580 10588 40872
rect 10622 40580 10628 40872
rect 10582 40568 10628 40580
rect 11640 40872 11686 40884
rect 11640 40580 11646 40872
rect 11680 40580 11686 40872
rect 11640 40568 11686 40580
rect 12698 40872 12744 40884
rect 12698 40580 12704 40872
rect 12738 40580 12744 40872
rect 12698 40568 12744 40580
rect 13756 40876 13802 40884
rect 14216 40876 14346 41534
rect 13756 40872 14346 40876
rect 13756 40580 13762 40872
rect 13796 40580 14346 40872
rect 13756 40574 14346 40580
rect 13756 40568 13802 40574
rect 7934 40536 8496 40568
rect 7934 40330 8018 40536
rect 1952 39770 1998 39782
rect 1952 39478 1958 39770
rect 1992 39478 1998 39770
rect 1952 39466 1998 39478
rect 3010 39770 3056 39782
rect 3010 39478 3016 39770
rect 3050 39478 3056 39770
rect 3010 39466 3056 39478
rect 4068 39770 4114 39782
rect 4068 39478 4074 39770
rect 4108 39478 4114 39770
rect 4068 39466 4114 39478
rect 5126 39770 5172 39782
rect 5126 39478 5132 39770
rect 5166 39478 5172 39770
rect 5126 39466 5172 39478
rect 6184 39770 6230 39782
rect 6184 39478 6190 39770
rect 6224 39478 6230 39770
rect 6184 39466 6230 39478
rect 7242 39770 7288 39782
rect 7242 39478 7248 39770
rect 7282 39478 7288 39770
rect 7242 39466 7288 39478
rect 1952 38676 1998 38688
rect 1952 38384 1958 38676
rect 1992 38384 1998 38676
rect 1952 38372 1998 38384
rect 3010 38676 3056 38688
rect 3010 38384 3016 38676
rect 3050 38384 3056 38676
rect 3010 38372 3056 38384
rect 4068 38676 4114 38688
rect 4068 38384 4074 38676
rect 4108 38384 4114 38676
rect 4068 38372 4114 38384
rect 5126 38676 5172 38688
rect 5126 38384 5132 38676
rect 5166 38384 5172 38676
rect 5126 38372 5172 38384
rect 6184 38676 6230 38688
rect 6184 38384 6190 38676
rect 6224 38384 6230 38676
rect 6184 38372 6230 38384
rect 7242 38676 7288 38688
rect 7242 38384 7248 38676
rect 7282 38384 7288 38676
rect 7242 38372 7288 38384
rect 1952 37236 1998 37248
rect 1952 36944 1958 37236
rect 1992 36944 1998 37236
rect 1952 36932 1998 36944
rect 3010 37236 3056 37248
rect 3010 36944 3016 37236
rect 3050 36944 3056 37236
rect 3010 36932 3056 36944
rect 4068 37236 4114 37248
rect 4068 36944 4074 37236
rect 4108 36944 4114 37236
rect 4068 36932 4114 36944
rect 5126 37236 5172 37248
rect 5126 36944 5132 37236
rect 5166 36944 5172 37236
rect 5126 36932 5172 36944
rect 6184 37236 6230 37248
rect 6184 36944 6190 37236
rect 6224 36944 6230 37236
rect 6184 36932 6230 36944
rect 7242 37236 7288 37248
rect 7242 36944 7248 37236
rect 7282 36944 7288 37236
rect 7242 36932 7288 36944
rect 1952 36142 1998 36154
rect 1952 35850 1958 36142
rect 1992 35850 1998 36142
rect 1952 35838 1998 35850
rect 3010 36142 3056 36154
rect 3010 35850 3016 36142
rect 3050 35850 3056 36142
rect 3010 35838 3056 35850
rect 4068 36142 4114 36154
rect 4068 35850 4074 36142
rect 4108 35850 4114 36142
rect 4068 35838 4114 35850
rect 5126 36142 5172 36154
rect 5126 35850 5132 36142
rect 5166 35850 5172 36142
rect 5126 35838 5172 35850
rect 6184 36142 6230 36154
rect 6184 35850 6190 36142
rect 6224 35850 6230 36142
rect 6184 35838 6230 35850
rect 7242 36142 7288 36154
rect 7242 35850 7248 36142
rect 7282 35850 7288 36142
rect 7242 35838 7288 35850
rect 1264 34506 1326 35702
rect 1420 34506 1560 35702
rect 7722 35710 8018 40330
rect 14216 40338 14346 40574
rect 14440 40338 14512 41534
rect 20748 41518 21044 41712
rect 21462 41666 21468 41958
rect 21502 41666 21508 41958
rect 21462 41654 21508 41666
rect 22520 41958 22566 41970
rect 22520 41666 22526 41958
rect 22560 41666 22566 41958
rect 22520 41654 22566 41666
rect 23578 41958 23624 41970
rect 23578 41666 23584 41958
rect 23618 41666 23624 41958
rect 23578 41654 23624 41666
rect 24636 41958 24682 41970
rect 24636 41666 24642 41958
rect 24676 41666 24682 41958
rect 24636 41654 24682 41666
rect 25694 41958 25740 41970
rect 25694 41666 25700 41958
rect 25734 41666 25740 41958
rect 25694 41654 25740 41666
rect 26752 41958 26798 41970
rect 26752 41666 26758 41958
rect 26792 41666 26798 41958
rect 27984 41682 27990 41974
rect 28024 41682 28030 41974
rect 27984 41670 28030 41682
rect 29042 41974 29088 41986
rect 29042 41682 29048 41974
rect 29082 41682 29088 41974
rect 29042 41670 29088 41682
rect 30100 41974 30146 41986
rect 30100 41682 30106 41974
rect 30140 41682 30146 41974
rect 30100 41670 30146 41682
rect 31158 41974 31204 41986
rect 31158 41682 31164 41974
rect 31198 41682 31204 41974
rect 31158 41670 31204 41682
rect 32216 41974 32262 41986
rect 32216 41682 32222 41974
rect 32256 41682 32262 41974
rect 32216 41670 32262 41682
rect 33274 41974 33320 41986
rect 33274 41682 33280 41974
rect 33314 41682 33320 41974
rect 33274 41670 33320 41682
rect 34494 41980 34540 41992
rect 34494 41688 34500 41980
rect 34534 41688 34540 41980
rect 34494 41676 34540 41688
rect 35552 41980 35598 41992
rect 35552 41688 35558 41980
rect 35592 41688 35598 41980
rect 35552 41676 35598 41688
rect 36610 41980 36656 41992
rect 36610 41688 36616 41980
rect 36650 41688 36656 41980
rect 36610 41676 36656 41688
rect 37668 41980 37714 41992
rect 37668 41688 37674 41980
rect 37708 41688 37714 41980
rect 37668 41676 37714 41688
rect 38726 41980 38772 41992
rect 38726 41688 38732 41980
rect 38766 41688 38772 41980
rect 38726 41676 38772 41688
rect 39784 41980 39830 41992
rect 39784 41688 39790 41980
rect 39824 41688 39830 41980
rect 39784 41676 39830 41688
rect 40984 41980 41030 41992
rect 40984 41688 40990 41980
rect 41024 41688 41030 41980
rect 40984 41676 41030 41688
rect 42042 41980 42088 41992
rect 42042 41688 42048 41980
rect 42082 41688 42088 41980
rect 42042 41676 42088 41688
rect 43100 41980 43146 41992
rect 43100 41688 43106 41980
rect 43140 41688 43146 41980
rect 43100 41676 43146 41688
rect 44158 41980 44204 41992
rect 44158 41688 44164 41980
rect 44198 41688 44204 41980
rect 44158 41676 44204 41688
rect 45216 41980 45262 41992
rect 45216 41688 45222 41980
rect 45256 41688 45262 41980
rect 45216 41676 45262 41688
rect 46274 41980 46320 41992
rect 46274 41688 46280 41980
rect 46314 41688 46320 41980
rect 47572 41710 47578 42002
rect 47612 41710 47618 42002
rect 47572 41698 47618 41710
rect 48630 42002 48676 42014
rect 48630 41710 48636 42002
rect 48670 41710 48676 42002
rect 48630 41698 48676 41710
rect 49688 42002 49734 42014
rect 49688 41710 49694 42002
rect 49728 41710 49734 42002
rect 49688 41698 49734 41710
rect 50746 42002 50792 42014
rect 50746 41710 50752 42002
rect 50786 41710 50792 42002
rect 50746 41698 50792 41710
rect 51804 42002 51850 42014
rect 51804 41710 51810 42002
rect 51844 41710 51850 42002
rect 51804 41698 51850 41710
rect 52862 42002 52908 42014
rect 52862 41710 52868 42002
rect 52902 41710 52908 42002
rect 54086 41724 54092 42016
rect 54126 41724 54132 42016
rect 54086 41712 54132 41724
rect 55144 42016 55190 42028
rect 55144 41724 55150 42016
rect 55184 41724 55190 42016
rect 55144 41712 55190 41724
rect 56202 42016 56248 42028
rect 56202 41724 56208 42016
rect 56242 41724 56248 42016
rect 56202 41712 56248 41724
rect 57260 42016 57306 42028
rect 57260 41724 57266 42016
rect 57300 41724 57306 42016
rect 57260 41712 57306 41724
rect 58318 42016 58364 42028
rect 58318 41724 58324 42016
rect 58358 41724 58364 42016
rect 58318 41712 58364 41724
rect 59376 42016 59422 42028
rect 59376 41724 59382 42016
rect 59416 41724 59422 42016
rect 59376 41712 59422 41724
rect 59530 41772 59934 41952
rect 52862 41698 52908 41710
rect 46274 41676 46320 41688
rect 26752 41654 26798 41666
rect 14972 40880 15018 40892
rect 14972 40588 14978 40880
rect 15012 40588 15018 40880
rect 14972 40576 15018 40588
rect 16030 40880 16076 40892
rect 16030 40588 16036 40880
rect 16070 40588 16076 40880
rect 16030 40576 16076 40588
rect 17088 40880 17134 40892
rect 17088 40588 17094 40880
rect 17128 40588 17134 40880
rect 17088 40576 17134 40588
rect 18146 40880 18192 40892
rect 18146 40588 18152 40880
rect 18186 40588 18192 40880
rect 18146 40576 18192 40588
rect 19204 40880 19250 40892
rect 19204 40588 19210 40880
rect 19244 40588 19250 40880
rect 19204 40576 19250 40588
rect 20262 40880 20308 40892
rect 20262 40588 20268 40880
rect 20302 40588 20308 40880
rect 20748 40840 20836 41518
rect 20262 40576 20308 40588
rect 20338 40538 20836 40840
rect 8466 39778 8512 39790
rect 8466 39486 8472 39778
rect 8506 39486 8512 39778
rect 8466 39474 8512 39486
rect 9524 39778 9570 39790
rect 9524 39486 9530 39778
rect 9564 39486 9570 39778
rect 9524 39474 9570 39486
rect 10582 39778 10628 39790
rect 10582 39486 10588 39778
rect 10622 39486 10628 39778
rect 10582 39474 10628 39486
rect 11640 39778 11686 39790
rect 11640 39486 11646 39778
rect 11680 39486 11686 39778
rect 11640 39474 11686 39486
rect 12698 39778 12744 39790
rect 12698 39486 12704 39778
rect 12738 39486 12744 39778
rect 12698 39474 12744 39486
rect 13756 39778 13802 39790
rect 13756 39486 13762 39778
rect 13796 39486 13802 39778
rect 13756 39474 13802 39486
rect 8466 38684 8512 38696
rect 8466 38392 8472 38684
rect 8506 38392 8512 38684
rect 8466 38380 8512 38392
rect 9524 38684 9570 38696
rect 9524 38392 9530 38684
rect 9564 38392 9570 38684
rect 9524 38380 9570 38392
rect 10582 38684 10628 38696
rect 10582 38392 10588 38684
rect 10622 38392 10628 38684
rect 10582 38380 10628 38392
rect 11640 38684 11686 38696
rect 11640 38392 11646 38684
rect 11680 38392 11686 38684
rect 11640 38380 11686 38392
rect 12698 38684 12744 38696
rect 12698 38392 12704 38684
rect 12738 38392 12744 38684
rect 12698 38380 12744 38392
rect 13756 38684 13802 38696
rect 13756 38392 13762 38684
rect 13796 38392 13802 38684
rect 13756 38380 13802 38392
rect 8466 37244 8512 37256
rect 8466 36952 8472 37244
rect 8506 36952 8512 37244
rect 8466 36940 8512 36952
rect 9524 37244 9570 37256
rect 9524 36952 9530 37244
rect 9564 36952 9570 37244
rect 9524 36940 9570 36952
rect 10582 37244 10628 37256
rect 10582 36952 10588 37244
rect 10622 36952 10628 37244
rect 10582 36940 10628 36952
rect 11640 37244 11686 37256
rect 11640 36952 11646 37244
rect 11680 36952 11686 37244
rect 11640 36940 11686 36952
rect 12698 37244 12744 37256
rect 12698 36952 12704 37244
rect 12738 36952 12744 37244
rect 12698 36940 12744 36952
rect 13756 37244 13802 37256
rect 13756 36952 13762 37244
rect 13796 36952 13802 37244
rect 13756 36940 13802 36952
rect 8466 36150 8512 36162
rect 8466 35858 8472 36150
rect 8506 35858 8512 36150
rect 8466 35846 8512 35858
rect 9524 36150 9570 36162
rect 9524 35858 9530 36150
rect 9564 35858 9570 36150
rect 9524 35846 9570 35858
rect 10582 36150 10628 36162
rect 10582 35858 10588 36150
rect 10622 35858 10628 36150
rect 10582 35846 10628 35858
rect 11640 36150 11686 36162
rect 11640 35858 11646 36150
rect 11680 35858 11686 36150
rect 11640 35846 11686 35858
rect 12698 36150 12744 36162
rect 12698 35858 12704 36150
rect 12738 35858 12744 36150
rect 12698 35846 12744 35858
rect 13756 36150 13802 36162
rect 13756 35858 13762 36150
rect 13796 35858 13802 36150
rect 13756 35846 13802 35858
rect 1952 35048 1998 35060
rect 1952 34756 1958 35048
rect 1992 34756 1998 35048
rect 1952 34744 1998 34756
rect 3010 35048 3056 35060
rect 3010 34756 3016 35048
rect 3050 34756 3056 35048
rect 3010 34744 3056 34756
rect 4068 35048 4114 35060
rect 4068 34756 4074 35048
rect 4108 34756 4114 35048
rect 4068 34744 4114 34756
rect 5126 35048 5172 35060
rect 5126 34756 5132 35048
rect 5166 34756 5172 35048
rect 5126 34744 5172 34756
rect 6184 35048 6230 35060
rect 6184 34756 6190 35048
rect 6224 34756 6230 35048
rect 6184 34744 6230 34756
rect 7242 35048 7288 35060
rect 7242 34756 7248 35048
rect 7282 34756 7288 35048
rect 7242 34744 7288 34756
rect 1264 29868 1560 34506
rect 7722 34514 7840 35710
rect 7934 34514 8018 35710
rect 14216 35718 14512 40338
rect 20748 40322 20836 40538
rect 20930 40322 21044 41518
rect 27336 41534 27486 41660
rect 27336 40970 27358 41534
rect 21462 40864 21508 40876
rect 21462 40572 21468 40864
rect 21502 40572 21508 40864
rect 21462 40560 21508 40572
rect 22520 40864 22566 40876
rect 22520 40572 22526 40864
rect 22560 40572 22566 40864
rect 22520 40560 22566 40572
rect 23578 40864 23624 40876
rect 23578 40572 23584 40864
rect 23618 40572 23624 40864
rect 23578 40560 23624 40572
rect 24636 40864 24682 40876
rect 24636 40572 24642 40864
rect 24676 40572 24682 40864
rect 24636 40560 24682 40572
rect 25694 40864 25740 40876
rect 25694 40572 25700 40864
rect 25734 40572 25740 40864
rect 25694 40560 25740 40572
rect 26752 40864 26798 40876
rect 26752 40572 26758 40864
rect 26792 40572 26798 40864
rect 26752 40560 26798 40572
rect 14972 39786 15018 39798
rect 14972 39494 14978 39786
rect 15012 39494 15018 39786
rect 14972 39482 15018 39494
rect 16030 39786 16076 39798
rect 16030 39494 16036 39786
rect 16070 39494 16076 39786
rect 16030 39482 16076 39494
rect 17088 39786 17134 39798
rect 17088 39494 17094 39786
rect 17128 39494 17134 39786
rect 17088 39482 17134 39494
rect 18146 39786 18192 39798
rect 18146 39494 18152 39786
rect 18186 39494 18192 39786
rect 18146 39482 18192 39494
rect 19204 39786 19250 39798
rect 19204 39494 19210 39786
rect 19244 39494 19250 39786
rect 19204 39482 19250 39494
rect 20262 39786 20308 39798
rect 20262 39494 20268 39786
rect 20302 39494 20308 39786
rect 20262 39482 20308 39494
rect 14972 38692 15018 38704
rect 14972 38400 14978 38692
rect 15012 38400 15018 38692
rect 14972 38388 15018 38400
rect 16030 38692 16076 38704
rect 16030 38400 16036 38692
rect 16070 38400 16076 38692
rect 16030 38388 16076 38400
rect 17088 38692 17134 38704
rect 17088 38400 17094 38692
rect 17128 38400 17134 38692
rect 17088 38388 17134 38400
rect 18146 38692 18192 38704
rect 18146 38400 18152 38692
rect 18186 38400 18192 38692
rect 18146 38388 18192 38400
rect 19204 38692 19250 38704
rect 19204 38400 19210 38692
rect 19244 38400 19250 38692
rect 19204 38388 19250 38400
rect 20262 38692 20308 38704
rect 20262 38400 20268 38692
rect 20302 38400 20308 38692
rect 20262 38388 20308 38400
rect 14972 37252 15018 37264
rect 14972 36960 14978 37252
rect 15012 36960 15018 37252
rect 14972 36948 15018 36960
rect 16030 37252 16076 37264
rect 16030 36960 16036 37252
rect 16070 36960 16076 37252
rect 16030 36948 16076 36960
rect 17088 37252 17134 37264
rect 17088 36960 17094 37252
rect 17128 36960 17134 37252
rect 17088 36948 17134 36960
rect 18146 37252 18192 37264
rect 18146 36960 18152 37252
rect 18186 36960 18192 37252
rect 18146 36948 18192 36960
rect 19204 37252 19250 37264
rect 19204 36960 19210 37252
rect 19244 36960 19250 37252
rect 19204 36948 19250 36960
rect 20262 37252 20308 37264
rect 20262 36960 20268 37252
rect 20302 36960 20308 37252
rect 20262 36948 20308 36960
rect 14972 36158 15018 36170
rect 14972 35866 14978 36158
rect 15012 35866 15018 36158
rect 14972 35854 15018 35866
rect 16030 36158 16076 36170
rect 16030 35866 16036 36158
rect 16070 35866 16076 36158
rect 16030 35854 16076 35866
rect 17088 36158 17134 36170
rect 17088 35866 17094 36158
rect 17128 35866 17134 36158
rect 17088 35854 17134 35866
rect 18146 36158 18192 36170
rect 18146 35866 18152 36158
rect 18186 35866 18192 36158
rect 18146 35854 18192 35866
rect 19204 36158 19250 36170
rect 19204 35866 19210 36158
rect 19244 35866 19250 36158
rect 19204 35854 19250 35866
rect 20262 36158 20308 36170
rect 20262 35866 20268 36158
rect 20302 35866 20308 36158
rect 20262 35854 20308 35866
rect 8466 35056 8512 35068
rect 8466 34764 8472 35056
rect 8506 34764 8512 35056
rect 8466 34752 8512 34764
rect 9524 35056 9570 35068
rect 9524 34764 9530 35056
rect 9564 34764 9570 35056
rect 9524 34752 9570 34764
rect 10582 35056 10628 35068
rect 10582 34764 10588 35056
rect 10622 34764 10628 35056
rect 10582 34752 10628 34764
rect 11640 35056 11686 35068
rect 11640 34764 11646 35056
rect 11680 34764 11686 35056
rect 11640 34752 11686 34764
rect 12698 35056 12744 35068
rect 12698 34764 12704 35056
rect 12738 34764 12744 35056
rect 12698 34752 12744 34764
rect 13756 35056 13802 35068
rect 13756 34764 13762 35056
rect 13796 34764 13802 35056
rect 13756 34752 13802 34764
rect 1952 33954 1998 33966
rect 1952 33662 1958 33954
rect 1992 33662 1998 33954
rect 1952 33650 1998 33662
rect 3010 33954 3056 33966
rect 3010 33662 3016 33954
rect 3050 33662 3056 33954
rect 3010 33650 3056 33662
rect 4068 33954 4114 33966
rect 4068 33662 4074 33954
rect 4108 33662 4114 33954
rect 4068 33650 4114 33662
rect 5126 33954 5172 33966
rect 5126 33662 5132 33954
rect 5166 33662 5172 33954
rect 5126 33650 5172 33662
rect 6184 33954 6230 33966
rect 6184 33662 6190 33954
rect 6224 33662 6230 33954
rect 6184 33650 6230 33662
rect 7242 33954 7288 33966
rect 7242 33662 7248 33954
rect 7282 33662 7288 33954
rect 7242 33650 7288 33662
rect 1952 32860 1998 32872
rect 1952 32568 1958 32860
rect 1992 32568 1998 32860
rect 1952 32556 1998 32568
rect 3010 32860 3056 32872
rect 3010 32568 3016 32860
rect 3050 32568 3056 32860
rect 3010 32556 3056 32568
rect 4068 32860 4114 32872
rect 4068 32568 4074 32860
rect 4108 32568 4114 32860
rect 4068 32556 4114 32568
rect 5126 32860 5172 32872
rect 5126 32568 5132 32860
rect 5166 32568 5172 32860
rect 5126 32556 5172 32568
rect 6184 32860 6230 32872
rect 6184 32568 6190 32860
rect 6224 32568 6230 32860
rect 6184 32556 6230 32568
rect 7242 32860 7288 32872
rect 7242 32568 7248 32860
rect 7282 32568 7288 32860
rect 7242 32556 7288 32568
rect 1952 31402 1998 31414
rect 1952 31110 1958 31402
rect 1992 31110 1998 31402
rect 1952 31098 1998 31110
rect 3010 31402 3056 31414
rect 3010 31110 3016 31402
rect 3050 31110 3056 31402
rect 3010 31098 3056 31110
rect 4068 31402 4114 31414
rect 4068 31110 4074 31402
rect 4108 31110 4114 31402
rect 4068 31098 4114 31110
rect 5126 31402 5172 31414
rect 5126 31110 5132 31402
rect 5166 31110 5172 31402
rect 5126 31098 5172 31110
rect 6184 31402 6230 31414
rect 6184 31110 6190 31402
rect 6224 31110 6230 31402
rect 6184 31098 6230 31110
rect 7242 31402 7288 31414
rect 7242 31110 7248 31402
rect 7282 31110 7288 31402
rect 7242 31098 7288 31110
rect 1952 30308 1998 30320
rect 1952 30016 1958 30308
rect 1992 30016 1998 30308
rect 1952 30004 1998 30016
rect 3010 30308 3056 30320
rect 3010 30016 3016 30308
rect 3050 30016 3056 30308
rect 3010 30004 3056 30016
rect 4068 30308 4114 30320
rect 4068 30016 4074 30308
rect 4108 30016 4114 30308
rect 4068 30004 4114 30016
rect 5126 30308 5172 30320
rect 5126 30016 5132 30308
rect 5166 30016 5172 30308
rect 5126 30004 5172 30016
rect 6184 30308 6230 30320
rect 6184 30016 6190 30308
rect 6224 30016 6230 30308
rect 6184 30004 6230 30016
rect 7242 30308 7288 30320
rect 7242 30016 7248 30308
rect 7282 30016 7288 30308
rect 7242 30004 7288 30016
rect 1264 28672 1326 29868
rect 1420 28672 1560 29868
rect 7722 29876 8018 34514
rect 14216 34522 14346 35718
rect 14440 34522 14512 35718
rect 20748 35702 21044 40322
rect 27278 40338 27358 40970
rect 27452 40970 27486 41534
rect 33846 41540 33996 41666
rect 27452 40338 27574 40970
rect 27984 40880 28030 40892
rect 27984 40588 27990 40880
rect 28024 40588 28030 40880
rect 27984 40576 28030 40588
rect 29042 40880 29088 40892
rect 29042 40588 29048 40880
rect 29082 40588 29088 40880
rect 29042 40576 29088 40588
rect 30100 40880 30146 40892
rect 30100 40588 30106 40880
rect 30140 40588 30146 40880
rect 30100 40576 30146 40588
rect 31158 40880 31204 40892
rect 31158 40588 31164 40880
rect 31198 40588 31204 40880
rect 31158 40576 31204 40588
rect 32216 40880 32262 40892
rect 32216 40588 32222 40880
rect 32256 40588 32262 40880
rect 32216 40576 32262 40588
rect 33274 40880 33320 40892
rect 33274 40588 33280 40880
rect 33314 40588 33320 40880
rect 33274 40576 33320 40588
rect 21462 39770 21508 39782
rect 21462 39478 21468 39770
rect 21502 39478 21508 39770
rect 21462 39466 21508 39478
rect 22520 39770 22566 39782
rect 22520 39478 22526 39770
rect 22560 39478 22566 39770
rect 22520 39466 22566 39478
rect 23578 39770 23624 39782
rect 23578 39478 23584 39770
rect 23618 39478 23624 39770
rect 23578 39466 23624 39478
rect 24636 39770 24682 39782
rect 24636 39478 24642 39770
rect 24676 39478 24682 39770
rect 24636 39466 24682 39478
rect 25694 39770 25740 39782
rect 25694 39478 25700 39770
rect 25734 39478 25740 39770
rect 25694 39466 25740 39478
rect 26752 39770 26798 39782
rect 26752 39478 26758 39770
rect 26792 39478 26798 39770
rect 26752 39466 26798 39478
rect 21462 38676 21508 38688
rect 21462 38384 21468 38676
rect 21502 38384 21508 38676
rect 21462 38372 21508 38384
rect 22520 38676 22566 38688
rect 22520 38384 22526 38676
rect 22560 38384 22566 38676
rect 22520 38372 22566 38384
rect 23578 38676 23624 38688
rect 23578 38384 23584 38676
rect 23618 38384 23624 38676
rect 23578 38372 23624 38384
rect 24636 38676 24682 38688
rect 24636 38384 24642 38676
rect 24676 38384 24682 38676
rect 24636 38372 24682 38384
rect 25694 38676 25740 38688
rect 25694 38384 25700 38676
rect 25734 38384 25740 38676
rect 25694 38372 25740 38384
rect 26752 38676 26798 38688
rect 26752 38384 26758 38676
rect 26792 38384 26798 38676
rect 26752 38372 26798 38384
rect 21462 37236 21508 37248
rect 21462 36944 21468 37236
rect 21502 36944 21508 37236
rect 21462 36932 21508 36944
rect 22520 37236 22566 37248
rect 22520 36944 22526 37236
rect 22560 36944 22566 37236
rect 22520 36932 22566 36944
rect 23578 37236 23624 37248
rect 23578 36944 23584 37236
rect 23618 36944 23624 37236
rect 23578 36932 23624 36944
rect 24636 37236 24682 37248
rect 24636 36944 24642 37236
rect 24676 36944 24682 37236
rect 24636 36932 24682 36944
rect 25694 37236 25740 37248
rect 25694 36944 25700 37236
rect 25734 36944 25740 37236
rect 25694 36932 25740 36944
rect 26752 37236 26798 37248
rect 26752 36944 26758 37236
rect 26792 36944 26798 37236
rect 26752 36932 26798 36944
rect 21462 36142 21508 36154
rect 21462 35850 21468 36142
rect 21502 35850 21508 36142
rect 21462 35838 21508 35850
rect 22520 36142 22566 36154
rect 22520 35850 22526 36142
rect 22560 35850 22566 36142
rect 22520 35838 22566 35850
rect 23578 36142 23624 36154
rect 23578 35850 23584 36142
rect 23618 35850 23624 36142
rect 23578 35838 23624 35850
rect 24636 36142 24682 36154
rect 24636 35850 24642 36142
rect 24676 35850 24682 36142
rect 24636 35838 24682 35850
rect 25694 36142 25740 36154
rect 25694 35850 25700 36142
rect 25734 35850 25740 36142
rect 25694 35838 25740 35850
rect 26752 36142 26798 36154
rect 26752 35850 26758 36142
rect 26792 35850 26798 36142
rect 26752 35838 26798 35850
rect 14972 35064 15018 35076
rect 14972 34772 14978 35064
rect 15012 34772 15018 35064
rect 14972 34760 15018 34772
rect 16030 35064 16076 35076
rect 16030 34772 16036 35064
rect 16070 34772 16076 35064
rect 16030 34760 16076 34772
rect 17088 35064 17134 35076
rect 17088 34772 17094 35064
rect 17128 34772 17134 35064
rect 17088 34760 17134 34772
rect 18146 35064 18192 35076
rect 18146 34772 18152 35064
rect 18186 34772 18192 35064
rect 18146 34760 18192 34772
rect 19204 35064 19250 35076
rect 19204 34772 19210 35064
rect 19244 34772 19250 35064
rect 19204 34760 19250 34772
rect 20262 35064 20308 35076
rect 20262 34772 20268 35064
rect 20302 34772 20308 35064
rect 20262 34760 20308 34772
rect 8466 33962 8512 33974
rect 8466 33670 8472 33962
rect 8506 33670 8512 33962
rect 8466 33658 8512 33670
rect 9524 33962 9570 33974
rect 9524 33670 9530 33962
rect 9564 33670 9570 33962
rect 9524 33658 9570 33670
rect 10582 33962 10628 33974
rect 10582 33670 10588 33962
rect 10622 33670 10628 33962
rect 10582 33658 10628 33670
rect 11640 33962 11686 33974
rect 11640 33670 11646 33962
rect 11680 33670 11686 33962
rect 11640 33658 11686 33670
rect 12698 33962 12744 33974
rect 12698 33670 12704 33962
rect 12738 33670 12744 33962
rect 12698 33658 12744 33670
rect 13756 33962 13802 33974
rect 13756 33670 13762 33962
rect 13796 33670 13802 33962
rect 13756 33658 13802 33670
rect 8466 32868 8512 32880
rect 8466 32576 8472 32868
rect 8506 32576 8512 32868
rect 8466 32564 8512 32576
rect 9524 32868 9570 32880
rect 9524 32576 9530 32868
rect 9564 32576 9570 32868
rect 9524 32564 9570 32576
rect 10582 32868 10628 32880
rect 10582 32576 10588 32868
rect 10622 32576 10628 32868
rect 10582 32564 10628 32576
rect 11640 32868 11686 32880
rect 11640 32576 11646 32868
rect 11680 32576 11686 32868
rect 11640 32564 11686 32576
rect 12698 32868 12744 32880
rect 12698 32576 12704 32868
rect 12738 32576 12744 32868
rect 12698 32564 12744 32576
rect 13756 32868 13802 32880
rect 13756 32576 13762 32868
rect 13796 32576 13802 32868
rect 13756 32564 13802 32576
rect 8466 31410 8512 31422
rect 8466 31118 8472 31410
rect 8506 31118 8512 31410
rect 8466 31106 8512 31118
rect 9524 31410 9570 31422
rect 9524 31118 9530 31410
rect 9564 31118 9570 31410
rect 9524 31106 9570 31118
rect 10582 31410 10628 31422
rect 10582 31118 10588 31410
rect 10622 31118 10628 31410
rect 10582 31106 10628 31118
rect 11640 31410 11686 31422
rect 11640 31118 11646 31410
rect 11680 31118 11686 31410
rect 11640 31106 11686 31118
rect 12698 31410 12744 31422
rect 12698 31118 12704 31410
rect 12738 31118 12744 31410
rect 12698 31106 12744 31118
rect 13756 31410 13802 31422
rect 13756 31118 13762 31410
rect 13796 31118 13802 31410
rect 13756 31106 13802 31118
rect 8466 30316 8512 30328
rect 8466 30024 8472 30316
rect 8506 30024 8512 30316
rect 8466 30012 8512 30024
rect 9524 30316 9570 30328
rect 9524 30024 9530 30316
rect 9564 30024 9570 30316
rect 9524 30012 9570 30024
rect 10582 30316 10628 30328
rect 10582 30024 10588 30316
rect 10622 30024 10628 30316
rect 10582 30012 10628 30024
rect 11640 30316 11686 30328
rect 11640 30024 11646 30316
rect 11680 30024 11686 30316
rect 11640 30012 11686 30024
rect 12698 30316 12744 30328
rect 12698 30024 12704 30316
rect 12738 30024 12744 30316
rect 12698 30012 12744 30024
rect 13756 30316 13802 30328
rect 13756 30024 13762 30316
rect 13796 30024 13802 30316
rect 13756 30012 13802 30024
rect 1952 29214 1998 29226
rect 1952 28922 1958 29214
rect 1992 28922 1998 29214
rect 1952 28910 1998 28922
rect 3010 29214 3056 29226
rect 3010 28922 3016 29214
rect 3050 28922 3056 29214
rect 3010 28910 3056 28922
rect 4068 29214 4114 29226
rect 4068 28922 4074 29214
rect 4108 28922 4114 29214
rect 4068 28910 4114 28922
rect 5126 29214 5172 29226
rect 5126 28922 5132 29214
rect 5166 28922 5172 29214
rect 5126 28910 5172 28922
rect 6184 29214 6230 29226
rect 6184 28922 6190 29214
rect 6224 28922 6230 29214
rect 6184 28910 6230 28922
rect 7242 29214 7288 29226
rect 7242 28922 7248 29214
rect 7282 28922 7288 29214
rect 7242 28910 7288 28922
rect 1264 24032 1560 28672
rect 7722 28680 7840 29876
rect 7934 28680 8018 29876
rect 14216 29884 14512 34522
rect 20748 34506 20836 35702
rect 20930 34506 21044 35702
rect 27278 35718 27574 40338
rect 33846 40344 33868 41540
rect 33962 40896 33996 41540
rect 40336 41540 40486 41666
rect 40336 41156 40358 41540
rect 33962 40344 34144 40896
rect 34494 40886 34540 40898
rect 34494 40594 34500 40886
rect 34534 40594 34540 40886
rect 34494 40582 34540 40594
rect 35552 40886 35598 40898
rect 35552 40594 35558 40886
rect 35592 40594 35598 40886
rect 35552 40582 35598 40594
rect 36610 40886 36656 40898
rect 36610 40594 36616 40886
rect 36650 40594 36656 40886
rect 36610 40582 36656 40594
rect 37668 40886 37714 40898
rect 37668 40594 37674 40886
rect 37708 40594 37714 40886
rect 37668 40582 37714 40594
rect 38726 40886 38772 40898
rect 38726 40594 38732 40886
rect 38766 40594 38772 40886
rect 38726 40582 38772 40594
rect 39784 40886 39830 40898
rect 39784 40594 39790 40886
rect 39824 40594 39830 40886
rect 39784 40582 39830 40594
rect 33846 40020 34144 40344
rect 27984 39786 28030 39798
rect 27984 39494 27990 39786
rect 28024 39494 28030 39786
rect 27984 39482 28030 39494
rect 29042 39786 29088 39798
rect 29042 39494 29048 39786
rect 29082 39494 29088 39786
rect 29042 39482 29088 39494
rect 30100 39786 30146 39798
rect 30100 39494 30106 39786
rect 30140 39494 30146 39786
rect 30100 39482 30146 39494
rect 31158 39786 31204 39798
rect 31158 39494 31164 39786
rect 31198 39494 31204 39786
rect 31158 39482 31204 39494
rect 32216 39786 32262 39798
rect 32216 39494 32222 39786
rect 32256 39494 32262 39786
rect 32216 39482 32262 39494
rect 33274 39786 33320 39798
rect 33274 39494 33280 39786
rect 33314 39494 33320 39786
rect 33274 39482 33320 39494
rect 27984 38692 28030 38704
rect 27984 38400 27990 38692
rect 28024 38400 28030 38692
rect 27984 38388 28030 38400
rect 29042 38692 29088 38704
rect 29042 38400 29048 38692
rect 29082 38400 29088 38692
rect 29042 38388 29088 38400
rect 30100 38692 30146 38704
rect 30100 38400 30106 38692
rect 30140 38400 30146 38692
rect 30100 38388 30146 38400
rect 31158 38692 31204 38704
rect 31158 38400 31164 38692
rect 31198 38400 31204 38692
rect 31158 38388 31204 38400
rect 32216 38692 32262 38704
rect 32216 38400 32222 38692
rect 32256 38400 32262 38692
rect 32216 38388 32262 38400
rect 33274 38692 33320 38704
rect 33274 38400 33280 38692
rect 33314 38400 33320 38692
rect 33274 38388 33320 38400
rect 27984 37252 28030 37264
rect 27984 36960 27990 37252
rect 28024 36960 28030 37252
rect 27984 36948 28030 36960
rect 29042 37252 29088 37264
rect 29042 36960 29048 37252
rect 29082 36960 29088 37252
rect 29042 36948 29088 36960
rect 30100 37252 30146 37264
rect 30100 36960 30106 37252
rect 30140 36960 30146 37252
rect 30100 36948 30146 36960
rect 31158 37252 31204 37264
rect 31158 36960 31164 37252
rect 31198 36960 31204 37252
rect 31158 36948 31204 36960
rect 32216 37252 32262 37264
rect 32216 36960 32222 37252
rect 32256 36960 32262 37252
rect 32216 36948 32262 36960
rect 33274 37252 33320 37264
rect 33274 36960 33280 37252
rect 33314 36960 33320 37252
rect 33274 36948 33320 36960
rect 27984 36158 28030 36170
rect 27984 35866 27990 36158
rect 28024 35866 28030 36158
rect 27984 35854 28030 35866
rect 29042 36158 29088 36170
rect 29042 35866 29048 36158
rect 29082 35866 29088 36158
rect 29042 35854 29088 35866
rect 30100 36158 30146 36170
rect 30100 35866 30106 36158
rect 30140 35866 30146 36158
rect 30100 35854 30146 35866
rect 31158 36158 31204 36170
rect 31158 35866 31164 36158
rect 31198 35866 31204 36158
rect 31158 35854 31204 35866
rect 32216 36158 32262 36170
rect 32216 35866 32222 36158
rect 32256 35866 32262 36158
rect 32216 35854 32262 35866
rect 33274 36158 33320 36170
rect 33274 35866 33280 36158
rect 33314 35866 33320 36158
rect 33274 35854 33320 35866
rect 33848 35850 34144 40020
rect 40304 40344 40358 41156
rect 40452 41156 40486 41540
rect 46924 41562 47074 41688
rect 40452 40344 40638 41156
rect 40984 40886 41030 40898
rect 40984 40594 40990 40886
rect 41024 40594 41030 40886
rect 40984 40582 41030 40594
rect 42042 40886 42088 40898
rect 42042 40594 42048 40886
rect 42082 40594 42088 40886
rect 42042 40582 42088 40594
rect 43100 40886 43146 40898
rect 43100 40594 43106 40886
rect 43140 40594 43146 40886
rect 43100 40582 43146 40594
rect 44158 40886 44204 40898
rect 44158 40594 44164 40886
rect 44198 40594 44204 40886
rect 44158 40582 44204 40594
rect 45216 40886 45262 40898
rect 45216 40594 45222 40886
rect 45256 40594 45262 40886
rect 45216 40582 45262 40594
rect 46274 40886 46320 40898
rect 46274 40594 46280 40886
rect 46314 40594 46320 40886
rect 46924 40858 46946 41562
rect 46274 40582 46320 40594
rect 34494 39792 34540 39804
rect 34494 39500 34500 39792
rect 34534 39500 34540 39792
rect 34494 39488 34540 39500
rect 35552 39792 35598 39804
rect 35552 39500 35558 39792
rect 35592 39500 35598 39792
rect 35552 39488 35598 39500
rect 36610 39792 36656 39804
rect 36610 39500 36616 39792
rect 36650 39500 36656 39792
rect 36610 39488 36656 39500
rect 37668 39792 37714 39804
rect 37668 39500 37674 39792
rect 37708 39500 37714 39792
rect 37668 39488 37714 39500
rect 38726 39792 38772 39804
rect 38726 39500 38732 39792
rect 38766 39500 38772 39792
rect 38726 39488 38772 39500
rect 39784 39792 39830 39804
rect 39784 39500 39790 39792
rect 39824 39500 39830 39792
rect 39784 39488 39830 39500
rect 34494 38698 34540 38710
rect 34494 38406 34500 38698
rect 34534 38406 34540 38698
rect 34494 38394 34540 38406
rect 35552 38698 35598 38710
rect 35552 38406 35558 38698
rect 35592 38406 35598 38698
rect 35552 38394 35598 38406
rect 36610 38698 36656 38710
rect 36610 38406 36616 38698
rect 36650 38406 36656 38698
rect 36610 38394 36656 38406
rect 37668 38698 37714 38710
rect 37668 38406 37674 38698
rect 37708 38406 37714 38698
rect 37668 38394 37714 38406
rect 38726 38698 38772 38710
rect 38726 38406 38732 38698
rect 38766 38406 38772 38698
rect 38726 38394 38772 38406
rect 39784 38698 39830 38710
rect 39784 38406 39790 38698
rect 39824 38406 39830 38698
rect 39784 38394 39830 38406
rect 34494 37258 34540 37270
rect 34494 36966 34500 37258
rect 34534 36966 34540 37258
rect 34494 36954 34540 36966
rect 35552 37258 35598 37270
rect 35552 36966 35558 37258
rect 35592 36966 35598 37258
rect 35552 36954 35598 36966
rect 36610 37258 36656 37270
rect 36610 36966 36616 37258
rect 36650 36966 36656 37258
rect 36610 36954 36656 36966
rect 37668 37258 37714 37270
rect 37668 36966 37674 37258
rect 37708 36966 37714 37258
rect 37668 36954 37714 36966
rect 38726 37258 38772 37270
rect 38726 36966 38732 37258
rect 38766 36966 38772 37258
rect 38726 36954 38772 36966
rect 39784 37258 39830 37270
rect 39784 36966 39790 37258
rect 39824 36966 39830 37258
rect 39784 36954 39830 36966
rect 34494 36164 34540 36176
rect 34494 35872 34500 36164
rect 34534 35872 34540 36164
rect 34494 35860 34540 35872
rect 35552 36164 35598 36176
rect 35552 35872 35558 36164
rect 35592 35872 35598 36164
rect 35552 35860 35598 35872
rect 36610 36164 36656 36176
rect 36610 35872 36616 36164
rect 36650 35872 36656 36164
rect 36610 35860 36656 35872
rect 37668 36164 37714 36176
rect 37668 35872 37674 36164
rect 37708 35872 37714 36164
rect 37668 35860 37714 35872
rect 38726 36164 38772 36176
rect 38726 35872 38732 36164
rect 38766 35872 38772 36164
rect 38726 35860 38772 35872
rect 39784 36164 39830 36176
rect 39784 35872 39790 36164
rect 39824 35872 39830 36164
rect 39784 35860 39830 35872
rect 21462 35048 21508 35060
rect 21462 34756 21468 35048
rect 21502 34756 21508 35048
rect 21462 34744 21508 34756
rect 22520 35048 22566 35060
rect 22520 34756 22526 35048
rect 22560 34756 22566 35048
rect 22520 34744 22566 34756
rect 23578 35048 23624 35060
rect 23578 34756 23584 35048
rect 23618 34756 23624 35048
rect 23578 34744 23624 34756
rect 24636 35048 24682 35060
rect 24636 34756 24642 35048
rect 24676 34756 24682 35048
rect 24636 34744 24682 34756
rect 25694 35048 25740 35060
rect 25694 34756 25700 35048
rect 25734 34756 25740 35048
rect 25694 34744 25740 34756
rect 26752 35048 26798 35060
rect 26752 34756 26758 35048
rect 26792 34756 26798 35048
rect 26752 34744 26798 34756
rect 14972 33970 15018 33982
rect 14972 33678 14978 33970
rect 15012 33678 15018 33970
rect 14972 33666 15018 33678
rect 16030 33970 16076 33982
rect 16030 33678 16036 33970
rect 16070 33678 16076 33970
rect 16030 33666 16076 33678
rect 17088 33970 17134 33982
rect 17088 33678 17094 33970
rect 17128 33678 17134 33970
rect 17088 33666 17134 33678
rect 18146 33970 18192 33982
rect 18146 33678 18152 33970
rect 18186 33678 18192 33970
rect 18146 33666 18192 33678
rect 19204 33970 19250 33982
rect 19204 33678 19210 33970
rect 19244 33678 19250 33970
rect 19204 33666 19250 33678
rect 20262 33970 20308 33982
rect 20262 33678 20268 33970
rect 20302 33678 20308 33970
rect 20262 33666 20308 33678
rect 14972 32876 15018 32888
rect 14972 32584 14978 32876
rect 15012 32584 15018 32876
rect 14972 32572 15018 32584
rect 16030 32876 16076 32888
rect 16030 32584 16036 32876
rect 16070 32584 16076 32876
rect 16030 32572 16076 32584
rect 17088 32876 17134 32888
rect 17088 32584 17094 32876
rect 17128 32584 17134 32876
rect 17088 32572 17134 32584
rect 18146 32876 18192 32888
rect 18146 32584 18152 32876
rect 18186 32584 18192 32876
rect 18146 32572 18192 32584
rect 19204 32876 19250 32888
rect 19204 32584 19210 32876
rect 19244 32584 19250 32876
rect 19204 32572 19250 32584
rect 20262 32876 20308 32888
rect 20262 32584 20268 32876
rect 20302 32584 20308 32876
rect 20262 32572 20308 32584
rect 14972 31418 15018 31430
rect 14972 31126 14978 31418
rect 15012 31126 15018 31418
rect 14972 31114 15018 31126
rect 16030 31418 16076 31430
rect 16030 31126 16036 31418
rect 16070 31126 16076 31418
rect 16030 31114 16076 31126
rect 17088 31418 17134 31430
rect 17088 31126 17094 31418
rect 17128 31126 17134 31418
rect 17088 31114 17134 31126
rect 18146 31418 18192 31430
rect 18146 31126 18152 31418
rect 18186 31126 18192 31418
rect 18146 31114 18192 31126
rect 19204 31418 19250 31430
rect 19204 31126 19210 31418
rect 19244 31126 19250 31418
rect 19204 31114 19250 31126
rect 20262 31418 20308 31430
rect 20262 31126 20268 31418
rect 20302 31126 20308 31418
rect 20262 31114 20308 31126
rect 14972 30324 15018 30336
rect 14972 30032 14978 30324
rect 15012 30032 15018 30324
rect 14972 30020 15018 30032
rect 16030 30324 16076 30336
rect 16030 30032 16036 30324
rect 16070 30032 16076 30324
rect 16030 30020 16076 30032
rect 17088 30324 17134 30336
rect 17088 30032 17094 30324
rect 17128 30032 17134 30324
rect 17088 30020 17134 30032
rect 18146 30324 18192 30336
rect 18146 30032 18152 30324
rect 18186 30032 18192 30324
rect 18146 30020 18192 30032
rect 19204 30324 19250 30336
rect 19204 30032 19210 30324
rect 19244 30032 19250 30324
rect 19204 30020 19250 30032
rect 20262 30324 20308 30336
rect 20262 30032 20268 30324
rect 20302 30032 20308 30324
rect 20262 30020 20308 30032
rect 8466 29222 8512 29234
rect 8466 28930 8472 29222
rect 8506 28930 8512 29222
rect 8466 28918 8512 28930
rect 9524 29222 9570 29234
rect 9524 28930 9530 29222
rect 9564 28930 9570 29222
rect 9524 28918 9570 28930
rect 10582 29222 10628 29234
rect 10582 28930 10588 29222
rect 10622 28930 10628 29222
rect 10582 28918 10628 28930
rect 11640 29222 11686 29234
rect 11640 28930 11646 29222
rect 11680 28930 11686 29222
rect 11640 28918 11686 28930
rect 12698 29222 12744 29234
rect 12698 28930 12704 29222
rect 12738 28930 12744 29222
rect 12698 28918 12744 28930
rect 13756 29222 13802 29234
rect 13756 28930 13762 29222
rect 13796 28930 13802 29222
rect 13756 28918 13802 28930
rect 1952 28120 1998 28132
rect 1952 27828 1958 28120
rect 1992 27828 1998 28120
rect 1952 27816 1998 27828
rect 3010 28120 3056 28132
rect 3010 27828 3016 28120
rect 3050 27828 3056 28120
rect 3010 27816 3056 27828
rect 4068 28120 4114 28132
rect 4068 27828 4074 28120
rect 4108 27828 4114 28120
rect 4068 27816 4114 27828
rect 5126 28120 5172 28132
rect 5126 27828 5132 28120
rect 5166 27828 5172 28120
rect 5126 27816 5172 27828
rect 6184 28120 6230 28132
rect 6184 27828 6190 28120
rect 6224 27828 6230 28120
rect 6184 27816 6230 27828
rect 7242 28120 7288 28132
rect 7242 27828 7248 28120
rect 7282 27828 7288 28120
rect 7242 27816 7288 27828
rect 1952 27026 1998 27038
rect 1952 26734 1958 27026
rect 1992 26734 1998 27026
rect 1952 26722 1998 26734
rect 3010 27026 3056 27038
rect 3010 26734 3016 27026
rect 3050 26734 3056 27026
rect 3010 26722 3056 26734
rect 4068 27026 4114 27038
rect 4068 26734 4074 27026
rect 4108 26734 4114 27026
rect 4068 26722 4114 26734
rect 5126 27026 5172 27038
rect 5126 26734 5132 27026
rect 5166 26734 5172 27026
rect 5126 26722 5172 26734
rect 6184 27026 6230 27038
rect 6184 26734 6190 27026
rect 6224 26734 6230 27026
rect 6184 26722 6230 26734
rect 7242 27026 7288 27038
rect 7242 26734 7248 27026
rect 7282 26734 7288 27026
rect 7242 26722 7288 26734
rect 1952 25566 1998 25578
rect 1952 25274 1958 25566
rect 1992 25274 1998 25566
rect 1952 25262 1998 25274
rect 3010 25566 3056 25578
rect 3010 25274 3016 25566
rect 3050 25274 3056 25566
rect 3010 25262 3056 25274
rect 4068 25566 4114 25578
rect 4068 25274 4074 25566
rect 4108 25274 4114 25566
rect 4068 25262 4114 25274
rect 5126 25566 5172 25578
rect 5126 25274 5132 25566
rect 5166 25274 5172 25566
rect 5126 25262 5172 25274
rect 6184 25566 6230 25578
rect 6184 25274 6190 25566
rect 6224 25274 6230 25566
rect 6184 25262 6230 25274
rect 7242 25566 7288 25578
rect 7242 25274 7248 25566
rect 7282 25274 7288 25566
rect 7242 25262 7288 25274
rect 1952 24472 1998 24484
rect 1952 24180 1958 24472
rect 1992 24180 1998 24472
rect 1952 24168 1998 24180
rect 3010 24472 3056 24484
rect 3010 24180 3016 24472
rect 3050 24180 3056 24472
rect 3010 24168 3056 24180
rect 4068 24472 4114 24484
rect 4068 24180 4074 24472
rect 4108 24180 4114 24472
rect 4068 24168 4114 24180
rect 5126 24472 5172 24484
rect 5126 24180 5132 24472
rect 5166 24180 5172 24472
rect 5126 24168 5172 24180
rect 6184 24472 6230 24484
rect 6184 24180 6190 24472
rect 6224 24180 6230 24472
rect 6184 24168 6230 24180
rect 7242 24472 7288 24484
rect 7242 24180 7248 24472
rect 7282 24180 7288 24472
rect 7242 24168 7288 24180
rect 1264 22836 1326 24032
rect 1420 22836 1560 24032
rect 7722 24040 8018 28680
rect 14216 28688 14346 29884
rect 14440 28688 14512 29884
rect 20748 29868 21044 34506
rect 27278 34522 27358 35718
rect 27452 34522 27574 35718
rect 33846 35724 34144 35850
rect 27984 35064 28030 35076
rect 27984 34772 27990 35064
rect 28024 34772 28030 35064
rect 27984 34760 28030 34772
rect 29042 35064 29088 35076
rect 29042 34772 29048 35064
rect 29082 34772 29088 35064
rect 29042 34760 29088 34772
rect 30100 35064 30146 35076
rect 30100 34772 30106 35064
rect 30140 34772 30146 35064
rect 30100 34760 30146 34772
rect 31158 35064 31204 35076
rect 31158 34772 31164 35064
rect 31198 34772 31204 35064
rect 31158 34760 31204 34772
rect 32216 35064 32262 35076
rect 32216 34772 32222 35064
rect 32256 34772 32262 35064
rect 32216 34760 32262 34772
rect 33274 35064 33320 35076
rect 33274 34772 33280 35064
rect 33314 34772 33320 35064
rect 33274 34760 33320 34772
rect 21462 33954 21508 33966
rect 21462 33662 21468 33954
rect 21502 33662 21508 33954
rect 21462 33650 21508 33662
rect 22520 33954 22566 33966
rect 22520 33662 22526 33954
rect 22560 33662 22566 33954
rect 22520 33650 22566 33662
rect 23578 33954 23624 33966
rect 23578 33662 23584 33954
rect 23618 33662 23624 33954
rect 23578 33650 23624 33662
rect 24636 33954 24682 33966
rect 24636 33662 24642 33954
rect 24676 33662 24682 33954
rect 24636 33650 24682 33662
rect 25694 33954 25740 33966
rect 25694 33662 25700 33954
rect 25734 33662 25740 33954
rect 25694 33650 25740 33662
rect 26752 33954 26798 33966
rect 26752 33662 26758 33954
rect 26792 33662 26798 33954
rect 26752 33650 26798 33662
rect 21462 32860 21508 32872
rect 21462 32568 21468 32860
rect 21502 32568 21508 32860
rect 21462 32556 21508 32568
rect 22520 32860 22566 32872
rect 22520 32568 22526 32860
rect 22560 32568 22566 32860
rect 22520 32556 22566 32568
rect 23578 32860 23624 32872
rect 23578 32568 23584 32860
rect 23618 32568 23624 32860
rect 23578 32556 23624 32568
rect 24636 32860 24682 32872
rect 24636 32568 24642 32860
rect 24676 32568 24682 32860
rect 24636 32556 24682 32568
rect 25694 32860 25740 32872
rect 25694 32568 25700 32860
rect 25734 32568 25740 32860
rect 25694 32556 25740 32568
rect 26752 32860 26798 32872
rect 26752 32568 26758 32860
rect 26792 32568 26798 32860
rect 26752 32556 26798 32568
rect 21462 31402 21508 31414
rect 21462 31110 21468 31402
rect 21502 31110 21508 31402
rect 21462 31098 21508 31110
rect 22520 31402 22566 31414
rect 22520 31110 22526 31402
rect 22560 31110 22566 31402
rect 22520 31098 22566 31110
rect 23578 31402 23624 31414
rect 23578 31110 23584 31402
rect 23618 31110 23624 31402
rect 23578 31098 23624 31110
rect 24636 31402 24682 31414
rect 24636 31110 24642 31402
rect 24676 31110 24682 31402
rect 24636 31098 24682 31110
rect 25694 31402 25740 31414
rect 25694 31110 25700 31402
rect 25734 31110 25740 31402
rect 25694 31098 25740 31110
rect 26752 31402 26798 31414
rect 26752 31110 26758 31402
rect 26792 31110 26798 31402
rect 26752 31098 26798 31110
rect 21462 30308 21508 30320
rect 21462 30016 21468 30308
rect 21502 30016 21508 30308
rect 21462 30004 21508 30016
rect 22520 30308 22566 30320
rect 22520 30016 22526 30308
rect 22560 30016 22566 30308
rect 22520 30004 22566 30016
rect 23578 30308 23624 30320
rect 23578 30016 23584 30308
rect 23618 30016 23624 30308
rect 23578 30004 23624 30016
rect 24636 30308 24682 30320
rect 24636 30016 24642 30308
rect 24676 30016 24682 30308
rect 24636 30004 24682 30016
rect 25694 30308 25740 30320
rect 25694 30016 25700 30308
rect 25734 30016 25740 30308
rect 25694 30004 25740 30016
rect 26752 30308 26798 30320
rect 26752 30016 26758 30308
rect 26792 30016 26798 30308
rect 26752 30004 26798 30016
rect 14972 29230 15018 29242
rect 14972 28938 14978 29230
rect 15012 28938 15018 29230
rect 14972 28926 15018 28938
rect 16030 29230 16076 29242
rect 16030 28938 16036 29230
rect 16070 28938 16076 29230
rect 16030 28926 16076 28938
rect 17088 29230 17134 29242
rect 17088 28938 17094 29230
rect 17128 28938 17134 29230
rect 17088 28926 17134 28938
rect 18146 29230 18192 29242
rect 18146 28938 18152 29230
rect 18186 28938 18192 29230
rect 18146 28926 18192 28938
rect 19204 29230 19250 29242
rect 19204 28938 19210 29230
rect 19244 28938 19250 29230
rect 19204 28926 19250 28938
rect 20262 29230 20308 29242
rect 20262 28938 20268 29230
rect 20302 28938 20308 29230
rect 20262 28926 20308 28938
rect 8466 28128 8512 28140
rect 8466 27836 8472 28128
rect 8506 27836 8512 28128
rect 8466 27824 8512 27836
rect 9524 28128 9570 28140
rect 9524 27836 9530 28128
rect 9564 27836 9570 28128
rect 9524 27824 9570 27836
rect 10582 28128 10628 28140
rect 10582 27836 10588 28128
rect 10622 27836 10628 28128
rect 10582 27824 10628 27836
rect 11640 28128 11686 28140
rect 11640 27836 11646 28128
rect 11680 27836 11686 28128
rect 11640 27824 11686 27836
rect 12698 28128 12744 28140
rect 12698 27836 12704 28128
rect 12738 27836 12744 28128
rect 12698 27824 12744 27836
rect 13756 28128 13802 28140
rect 13756 27836 13762 28128
rect 13796 27836 13802 28128
rect 13756 27824 13802 27836
rect 8466 27034 8512 27046
rect 8466 26742 8472 27034
rect 8506 26742 8512 27034
rect 8466 26730 8512 26742
rect 9524 27034 9570 27046
rect 9524 26742 9530 27034
rect 9564 26742 9570 27034
rect 9524 26730 9570 26742
rect 10582 27034 10628 27046
rect 10582 26742 10588 27034
rect 10622 26742 10628 27034
rect 10582 26730 10628 26742
rect 11640 27034 11686 27046
rect 11640 26742 11646 27034
rect 11680 26742 11686 27034
rect 11640 26730 11686 26742
rect 12698 27034 12744 27046
rect 12698 26742 12704 27034
rect 12738 26742 12744 27034
rect 12698 26730 12744 26742
rect 13756 27034 13802 27046
rect 13756 26742 13762 27034
rect 13796 26742 13802 27034
rect 13756 26730 13802 26742
rect 8466 25574 8512 25586
rect 8466 25282 8472 25574
rect 8506 25282 8512 25574
rect 8466 25270 8512 25282
rect 9524 25574 9570 25586
rect 9524 25282 9530 25574
rect 9564 25282 9570 25574
rect 9524 25270 9570 25282
rect 10582 25574 10628 25586
rect 10582 25282 10588 25574
rect 10622 25282 10628 25574
rect 10582 25270 10628 25282
rect 11640 25574 11686 25586
rect 11640 25282 11646 25574
rect 11680 25282 11686 25574
rect 11640 25270 11686 25282
rect 12698 25574 12744 25586
rect 12698 25282 12704 25574
rect 12738 25282 12744 25574
rect 12698 25270 12744 25282
rect 13756 25574 13802 25586
rect 13756 25282 13762 25574
rect 13796 25282 13802 25574
rect 13756 25270 13802 25282
rect 8466 24480 8512 24492
rect 8466 24188 8472 24480
rect 8506 24188 8512 24480
rect 8466 24176 8512 24188
rect 9524 24480 9570 24492
rect 9524 24188 9530 24480
rect 9564 24188 9570 24480
rect 9524 24176 9570 24188
rect 10582 24480 10628 24492
rect 10582 24188 10588 24480
rect 10622 24188 10628 24480
rect 10582 24176 10628 24188
rect 11640 24480 11686 24492
rect 11640 24188 11646 24480
rect 11680 24188 11686 24480
rect 11640 24176 11686 24188
rect 12698 24480 12744 24492
rect 12698 24188 12704 24480
rect 12738 24188 12744 24480
rect 12698 24176 12744 24188
rect 13756 24480 13802 24492
rect 13756 24188 13762 24480
rect 13796 24188 13802 24480
rect 13756 24176 13802 24188
rect 1952 23378 1998 23390
rect 1952 23086 1958 23378
rect 1992 23086 1998 23378
rect 1952 23074 1998 23086
rect 3010 23378 3056 23390
rect 3010 23086 3016 23378
rect 3050 23086 3056 23378
rect 3010 23074 3056 23086
rect 4068 23378 4114 23390
rect 4068 23086 4074 23378
rect 4108 23086 4114 23378
rect 4068 23074 4114 23086
rect 5126 23378 5172 23390
rect 5126 23086 5132 23378
rect 5166 23086 5172 23378
rect 5126 23074 5172 23086
rect 6184 23378 6230 23390
rect 6184 23086 6190 23378
rect 6224 23086 6230 23378
rect 6184 23074 6230 23086
rect 7242 23378 7288 23390
rect 7242 23086 7248 23378
rect 7282 23086 7288 23378
rect 7242 23074 7288 23086
rect 1264 18168 1560 22836
rect 7722 22844 7840 24040
rect 7934 22844 8018 24040
rect 14216 24048 14512 28688
rect 20748 28672 20836 29868
rect 20930 28672 21044 29868
rect 27278 29884 27574 34522
rect 33846 34528 33868 35724
rect 33962 34528 34144 35724
rect 40304 35724 40638 40344
rect 46836 40366 46946 40858
rect 47040 40858 47074 41562
rect 53438 41576 53588 41702
rect 47572 40908 47618 40920
rect 47040 40366 47170 40858
rect 47572 40616 47578 40908
rect 47612 40616 47618 40908
rect 47572 40604 47618 40616
rect 48630 40908 48676 40920
rect 48630 40616 48636 40908
rect 48670 40616 48676 40908
rect 48630 40604 48676 40616
rect 49688 40908 49734 40920
rect 49688 40616 49694 40908
rect 49728 40616 49734 40908
rect 49688 40604 49734 40616
rect 50746 40908 50792 40920
rect 50746 40616 50752 40908
rect 50786 40616 50792 40908
rect 50746 40604 50792 40616
rect 51804 40908 51850 40920
rect 51804 40616 51810 40908
rect 51844 40616 51850 40908
rect 51804 40604 51850 40616
rect 52862 40908 52908 40920
rect 52862 40616 52868 40908
rect 52902 40616 52908 40908
rect 52862 40604 52908 40616
rect 40984 39792 41030 39804
rect 40984 39500 40990 39792
rect 41024 39500 41030 39792
rect 40984 39488 41030 39500
rect 42042 39792 42088 39804
rect 42042 39500 42048 39792
rect 42082 39500 42088 39792
rect 42042 39488 42088 39500
rect 43100 39792 43146 39804
rect 43100 39500 43106 39792
rect 43140 39500 43146 39792
rect 43100 39488 43146 39500
rect 44158 39792 44204 39804
rect 44158 39500 44164 39792
rect 44198 39500 44204 39792
rect 44158 39488 44204 39500
rect 45216 39792 45262 39804
rect 45216 39500 45222 39792
rect 45256 39500 45262 39792
rect 45216 39488 45262 39500
rect 46274 39792 46320 39804
rect 46274 39500 46280 39792
rect 46314 39500 46320 39792
rect 46274 39488 46320 39500
rect 40984 38698 41030 38710
rect 40984 38406 40990 38698
rect 41024 38406 41030 38698
rect 40984 38394 41030 38406
rect 42042 38698 42088 38710
rect 42042 38406 42048 38698
rect 42082 38406 42088 38698
rect 42042 38394 42088 38406
rect 43100 38698 43146 38710
rect 43100 38406 43106 38698
rect 43140 38406 43146 38698
rect 43100 38394 43146 38406
rect 44158 38698 44204 38710
rect 44158 38406 44164 38698
rect 44198 38406 44204 38698
rect 44158 38394 44204 38406
rect 45216 38698 45262 38710
rect 45216 38406 45222 38698
rect 45256 38406 45262 38698
rect 45216 38394 45262 38406
rect 46274 38698 46320 38710
rect 46274 38406 46280 38698
rect 46314 38406 46320 38698
rect 46274 38394 46320 38406
rect 40984 37258 41030 37270
rect 40984 36966 40990 37258
rect 41024 36966 41030 37258
rect 40984 36954 41030 36966
rect 42042 37258 42088 37270
rect 42042 36966 42048 37258
rect 42082 36966 42088 37258
rect 42042 36954 42088 36966
rect 43100 37258 43146 37270
rect 43100 36966 43106 37258
rect 43140 36966 43146 37258
rect 43100 36954 43146 36966
rect 44158 37258 44204 37270
rect 44158 36966 44164 37258
rect 44198 36966 44204 37258
rect 44158 36954 44204 36966
rect 45216 37258 45262 37270
rect 45216 36966 45222 37258
rect 45256 36966 45262 37258
rect 45216 36954 45262 36966
rect 46274 37258 46320 37270
rect 46274 36966 46280 37258
rect 46314 36966 46320 37258
rect 46274 36954 46320 36966
rect 40984 36164 41030 36176
rect 40984 35872 40990 36164
rect 41024 35872 41030 36164
rect 40984 35860 41030 35872
rect 42042 36164 42088 36176
rect 42042 35872 42048 36164
rect 42082 35872 42088 36164
rect 42042 35860 42088 35872
rect 43100 36164 43146 36176
rect 43100 35872 43106 36164
rect 43140 35872 43146 36164
rect 43100 35860 43146 35872
rect 44158 36164 44204 36176
rect 44158 35872 44164 36164
rect 44198 35872 44204 36164
rect 44158 35860 44204 35872
rect 45216 36164 45262 36176
rect 45216 35872 45222 36164
rect 45256 35872 45262 36164
rect 45216 35860 45262 35872
rect 46274 36164 46320 36176
rect 46274 35872 46280 36164
rect 46314 35872 46320 36164
rect 46274 35860 46320 35872
rect 34494 35070 34540 35082
rect 34494 34778 34500 35070
rect 34534 34778 34540 35070
rect 34494 34766 34540 34778
rect 35552 35070 35598 35082
rect 35552 34778 35558 35070
rect 35592 34778 35598 35070
rect 35552 34766 35598 34778
rect 36610 35070 36656 35082
rect 36610 34778 36616 35070
rect 36650 34778 36656 35070
rect 36610 34766 36656 34778
rect 37668 35070 37714 35082
rect 37668 34778 37674 35070
rect 37708 34778 37714 35070
rect 37668 34766 37714 34778
rect 38726 35070 38772 35082
rect 38726 34778 38732 35070
rect 38766 34778 38772 35070
rect 38726 34766 38772 34778
rect 39784 35070 39830 35082
rect 39784 34778 39790 35070
rect 39824 34778 39830 35070
rect 39784 34766 39830 34778
rect 33846 34204 34144 34528
rect 27984 33970 28030 33982
rect 27984 33678 27990 33970
rect 28024 33678 28030 33970
rect 27984 33666 28030 33678
rect 29042 33970 29088 33982
rect 29042 33678 29048 33970
rect 29082 33678 29088 33970
rect 29042 33666 29088 33678
rect 30100 33970 30146 33982
rect 30100 33678 30106 33970
rect 30140 33678 30146 33970
rect 30100 33666 30146 33678
rect 31158 33970 31204 33982
rect 31158 33678 31164 33970
rect 31198 33678 31204 33970
rect 31158 33666 31204 33678
rect 32216 33970 32262 33982
rect 32216 33678 32222 33970
rect 32256 33678 32262 33970
rect 32216 33666 32262 33678
rect 33274 33970 33320 33982
rect 33274 33678 33280 33970
rect 33314 33678 33320 33970
rect 33274 33666 33320 33678
rect 27984 32876 28030 32888
rect 27984 32584 27990 32876
rect 28024 32584 28030 32876
rect 27984 32572 28030 32584
rect 29042 32876 29088 32888
rect 29042 32584 29048 32876
rect 29082 32584 29088 32876
rect 29042 32572 29088 32584
rect 30100 32876 30146 32888
rect 30100 32584 30106 32876
rect 30140 32584 30146 32876
rect 30100 32572 30146 32584
rect 31158 32876 31204 32888
rect 31158 32584 31164 32876
rect 31198 32584 31204 32876
rect 31158 32572 31204 32584
rect 32216 32876 32262 32888
rect 32216 32584 32222 32876
rect 32256 32584 32262 32876
rect 32216 32572 32262 32584
rect 33274 32876 33320 32888
rect 33274 32584 33280 32876
rect 33314 32584 33320 32876
rect 33274 32572 33320 32584
rect 27984 31418 28030 31430
rect 27984 31126 27990 31418
rect 28024 31126 28030 31418
rect 27984 31114 28030 31126
rect 29042 31418 29088 31430
rect 29042 31126 29048 31418
rect 29082 31126 29088 31418
rect 29042 31114 29088 31126
rect 30100 31418 30146 31430
rect 30100 31126 30106 31418
rect 30140 31126 30146 31418
rect 30100 31114 30146 31126
rect 31158 31418 31204 31430
rect 31158 31126 31164 31418
rect 31198 31126 31204 31418
rect 31158 31114 31204 31126
rect 32216 31418 32262 31430
rect 32216 31126 32222 31418
rect 32256 31126 32262 31418
rect 32216 31114 32262 31126
rect 33274 31418 33320 31430
rect 33274 31126 33280 31418
rect 33314 31126 33320 31418
rect 33274 31114 33320 31126
rect 27984 30324 28030 30336
rect 27984 30032 27990 30324
rect 28024 30032 28030 30324
rect 27984 30020 28030 30032
rect 29042 30324 29088 30336
rect 29042 30032 29048 30324
rect 29082 30032 29088 30324
rect 29042 30020 29088 30032
rect 30100 30324 30146 30336
rect 30100 30032 30106 30324
rect 30140 30032 30146 30324
rect 30100 30020 30146 30032
rect 31158 30324 31204 30336
rect 31158 30032 31164 30324
rect 31198 30032 31204 30324
rect 31158 30020 31204 30032
rect 32216 30324 32262 30336
rect 32216 30032 32222 30324
rect 32256 30032 32262 30324
rect 32216 30020 32262 30032
rect 33274 30324 33320 30336
rect 33274 30032 33280 30324
rect 33314 30032 33320 30324
rect 33274 30020 33320 30032
rect 33848 30016 34144 34204
rect 40304 34528 40358 35724
rect 40452 34528 40638 35724
rect 46836 35746 47170 40366
rect 53438 40380 53460 41576
rect 53554 41008 53588 41576
rect 53554 40380 53776 41008
rect 54086 40922 54132 40934
rect 54086 40630 54092 40922
rect 54126 40630 54132 40922
rect 54086 40618 54132 40630
rect 55144 40922 55190 40934
rect 55144 40630 55150 40922
rect 55184 40630 55190 40922
rect 55144 40618 55190 40630
rect 56202 40922 56248 40934
rect 56202 40630 56208 40922
rect 56242 40630 56248 40922
rect 56202 40618 56248 40630
rect 57260 40922 57306 40934
rect 57260 40630 57266 40922
rect 57300 40630 57306 40922
rect 57260 40618 57306 40630
rect 58318 40922 58364 40934
rect 58318 40630 58324 40922
rect 58358 40630 58364 40922
rect 58318 40618 58364 40630
rect 59376 40922 59422 40934
rect 59376 40630 59382 40922
rect 59416 40630 59422 40922
rect 59376 40618 59422 40630
rect 53438 40056 53776 40380
rect 59530 40204 59572 41772
rect 59836 41292 59934 41772
rect 62148 41604 62194 42532
rect 62116 41292 62194 41604
rect 59836 41040 62194 41292
rect 59836 40204 60012 41040
rect 59530 40066 60012 40204
rect 47572 39814 47618 39826
rect 47572 39522 47578 39814
rect 47612 39522 47618 39814
rect 47572 39510 47618 39522
rect 48630 39814 48676 39826
rect 48630 39522 48636 39814
rect 48670 39522 48676 39814
rect 48630 39510 48676 39522
rect 49688 39814 49734 39826
rect 49688 39522 49694 39814
rect 49728 39522 49734 39814
rect 49688 39510 49734 39522
rect 50746 39814 50792 39826
rect 50746 39522 50752 39814
rect 50786 39522 50792 39814
rect 50746 39510 50792 39522
rect 51804 39814 51850 39826
rect 51804 39522 51810 39814
rect 51844 39522 51850 39814
rect 51804 39510 51850 39522
rect 52862 39814 52908 39826
rect 52862 39522 52868 39814
rect 52902 39522 52908 39814
rect 52862 39510 52908 39522
rect 47572 38720 47618 38732
rect 47572 38428 47578 38720
rect 47612 38428 47618 38720
rect 47572 38416 47618 38428
rect 48630 38720 48676 38732
rect 48630 38428 48636 38720
rect 48670 38428 48676 38720
rect 48630 38416 48676 38428
rect 49688 38720 49734 38732
rect 49688 38428 49694 38720
rect 49728 38428 49734 38720
rect 49688 38416 49734 38428
rect 50746 38720 50792 38732
rect 50746 38428 50752 38720
rect 50786 38428 50792 38720
rect 50746 38416 50792 38428
rect 51804 38720 51850 38732
rect 51804 38428 51810 38720
rect 51844 38428 51850 38720
rect 51804 38416 51850 38428
rect 52862 38720 52908 38732
rect 52862 38428 52868 38720
rect 52902 38428 52908 38720
rect 52862 38416 52908 38428
rect 47572 37280 47618 37292
rect 47572 36988 47578 37280
rect 47612 36988 47618 37280
rect 47572 36976 47618 36988
rect 48630 37280 48676 37292
rect 48630 36988 48636 37280
rect 48670 36988 48676 37280
rect 48630 36976 48676 36988
rect 49688 37280 49734 37292
rect 49688 36988 49694 37280
rect 49728 36988 49734 37280
rect 49688 36976 49734 36988
rect 50746 37280 50792 37292
rect 50746 36988 50752 37280
rect 50786 36988 50792 37280
rect 50746 36976 50792 36988
rect 51804 37280 51850 37292
rect 51804 36988 51810 37280
rect 51844 36988 51850 37280
rect 51804 36976 51850 36988
rect 52862 37280 52908 37292
rect 52862 36988 52868 37280
rect 52902 36988 52908 37280
rect 52862 36976 52908 36988
rect 47572 36186 47618 36198
rect 47572 35894 47578 36186
rect 47612 35894 47618 36186
rect 47572 35882 47618 35894
rect 48630 36186 48676 36198
rect 48630 35894 48636 36186
rect 48670 35894 48676 36186
rect 48630 35882 48676 35894
rect 49688 36186 49734 36198
rect 49688 35894 49694 36186
rect 49728 35894 49734 36186
rect 49688 35882 49734 35894
rect 50746 36186 50792 36198
rect 50746 35894 50752 36186
rect 50786 35894 50792 36186
rect 50746 35882 50792 35894
rect 51804 36186 51850 36198
rect 51804 35894 51810 36186
rect 51844 35894 51850 36186
rect 51804 35882 51850 35894
rect 52862 36186 52908 36198
rect 52862 35894 52868 36186
rect 52902 35894 52908 36186
rect 52862 35882 52908 35894
rect 53442 35886 53776 40056
rect 54086 39828 54132 39840
rect 54086 39536 54092 39828
rect 54126 39536 54132 39828
rect 54086 39524 54132 39536
rect 55144 39828 55190 39840
rect 55144 39536 55150 39828
rect 55184 39536 55190 39828
rect 55144 39524 55190 39536
rect 56202 39828 56248 39840
rect 56202 39536 56208 39828
rect 56242 39536 56248 39828
rect 56202 39524 56248 39536
rect 57260 39828 57306 39840
rect 57260 39536 57266 39828
rect 57300 39536 57306 39828
rect 57260 39524 57306 39536
rect 58318 39828 58364 39840
rect 58318 39536 58324 39828
rect 58358 39536 58364 39828
rect 58318 39524 58364 39536
rect 59376 39828 59422 39840
rect 59376 39536 59382 39828
rect 59416 39536 59422 39828
rect 59376 39524 59422 39536
rect 54086 38734 54132 38746
rect 54086 38442 54092 38734
rect 54126 38442 54132 38734
rect 54086 38430 54132 38442
rect 55144 38734 55190 38746
rect 55144 38442 55150 38734
rect 55184 38442 55190 38734
rect 55144 38430 55190 38442
rect 56202 38734 56248 38746
rect 56202 38442 56208 38734
rect 56242 38442 56248 38734
rect 56202 38430 56248 38442
rect 57260 38734 57306 38746
rect 57260 38442 57266 38734
rect 57300 38442 57306 38734
rect 57260 38430 57306 38442
rect 58318 38734 58364 38746
rect 58318 38442 58324 38734
rect 58358 38442 58364 38734
rect 58318 38430 58364 38442
rect 59376 38734 59422 38746
rect 59376 38442 59382 38734
rect 59416 38442 59422 38734
rect 59376 38430 59422 38442
rect 54086 37294 54132 37306
rect 54086 37002 54092 37294
rect 54126 37002 54132 37294
rect 54086 36990 54132 37002
rect 55144 37294 55190 37306
rect 55144 37002 55150 37294
rect 55184 37002 55190 37294
rect 55144 36990 55190 37002
rect 56202 37294 56248 37306
rect 56202 37002 56208 37294
rect 56242 37002 56248 37294
rect 56202 36990 56248 37002
rect 57260 37294 57306 37306
rect 57260 37002 57266 37294
rect 57300 37002 57306 37294
rect 57260 36990 57306 37002
rect 58318 37294 58364 37306
rect 58318 37002 58324 37294
rect 58358 37002 58364 37294
rect 58318 36990 58364 37002
rect 59376 37294 59422 37306
rect 59376 37002 59382 37294
rect 59416 37002 59422 37294
rect 59376 36990 59422 37002
rect 54086 36200 54132 36212
rect 54086 35908 54092 36200
rect 54126 35908 54132 36200
rect 54086 35896 54132 35908
rect 55144 36200 55190 36212
rect 55144 35908 55150 36200
rect 55184 35908 55190 36200
rect 55144 35896 55190 35908
rect 56202 36200 56248 36212
rect 56202 35908 56208 36200
rect 56242 35908 56248 36200
rect 56202 35896 56248 35908
rect 57260 36200 57306 36212
rect 57260 35908 57266 36200
rect 57300 35908 57306 36200
rect 57260 35896 57306 35908
rect 58318 36200 58364 36212
rect 58318 35908 58324 36200
rect 58358 35908 58364 36200
rect 58318 35896 58364 35908
rect 59376 36200 59422 36212
rect 59376 35908 59382 36200
rect 59416 35908 59422 36200
rect 59680 36084 60012 40066
rect 62116 41028 62194 41040
rect 62288 41028 62360 42532
rect 65942 42534 66154 42702
rect 62502 42414 62548 42426
rect 62502 42242 62508 42414
rect 62542 42242 62548 42414
rect 62502 42230 62548 42242
rect 63160 42414 63206 42426
rect 63160 42242 63166 42414
rect 63200 42242 63206 42414
rect 63160 42230 63206 42242
rect 63818 42414 63864 42426
rect 63818 42242 63824 42414
rect 63858 42242 63864 42414
rect 63818 42230 63864 42242
rect 64476 42414 64522 42426
rect 64476 42242 64482 42414
rect 64516 42242 64522 42414
rect 64476 42230 64522 42242
rect 65134 42414 65180 42426
rect 65134 42242 65140 42414
rect 65174 42242 65180 42414
rect 65134 42230 65180 42242
rect 65792 42414 65838 42426
rect 65792 42242 65798 42414
rect 65832 42242 65838 42414
rect 65792 42230 65838 42242
rect 62502 41720 62548 41732
rect 62502 41548 62508 41720
rect 62542 41548 62548 41720
rect 62502 41536 62548 41548
rect 63160 41720 63206 41732
rect 63160 41548 63166 41720
rect 63200 41548 63206 41720
rect 63160 41536 63206 41548
rect 63818 41720 63864 41732
rect 63818 41548 63824 41720
rect 63858 41548 63864 41720
rect 63818 41536 63864 41548
rect 64476 41720 64522 41732
rect 64476 41548 64482 41720
rect 64516 41548 64522 41720
rect 64476 41536 64522 41548
rect 65134 41720 65180 41732
rect 65134 41548 65140 41720
rect 65174 41548 65180 41720
rect 65134 41536 65180 41548
rect 65792 41720 65838 41732
rect 65792 41548 65798 41720
rect 65832 41548 65838 41720
rect 65792 41536 65838 41548
rect 62116 40790 62360 41028
rect 62502 41026 62548 41038
rect 62502 40854 62508 41026
rect 62542 40854 62548 41026
rect 62502 40842 62548 40854
rect 63160 41026 63206 41038
rect 63160 40854 63166 41026
rect 63200 40854 63206 41026
rect 63160 40842 63206 40854
rect 63818 41026 63864 41038
rect 63818 40854 63824 41026
rect 63858 40854 63864 41026
rect 63818 40842 63864 40854
rect 64476 41026 64522 41038
rect 64476 40854 64482 41026
rect 64516 40854 64522 41026
rect 64476 40842 64522 40854
rect 65134 41026 65180 41038
rect 65134 40854 65140 41026
rect 65174 40854 65180 41026
rect 65134 40842 65180 40854
rect 65792 41026 65838 41038
rect 65792 40854 65798 41026
rect 65832 40854 65838 41026
rect 65792 40842 65838 40854
rect 65942 41030 65988 42534
rect 66082 42408 66154 42534
rect 69750 42548 69962 42716
rect 69750 42468 69796 42548
rect 66296 42416 66342 42428
rect 66082 41030 66228 42408
rect 66296 42244 66302 42416
rect 66336 42244 66342 42416
rect 66296 42232 66342 42244
rect 66954 42416 67000 42428
rect 66954 42244 66960 42416
rect 66994 42244 67000 42416
rect 66954 42232 67000 42244
rect 67612 42416 67658 42428
rect 67612 42244 67618 42416
rect 67652 42244 67658 42416
rect 67612 42232 67658 42244
rect 68270 42416 68316 42428
rect 68270 42244 68276 42416
rect 68310 42244 68316 42416
rect 68270 42232 68316 42244
rect 68928 42416 68974 42428
rect 68928 42244 68934 42416
rect 68968 42244 68974 42416
rect 68928 42232 68974 42244
rect 69586 42416 69632 42428
rect 69586 42244 69592 42416
rect 69626 42244 69632 42416
rect 69586 42232 69632 42244
rect 66296 41722 66342 41734
rect 66296 41550 66302 41722
rect 66336 41550 66342 41722
rect 66296 41538 66342 41550
rect 66954 41722 67000 41734
rect 66954 41550 66960 41722
rect 66994 41550 67000 41722
rect 66954 41538 67000 41550
rect 67612 41722 67658 41734
rect 67612 41550 67618 41722
rect 67652 41550 67658 41722
rect 67612 41538 67658 41550
rect 68270 41722 68316 41734
rect 68270 41550 68276 41722
rect 68310 41550 68316 41722
rect 68270 41538 68316 41550
rect 68928 41722 68974 41734
rect 68928 41550 68934 41722
rect 68968 41550 68974 41722
rect 68928 41538 68974 41550
rect 69586 41722 69632 41734
rect 69586 41550 69592 41722
rect 69626 41550 69632 41722
rect 69586 41538 69632 41550
rect 69708 41044 69796 42468
rect 69890 42468 69962 42548
rect 73610 42542 73646 42876
rect 69890 41044 69984 42468
rect 70104 42430 70150 42442
rect 70104 42258 70110 42430
rect 70144 42258 70150 42430
rect 70104 42246 70150 42258
rect 70762 42430 70808 42442
rect 70762 42258 70768 42430
rect 70802 42258 70808 42430
rect 70762 42246 70808 42258
rect 71420 42430 71466 42442
rect 71420 42258 71426 42430
rect 71460 42258 71466 42430
rect 71420 42246 71466 42258
rect 72078 42430 72124 42442
rect 72078 42258 72084 42430
rect 72118 42258 72124 42430
rect 72078 42246 72124 42258
rect 72736 42430 72782 42442
rect 72736 42258 72742 42430
rect 72776 42258 72782 42430
rect 72736 42246 72782 42258
rect 73394 42430 73440 42442
rect 73394 42258 73400 42430
rect 73434 42258 73440 42430
rect 73394 42246 73440 42258
rect 70104 41736 70150 41748
rect 70104 41564 70110 41736
rect 70144 41564 70150 41736
rect 70104 41552 70150 41564
rect 70762 41736 70808 41748
rect 70762 41564 70768 41736
rect 70802 41564 70808 41736
rect 70762 41552 70808 41564
rect 71420 41736 71466 41748
rect 71420 41564 71426 41736
rect 71460 41564 71466 41736
rect 71420 41552 71466 41564
rect 72078 41736 72124 41748
rect 72078 41564 72084 41736
rect 72118 41564 72124 41736
rect 72078 41552 72124 41564
rect 72736 41736 72782 41748
rect 72736 41564 72742 41736
rect 72776 41564 72782 41736
rect 72736 41552 72782 41564
rect 73394 41736 73440 41748
rect 73394 41564 73400 41736
rect 73434 41564 73440 41736
rect 73394 41552 73440 41564
rect 65942 40792 66228 41030
rect 66296 41028 66342 41040
rect 66296 40856 66302 41028
rect 66336 40856 66342 41028
rect 66296 40844 66342 40856
rect 66954 41028 67000 41040
rect 66954 40856 66960 41028
rect 66994 40856 67000 41028
rect 66954 40844 67000 40856
rect 67612 41028 67658 41040
rect 67612 40856 67618 41028
rect 67652 40856 67658 41028
rect 67612 40844 67658 40856
rect 68270 41028 68316 41040
rect 68270 40856 68276 41028
rect 68310 40856 68316 41028
rect 68270 40844 68316 40856
rect 68928 41028 68974 41040
rect 68928 40856 68934 41028
rect 68968 40856 68974 41028
rect 68928 40844 68974 40856
rect 69586 41028 69632 41040
rect 69586 40856 69592 41028
rect 69626 40856 69632 41028
rect 69586 40844 69632 40856
rect 62116 39622 62296 40790
rect 62502 40332 62548 40344
rect 62502 40160 62508 40332
rect 62542 40160 62548 40332
rect 62502 40148 62548 40160
rect 63160 40332 63206 40344
rect 63160 40160 63166 40332
rect 63200 40160 63206 40332
rect 63160 40148 63206 40160
rect 63818 40332 63864 40344
rect 63818 40160 63824 40332
rect 63858 40160 63864 40332
rect 63818 40148 63864 40160
rect 64476 40332 64522 40344
rect 64476 40160 64482 40332
rect 64516 40160 64522 40332
rect 64476 40148 64522 40160
rect 65134 40332 65180 40344
rect 65134 40160 65140 40332
rect 65174 40160 65180 40332
rect 65134 40148 65180 40160
rect 65792 40332 65838 40344
rect 65792 40160 65798 40332
rect 65832 40160 65838 40332
rect 65792 40148 65838 40160
rect 65952 39622 66228 40792
rect 66296 40334 66342 40346
rect 66296 40162 66302 40334
rect 66336 40162 66342 40334
rect 66296 40150 66342 40162
rect 66954 40334 67000 40346
rect 66954 40162 66960 40334
rect 66994 40162 67000 40334
rect 66954 40150 67000 40162
rect 67612 40334 67658 40346
rect 67612 40162 67618 40334
rect 67652 40162 67658 40334
rect 67612 40150 67658 40162
rect 68270 40334 68316 40346
rect 68270 40162 68276 40334
rect 68310 40162 68316 40334
rect 68270 40150 68316 40162
rect 68928 40334 68974 40346
rect 68928 40162 68934 40334
rect 68968 40162 68974 40334
rect 68928 40150 68974 40162
rect 69586 40334 69632 40346
rect 69586 40162 69592 40334
rect 69626 40162 69632 40334
rect 69586 40150 69632 40162
rect 69708 39622 69984 41044
rect 70104 41042 70150 41054
rect 70104 40870 70110 41042
rect 70144 40870 70150 41042
rect 70104 40858 70150 40870
rect 70762 41042 70808 41054
rect 70762 40870 70768 41042
rect 70802 40870 70808 41042
rect 70762 40858 70808 40870
rect 71420 41042 71466 41054
rect 71420 40870 71426 41042
rect 71460 40870 71466 41042
rect 71420 40858 71466 40870
rect 72078 41042 72124 41054
rect 72078 40870 72084 41042
rect 72118 40870 72124 41042
rect 72078 40858 72124 40870
rect 72736 41042 72782 41054
rect 72736 40870 72742 41042
rect 72776 40870 72782 41042
rect 72736 40858 72782 40870
rect 73394 41042 73440 41054
rect 73394 40870 73400 41042
rect 73434 40870 73440 41042
rect 73394 40858 73440 40870
rect 73598 40970 73646 42542
rect 73876 40970 73950 42876
rect 79424 41422 79538 43084
rect 80598 41576 80954 46204
rect 88542 42666 88552 43684
rect 89804 42666 89814 43684
rect 79422 41196 80188 41422
rect 73598 40668 73950 40970
rect 70104 40348 70150 40360
rect 70104 40176 70110 40348
rect 70144 40176 70150 40348
rect 70104 40164 70150 40176
rect 70762 40348 70808 40360
rect 70762 40176 70768 40348
rect 70802 40176 70808 40348
rect 70762 40164 70808 40176
rect 71420 40348 71466 40360
rect 71420 40176 71426 40348
rect 71460 40176 71466 40348
rect 71420 40164 71466 40176
rect 72078 40348 72124 40360
rect 72078 40176 72084 40348
rect 72118 40176 72124 40348
rect 72078 40164 72124 40176
rect 72736 40348 72782 40360
rect 72736 40176 72742 40348
rect 72776 40176 72782 40348
rect 72736 40164 72782 40176
rect 73394 40348 73440 40360
rect 73394 40176 73400 40348
rect 73434 40176 73440 40348
rect 73394 40164 73440 40176
rect 73598 39634 73874 40668
rect 76654 39634 76954 39646
rect 73508 39622 76954 39634
rect 62116 39454 76954 39622
rect 62140 39418 73870 39454
rect 65952 39370 66228 39418
rect 76654 39082 76954 39454
rect 78496 39506 78834 39528
rect 78496 39416 78570 39506
rect 78774 39416 78834 39506
rect 78496 39386 78834 39416
rect 80106 39474 80188 41196
rect 80598 39582 80952 41576
rect 86688 40886 87154 40908
rect 88846 40886 89414 42666
rect 86626 40396 89414 40886
rect 80598 39522 81140 39582
rect 80106 39470 80530 39474
rect 80598 39470 80908 39522
rect 80106 39410 80534 39470
rect 77164 39094 77210 39106
rect 59376 35896 59422 35908
rect 40984 35070 41030 35082
rect 40984 34778 40990 35070
rect 41024 34778 41030 35070
rect 40984 34766 41030 34778
rect 42042 35070 42088 35082
rect 42042 34778 42048 35070
rect 42082 34778 42088 35070
rect 42042 34766 42088 34778
rect 43100 35070 43146 35082
rect 43100 34778 43106 35070
rect 43140 34778 43146 35070
rect 43100 34766 43146 34778
rect 44158 35070 44204 35082
rect 44158 34778 44164 35070
rect 44198 34778 44204 35070
rect 44158 34766 44204 34778
rect 45216 35070 45262 35082
rect 45216 34778 45222 35070
rect 45256 34778 45262 35070
rect 45216 34766 45262 34778
rect 46274 35070 46320 35082
rect 46274 34778 46280 35070
rect 46314 34778 46320 35070
rect 46274 34766 46320 34778
rect 34494 33976 34540 33988
rect 34494 33684 34500 33976
rect 34534 33684 34540 33976
rect 34494 33672 34540 33684
rect 35552 33976 35598 33988
rect 35552 33684 35558 33976
rect 35592 33684 35598 33976
rect 35552 33672 35598 33684
rect 36610 33976 36656 33988
rect 36610 33684 36616 33976
rect 36650 33684 36656 33976
rect 36610 33672 36656 33684
rect 37668 33976 37714 33988
rect 37668 33684 37674 33976
rect 37708 33684 37714 33976
rect 37668 33672 37714 33684
rect 38726 33976 38772 33988
rect 38726 33684 38732 33976
rect 38766 33684 38772 33976
rect 38726 33672 38772 33684
rect 39784 33976 39830 33988
rect 39784 33684 39790 33976
rect 39824 33684 39830 33976
rect 39784 33672 39830 33684
rect 34494 32882 34540 32894
rect 34494 32590 34500 32882
rect 34534 32590 34540 32882
rect 34494 32578 34540 32590
rect 35552 32882 35598 32894
rect 35552 32590 35558 32882
rect 35592 32590 35598 32882
rect 35552 32578 35598 32590
rect 36610 32882 36656 32894
rect 36610 32590 36616 32882
rect 36650 32590 36656 32882
rect 36610 32578 36656 32590
rect 37668 32882 37714 32894
rect 37668 32590 37674 32882
rect 37708 32590 37714 32882
rect 37668 32578 37714 32590
rect 38726 32882 38772 32894
rect 38726 32590 38732 32882
rect 38766 32590 38772 32882
rect 38726 32578 38772 32590
rect 39784 32882 39830 32894
rect 39784 32590 39790 32882
rect 39824 32590 39830 32882
rect 39784 32578 39830 32590
rect 34494 31424 34540 31436
rect 34494 31132 34500 31424
rect 34534 31132 34540 31424
rect 34494 31120 34540 31132
rect 35552 31424 35598 31436
rect 35552 31132 35558 31424
rect 35592 31132 35598 31424
rect 35552 31120 35598 31132
rect 36610 31424 36656 31436
rect 36610 31132 36616 31424
rect 36650 31132 36656 31424
rect 36610 31120 36656 31132
rect 37668 31424 37714 31436
rect 37668 31132 37674 31424
rect 37708 31132 37714 31424
rect 37668 31120 37714 31132
rect 38726 31424 38772 31436
rect 38726 31132 38732 31424
rect 38766 31132 38772 31424
rect 38726 31120 38772 31132
rect 39784 31424 39830 31436
rect 39784 31132 39790 31424
rect 39824 31132 39830 31424
rect 39784 31120 39830 31132
rect 34494 30330 34540 30342
rect 34494 30038 34500 30330
rect 34534 30038 34540 30330
rect 34494 30026 34540 30038
rect 35552 30330 35598 30342
rect 35552 30038 35558 30330
rect 35592 30038 35598 30330
rect 35552 30026 35598 30038
rect 36610 30330 36656 30342
rect 36610 30038 36616 30330
rect 36650 30038 36656 30330
rect 36610 30026 36656 30038
rect 37668 30330 37714 30342
rect 37668 30038 37674 30330
rect 37708 30038 37714 30330
rect 37668 30026 37714 30038
rect 38726 30330 38772 30342
rect 38726 30038 38732 30330
rect 38766 30038 38772 30330
rect 38726 30026 38772 30038
rect 39784 30330 39830 30342
rect 39784 30038 39790 30330
rect 39824 30038 39830 30330
rect 39784 30026 39830 30038
rect 21462 29214 21508 29226
rect 21462 28922 21468 29214
rect 21502 28922 21508 29214
rect 21462 28910 21508 28922
rect 22520 29214 22566 29226
rect 22520 28922 22526 29214
rect 22560 28922 22566 29214
rect 22520 28910 22566 28922
rect 23578 29214 23624 29226
rect 23578 28922 23584 29214
rect 23618 28922 23624 29214
rect 23578 28910 23624 28922
rect 24636 29214 24682 29226
rect 24636 28922 24642 29214
rect 24676 28922 24682 29214
rect 24636 28910 24682 28922
rect 25694 29214 25740 29226
rect 25694 28922 25700 29214
rect 25734 28922 25740 29214
rect 25694 28910 25740 28922
rect 26752 29214 26798 29226
rect 26752 28922 26758 29214
rect 26792 28922 26798 29214
rect 26752 28910 26798 28922
rect 14972 28136 15018 28148
rect 14972 27844 14978 28136
rect 15012 27844 15018 28136
rect 14972 27832 15018 27844
rect 16030 28136 16076 28148
rect 16030 27844 16036 28136
rect 16070 27844 16076 28136
rect 16030 27832 16076 27844
rect 17088 28136 17134 28148
rect 17088 27844 17094 28136
rect 17128 27844 17134 28136
rect 17088 27832 17134 27844
rect 18146 28136 18192 28148
rect 18146 27844 18152 28136
rect 18186 27844 18192 28136
rect 18146 27832 18192 27844
rect 19204 28136 19250 28148
rect 19204 27844 19210 28136
rect 19244 27844 19250 28136
rect 19204 27832 19250 27844
rect 20262 28136 20308 28148
rect 20262 27844 20268 28136
rect 20302 27844 20308 28136
rect 20262 27832 20308 27844
rect 14972 27042 15018 27054
rect 14972 26750 14978 27042
rect 15012 26750 15018 27042
rect 14972 26738 15018 26750
rect 16030 27042 16076 27054
rect 16030 26750 16036 27042
rect 16070 26750 16076 27042
rect 16030 26738 16076 26750
rect 17088 27042 17134 27054
rect 17088 26750 17094 27042
rect 17128 26750 17134 27042
rect 17088 26738 17134 26750
rect 18146 27042 18192 27054
rect 18146 26750 18152 27042
rect 18186 26750 18192 27042
rect 18146 26738 18192 26750
rect 19204 27042 19250 27054
rect 19204 26750 19210 27042
rect 19244 26750 19250 27042
rect 19204 26738 19250 26750
rect 20262 27042 20308 27054
rect 20262 26750 20268 27042
rect 20302 26750 20308 27042
rect 20262 26738 20308 26750
rect 14972 25582 15018 25594
rect 14972 25290 14978 25582
rect 15012 25290 15018 25582
rect 14972 25278 15018 25290
rect 16030 25582 16076 25594
rect 16030 25290 16036 25582
rect 16070 25290 16076 25582
rect 16030 25278 16076 25290
rect 17088 25582 17134 25594
rect 17088 25290 17094 25582
rect 17128 25290 17134 25582
rect 17088 25278 17134 25290
rect 18146 25582 18192 25594
rect 18146 25290 18152 25582
rect 18186 25290 18192 25582
rect 18146 25278 18192 25290
rect 19204 25582 19250 25594
rect 19204 25290 19210 25582
rect 19244 25290 19250 25582
rect 19204 25278 19250 25290
rect 20262 25582 20308 25594
rect 20262 25290 20268 25582
rect 20302 25290 20308 25582
rect 20262 25278 20308 25290
rect 14972 24488 15018 24500
rect 14972 24196 14978 24488
rect 15012 24196 15018 24488
rect 14972 24184 15018 24196
rect 16030 24488 16076 24500
rect 16030 24196 16036 24488
rect 16070 24196 16076 24488
rect 16030 24184 16076 24196
rect 17088 24488 17134 24500
rect 17088 24196 17094 24488
rect 17128 24196 17134 24488
rect 17088 24184 17134 24196
rect 18146 24488 18192 24500
rect 18146 24196 18152 24488
rect 18186 24196 18192 24488
rect 18146 24184 18192 24196
rect 19204 24488 19250 24500
rect 19204 24196 19210 24488
rect 19244 24196 19250 24488
rect 19204 24184 19250 24196
rect 20262 24488 20308 24500
rect 20262 24196 20268 24488
rect 20302 24196 20308 24488
rect 20262 24184 20308 24196
rect 8466 23386 8512 23398
rect 8466 23094 8472 23386
rect 8506 23094 8512 23386
rect 8466 23082 8512 23094
rect 9524 23386 9570 23398
rect 9524 23094 9530 23386
rect 9564 23094 9570 23386
rect 9524 23082 9570 23094
rect 10582 23386 10628 23398
rect 10582 23094 10588 23386
rect 10622 23094 10628 23386
rect 10582 23082 10628 23094
rect 11640 23386 11686 23398
rect 11640 23094 11646 23386
rect 11680 23094 11686 23386
rect 11640 23082 11686 23094
rect 12698 23386 12744 23398
rect 12698 23094 12704 23386
rect 12738 23094 12744 23386
rect 12698 23082 12744 23094
rect 13756 23386 13802 23398
rect 13756 23094 13762 23386
rect 13796 23094 13802 23386
rect 13756 23082 13802 23094
rect 1952 22284 1998 22296
rect 1952 21992 1958 22284
rect 1992 21992 1998 22284
rect 1952 21980 1998 21992
rect 3010 22284 3056 22296
rect 3010 21992 3016 22284
rect 3050 21992 3056 22284
rect 3010 21980 3056 21992
rect 4068 22284 4114 22296
rect 4068 21992 4074 22284
rect 4108 21992 4114 22284
rect 4068 21980 4114 21992
rect 5126 22284 5172 22296
rect 5126 21992 5132 22284
rect 5166 21992 5172 22284
rect 5126 21980 5172 21992
rect 6184 22284 6230 22296
rect 6184 21992 6190 22284
rect 6224 21992 6230 22284
rect 6184 21980 6230 21992
rect 7242 22284 7288 22296
rect 7242 21992 7248 22284
rect 7282 21992 7288 22284
rect 7242 21980 7288 21992
rect 1952 21190 1998 21202
rect 1952 20898 1958 21190
rect 1992 20898 1998 21190
rect 1952 20886 1998 20898
rect 3010 21190 3056 21202
rect 3010 20898 3016 21190
rect 3050 20898 3056 21190
rect 3010 20886 3056 20898
rect 4068 21190 4114 21202
rect 4068 20898 4074 21190
rect 4108 20898 4114 21190
rect 4068 20886 4114 20898
rect 5126 21190 5172 21202
rect 5126 20898 5132 21190
rect 5166 20898 5172 21190
rect 5126 20886 5172 20898
rect 6184 21190 6230 21202
rect 6184 20898 6190 21190
rect 6224 20898 6230 21190
rect 6184 20886 6230 20898
rect 7242 21190 7288 21202
rect 7242 20898 7248 21190
rect 7282 20898 7288 21190
rect 7242 20886 7288 20898
rect 1952 19702 1998 19714
rect 1952 19410 1958 19702
rect 1992 19410 1998 19702
rect 1952 19398 1998 19410
rect 3010 19702 3056 19714
rect 3010 19410 3016 19702
rect 3050 19410 3056 19702
rect 3010 19398 3056 19410
rect 4068 19702 4114 19714
rect 4068 19410 4074 19702
rect 4108 19410 4114 19702
rect 4068 19398 4114 19410
rect 5126 19702 5172 19714
rect 5126 19410 5132 19702
rect 5166 19410 5172 19702
rect 5126 19398 5172 19410
rect 6184 19702 6230 19714
rect 6184 19410 6190 19702
rect 6224 19410 6230 19702
rect 6184 19398 6230 19410
rect 7242 19702 7288 19714
rect 7242 19410 7248 19702
rect 7282 19410 7288 19702
rect 7242 19398 7288 19410
rect 1952 18608 1998 18620
rect 1952 18316 1958 18608
rect 1992 18316 1998 18608
rect 1952 18304 1998 18316
rect 3010 18608 3056 18620
rect 3010 18316 3016 18608
rect 3050 18316 3056 18608
rect 3010 18304 3056 18316
rect 4068 18608 4114 18620
rect 4068 18316 4074 18608
rect 4108 18316 4114 18608
rect 4068 18304 4114 18316
rect 5126 18608 5172 18620
rect 5126 18316 5132 18608
rect 5166 18316 5172 18608
rect 5126 18304 5172 18316
rect 6184 18608 6230 18620
rect 6184 18316 6190 18608
rect 6224 18316 6230 18608
rect 6184 18304 6230 18316
rect 7242 18608 7288 18620
rect 7242 18316 7248 18608
rect 7282 18316 7288 18608
rect 7242 18304 7288 18316
rect 1264 16972 1326 18168
rect 1420 16972 1560 18168
rect 7722 18176 8018 22844
rect 14216 22852 14346 24048
rect 14440 22852 14512 24048
rect 20748 24032 21044 28672
rect 27278 28688 27358 29884
rect 27452 28688 27574 29884
rect 33846 29890 34144 30016
rect 27984 29230 28030 29242
rect 27984 28938 27990 29230
rect 28024 28938 28030 29230
rect 27984 28926 28030 28938
rect 29042 29230 29088 29242
rect 29042 28938 29048 29230
rect 29082 28938 29088 29230
rect 29042 28926 29088 28938
rect 30100 29230 30146 29242
rect 30100 28938 30106 29230
rect 30140 28938 30146 29230
rect 30100 28926 30146 28938
rect 31158 29230 31204 29242
rect 31158 28938 31164 29230
rect 31198 28938 31204 29230
rect 31158 28926 31204 28938
rect 32216 29230 32262 29242
rect 32216 28938 32222 29230
rect 32256 28938 32262 29230
rect 32216 28926 32262 28938
rect 33274 29230 33320 29242
rect 33274 28938 33280 29230
rect 33314 28938 33320 29230
rect 33274 28926 33320 28938
rect 21462 28120 21508 28132
rect 21462 27828 21468 28120
rect 21502 27828 21508 28120
rect 21462 27816 21508 27828
rect 22520 28120 22566 28132
rect 22520 27828 22526 28120
rect 22560 27828 22566 28120
rect 22520 27816 22566 27828
rect 23578 28120 23624 28132
rect 23578 27828 23584 28120
rect 23618 27828 23624 28120
rect 23578 27816 23624 27828
rect 24636 28120 24682 28132
rect 24636 27828 24642 28120
rect 24676 27828 24682 28120
rect 24636 27816 24682 27828
rect 25694 28120 25740 28132
rect 25694 27828 25700 28120
rect 25734 27828 25740 28120
rect 25694 27816 25740 27828
rect 26752 28120 26798 28132
rect 26752 27828 26758 28120
rect 26792 27828 26798 28120
rect 26752 27816 26798 27828
rect 21462 27026 21508 27038
rect 21462 26734 21468 27026
rect 21502 26734 21508 27026
rect 21462 26722 21508 26734
rect 22520 27026 22566 27038
rect 22520 26734 22526 27026
rect 22560 26734 22566 27026
rect 22520 26722 22566 26734
rect 23578 27026 23624 27038
rect 23578 26734 23584 27026
rect 23618 26734 23624 27026
rect 23578 26722 23624 26734
rect 24636 27026 24682 27038
rect 24636 26734 24642 27026
rect 24676 26734 24682 27026
rect 24636 26722 24682 26734
rect 25694 27026 25740 27038
rect 25694 26734 25700 27026
rect 25734 26734 25740 27026
rect 25694 26722 25740 26734
rect 26752 27026 26798 27038
rect 26752 26734 26758 27026
rect 26792 26734 26798 27026
rect 26752 26722 26798 26734
rect 21462 25566 21508 25578
rect 21462 25274 21468 25566
rect 21502 25274 21508 25566
rect 21462 25262 21508 25274
rect 22520 25566 22566 25578
rect 22520 25274 22526 25566
rect 22560 25274 22566 25566
rect 22520 25262 22566 25274
rect 23578 25566 23624 25578
rect 23578 25274 23584 25566
rect 23618 25274 23624 25566
rect 23578 25262 23624 25274
rect 24636 25566 24682 25578
rect 24636 25274 24642 25566
rect 24676 25274 24682 25566
rect 24636 25262 24682 25274
rect 25694 25566 25740 25578
rect 25694 25274 25700 25566
rect 25734 25274 25740 25566
rect 25694 25262 25740 25274
rect 26752 25566 26798 25578
rect 26752 25274 26758 25566
rect 26792 25274 26798 25566
rect 26752 25262 26798 25274
rect 21462 24472 21508 24484
rect 21462 24180 21468 24472
rect 21502 24180 21508 24472
rect 21462 24168 21508 24180
rect 22520 24472 22566 24484
rect 22520 24180 22526 24472
rect 22560 24180 22566 24472
rect 22520 24168 22566 24180
rect 23578 24472 23624 24484
rect 23578 24180 23584 24472
rect 23618 24180 23624 24472
rect 23578 24168 23624 24180
rect 24636 24472 24682 24484
rect 24636 24180 24642 24472
rect 24676 24180 24682 24472
rect 24636 24168 24682 24180
rect 25694 24472 25740 24484
rect 25694 24180 25700 24472
rect 25734 24180 25740 24472
rect 25694 24168 25740 24180
rect 26752 24472 26798 24484
rect 26752 24180 26758 24472
rect 26792 24180 26798 24472
rect 26752 24168 26798 24180
rect 14972 23394 15018 23406
rect 14972 23102 14978 23394
rect 15012 23102 15018 23394
rect 14972 23090 15018 23102
rect 16030 23394 16076 23406
rect 16030 23102 16036 23394
rect 16070 23102 16076 23394
rect 16030 23090 16076 23102
rect 17088 23394 17134 23406
rect 17088 23102 17094 23394
rect 17128 23102 17134 23394
rect 17088 23090 17134 23102
rect 18146 23394 18192 23406
rect 18146 23102 18152 23394
rect 18186 23102 18192 23394
rect 18146 23090 18192 23102
rect 19204 23394 19250 23406
rect 19204 23102 19210 23394
rect 19244 23102 19250 23394
rect 19204 23090 19250 23102
rect 20262 23394 20308 23406
rect 20262 23102 20268 23394
rect 20302 23102 20308 23394
rect 20262 23090 20308 23102
rect 8466 22292 8512 22304
rect 8466 22000 8472 22292
rect 8506 22000 8512 22292
rect 8466 21988 8512 22000
rect 9524 22292 9570 22304
rect 9524 22000 9530 22292
rect 9564 22000 9570 22292
rect 9524 21988 9570 22000
rect 10582 22292 10628 22304
rect 10582 22000 10588 22292
rect 10622 22000 10628 22292
rect 10582 21988 10628 22000
rect 11640 22292 11686 22304
rect 11640 22000 11646 22292
rect 11680 22000 11686 22292
rect 11640 21988 11686 22000
rect 12698 22292 12744 22304
rect 12698 22000 12704 22292
rect 12738 22000 12744 22292
rect 12698 21988 12744 22000
rect 13756 22292 13802 22304
rect 13756 22000 13762 22292
rect 13796 22000 13802 22292
rect 13756 21988 13802 22000
rect 8466 21198 8512 21210
rect 8466 20906 8472 21198
rect 8506 20906 8512 21198
rect 8466 20894 8512 20906
rect 9524 21198 9570 21210
rect 9524 20906 9530 21198
rect 9564 20906 9570 21198
rect 9524 20894 9570 20906
rect 10582 21198 10628 21210
rect 10582 20906 10588 21198
rect 10622 20906 10628 21198
rect 10582 20894 10628 20906
rect 11640 21198 11686 21210
rect 11640 20906 11646 21198
rect 11680 20906 11686 21198
rect 11640 20894 11686 20906
rect 12698 21198 12744 21210
rect 12698 20906 12704 21198
rect 12738 20906 12744 21198
rect 12698 20894 12744 20906
rect 13756 21198 13802 21210
rect 13756 20906 13762 21198
rect 13796 20906 13802 21198
rect 13756 20894 13802 20906
rect 8466 19710 8512 19722
rect 8466 19418 8472 19710
rect 8506 19418 8512 19710
rect 8466 19406 8512 19418
rect 9524 19710 9570 19722
rect 9524 19418 9530 19710
rect 9564 19418 9570 19710
rect 9524 19406 9570 19418
rect 10582 19710 10628 19722
rect 10582 19418 10588 19710
rect 10622 19418 10628 19710
rect 10582 19406 10628 19418
rect 11640 19710 11686 19722
rect 11640 19418 11646 19710
rect 11680 19418 11686 19710
rect 11640 19406 11686 19418
rect 12698 19710 12744 19722
rect 12698 19418 12704 19710
rect 12738 19418 12744 19710
rect 12698 19406 12744 19418
rect 13756 19710 13802 19722
rect 13756 19418 13762 19710
rect 13796 19418 13802 19710
rect 13756 19406 13802 19418
rect 8466 18616 8512 18628
rect 8466 18324 8472 18616
rect 8506 18324 8512 18616
rect 8466 18312 8512 18324
rect 9524 18616 9570 18628
rect 9524 18324 9530 18616
rect 9564 18324 9570 18616
rect 9524 18312 9570 18324
rect 10582 18616 10628 18628
rect 10582 18324 10588 18616
rect 10622 18324 10628 18616
rect 10582 18312 10628 18324
rect 11640 18616 11686 18628
rect 11640 18324 11646 18616
rect 11680 18324 11686 18616
rect 11640 18312 11686 18324
rect 12698 18616 12744 18628
rect 12698 18324 12704 18616
rect 12738 18324 12744 18616
rect 12698 18312 12744 18324
rect 13756 18616 13802 18628
rect 13756 18324 13762 18616
rect 13796 18324 13802 18616
rect 13756 18312 13802 18324
rect 1952 17514 1998 17526
rect 1952 17222 1958 17514
rect 1992 17222 1998 17514
rect 1952 17210 1998 17222
rect 3010 17514 3056 17526
rect 3010 17222 3016 17514
rect 3050 17222 3056 17514
rect 3010 17210 3056 17222
rect 4068 17514 4114 17526
rect 4068 17222 4074 17514
rect 4108 17222 4114 17514
rect 4068 17210 4114 17222
rect 5126 17514 5172 17526
rect 5126 17222 5132 17514
rect 5166 17222 5172 17514
rect 5126 17210 5172 17222
rect 6184 17514 6230 17526
rect 6184 17222 6190 17514
rect 6224 17222 6230 17514
rect 6184 17210 6230 17222
rect 7242 17514 7288 17526
rect 7242 17222 7248 17514
rect 7282 17222 7288 17514
rect 7242 17210 7288 17222
rect 1264 12312 1560 16972
rect 7722 16980 7840 18176
rect 7934 16980 8018 18176
rect 14216 18184 14512 22852
rect 20748 22836 20836 24032
rect 20930 22836 21044 24032
rect 27278 24048 27574 28688
rect 33846 28694 33868 29890
rect 33962 28694 34144 29890
rect 40304 29890 40638 34528
rect 46836 34550 46946 35746
rect 47040 34550 47170 35746
rect 53438 35760 53776 35886
rect 47572 35092 47618 35104
rect 47572 34800 47578 35092
rect 47612 34800 47618 35092
rect 47572 34788 47618 34800
rect 48630 35092 48676 35104
rect 48630 34800 48636 35092
rect 48670 34800 48676 35092
rect 48630 34788 48676 34800
rect 49688 35092 49734 35104
rect 49688 34800 49694 35092
rect 49728 34800 49734 35092
rect 49688 34788 49734 34800
rect 50746 35092 50792 35104
rect 50746 34800 50752 35092
rect 50786 34800 50792 35092
rect 50746 34788 50792 34800
rect 51804 35092 51850 35104
rect 51804 34800 51810 35092
rect 51844 34800 51850 35092
rect 51804 34788 51850 34800
rect 52862 35092 52908 35104
rect 52862 34800 52868 35092
rect 52902 34800 52908 35092
rect 52862 34788 52908 34800
rect 40984 33976 41030 33988
rect 40984 33684 40990 33976
rect 41024 33684 41030 33976
rect 40984 33672 41030 33684
rect 42042 33976 42088 33988
rect 42042 33684 42048 33976
rect 42082 33684 42088 33976
rect 42042 33672 42088 33684
rect 43100 33976 43146 33988
rect 43100 33684 43106 33976
rect 43140 33684 43146 33976
rect 43100 33672 43146 33684
rect 44158 33976 44204 33988
rect 44158 33684 44164 33976
rect 44198 33684 44204 33976
rect 44158 33672 44204 33684
rect 45216 33976 45262 33988
rect 45216 33684 45222 33976
rect 45256 33684 45262 33976
rect 45216 33672 45262 33684
rect 46274 33976 46320 33988
rect 46274 33684 46280 33976
rect 46314 33684 46320 33976
rect 46274 33672 46320 33684
rect 40984 32882 41030 32894
rect 40984 32590 40990 32882
rect 41024 32590 41030 32882
rect 40984 32578 41030 32590
rect 42042 32882 42088 32894
rect 42042 32590 42048 32882
rect 42082 32590 42088 32882
rect 42042 32578 42088 32590
rect 43100 32882 43146 32894
rect 43100 32590 43106 32882
rect 43140 32590 43146 32882
rect 43100 32578 43146 32590
rect 44158 32882 44204 32894
rect 44158 32590 44164 32882
rect 44198 32590 44204 32882
rect 44158 32578 44204 32590
rect 45216 32882 45262 32894
rect 45216 32590 45222 32882
rect 45256 32590 45262 32882
rect 45216 32578 45262 32590
rect 46274 32882 46320 32894
rect 46274 32590 46280 32882
rect 46314 32590 46320 32882
rect 46274 32578 46320 32590
rect 40984 31424 41030 31436
rect 40984 31132 40990 31424
rect 41024 31132 41030 31424
rect 40984 31120 41030 31132
rect 42042 31424 42088 31436
rect 42042 31132 42048 31424
rect 42082 31132 42088 31424
rect 42042 31120 42088 31132
rect 43100 31424 43146 31436
rect 43100 31132 43106 31424
rect 43140 31132 43146 31424
rect 43100 31120 43146 31132
rect 44158 31424 44204 31436
rect 44158 31132 44164 31424
rect 44198 31132 44204 31424
rect 44158 31120 44204 31132
rect 45216 31424 45262 31436
rect 45216 31132 45222 31424
rect 45256 31132 45262 31424
rect 45216 31120 45262 31132
rect 46274 31424 46320 31436
rect 46274 31132 46280 31424
rect 46314 31132 46320 31424
rect 46274 31120 46320 31132
rect 40984 30330 41030 30342
rect 40984 30038 40990 30330
rect 41024 30038 41030 30330
rect 40984 30026 41030 30038
rect 42042 30330 42088 30342
rect 42042 30038 42048 30330
rect 42082 30038 42088 30330
rect 42042 30026 42088 30038
rect 43100 30330 43146 30342
rect 43100 30038 43106 30330
rect 43140 30038 43146 30330
rect 43100 30026 43146 30038
rect 44158 30330 44204 30342
rect 44158 30038 44164 30330
rect 44198 30038 44204 30330
rect 44158 30026 44204 30038
rect 45216 30330 45262 30342
rect 45216 30038 45222 30330
rect 45256 30038 45262 30330
rect 45216 30026 45262 30038
rect 46274 30330 46320 30342
rect 46274 30038 46280 30330
rect 46314 30038 46320 30330
rect 46274 30026 46320 30038
rect 34494 29236 34540 29248
rect 34494 28944 34500 29236
rect 34534 28944 34540 29236
rect 34494 28932 34540 28944
rect 35552 29236 35598 29248
rect 35552 28944 35558 29236
rect 35592 28944 35598 29236
rect 35552 28932 35598 28944
rect 36610 29236 36656 29248
rect 36610 28944 36616 29236
rect 36650 28944 36656 29236
rect 36610 28932 36656 28944
rect 37668 29236 37714 29248
rect 37668 28944 37674 29236
rect 37708 28944 37714 29236
rect 37668 28932 37714 28944
rect 38726 29236 38772 29248
rect 38726 28944 38732 29236
rect 38766 28944 38772 29236
rect 38726 28932 38772 28944
rect 39784 29236 39830 29248
rect 39784 28944 39790 29236
rect 39824 28944 39830 29236
rect 39784 28932 39830 28944
rect 33846 28370 34144 28694
rect 27984 28136 28030 28148
rect 27984 27844 27990 28136
rect 28024 27844 28030 28136
rect 27984 27832 28030 27844
rect 29042 28136 29088 28148
rect 29042 27844 29048 28136
rect 29082 27844 29088 28136
rect 29042 27832 29088 27844
rect 30100 28136 30146 28148
rect 30100 27844 30106 28136
rect 30140 27844 30146 28136
rect 30100 27832 30146 27844
rect 31158 28136 31204 28148
rect 31158 27844 31164 28136
rect 31198 27844 31204 28136
rect 31158 27832 31204 27844
rect 32216 28136 32262 28148
rect 32216 27844 32222 28136
rect 32256 27844 32262 28136
rect 32216 27832 32262 27844
rect 33274 28136 33320 28148
rect 33274 27844 33280 28136
rect 33314 27844 33320 28136
rect 33274 27832 33320 27844
rect 27984 27042 28030 27054
rect 27984 26750 27990 27042
rect 28024 26750 28030 27042
rect 27984 26738 28030 26750
rect 29042 27042 29088 27054
rect 29042 26750 29048 27042
rect 29082 26750 29088 27042
rect 29042 26738 29088 26750
rect 30100 27042 30146 27054
rect 30100 26750 30106 27042
rect 30140 26750 30146 27042
rect 30100 26738 30146 26750
rect 31158 27042 31204 27054
rect 31158 26750 31164 27042
rect 31198 26750 31204 27042
rect 31158 26738 31204 26750
rect 32216 27042 32262 27054
rect 32216 26750 32222 27042
rect 32256 26750 32262 27042
rect 32216 26738 32262 26750
rect 33274 27042 33320 27054
rect 33274 26750 33280 27042
rect 33314 26750 33320 27042
rect 33274 26738 33320 26750
rect 27984 25582 28030 25594
rect 27984 25290 27990 25582
rect 28024 25290 28030 25582
rect 27984 25278 28030 25290
rect 29042 25582 29088 25594
rect 29042 25290 29048 25582
rect 29082 25290 29088 25582
rect 29042 25278 29088 25290
rect 30100 25582 30146 25594
rect 30100 25290 30106 25582
rect 30140 25290 30146 25582
rect 30100 25278 30146 25290
rect 31158 25582 31204 25594
rect 31158 25290 31164 25582
rect 31198 25290 31204 25582
rect 31158 25278 31204 25290
rect 32216 25582 32262 25594
rect 32216 25290 32222 25582
rect 32256 25290 32262 25582
rect 32216 25278 32262 25290
rect 33274 25582 33320 25594
rect 33274 25290 33280 25582
rect 33314 25290 33320 25582
rect 33274 25278 33320 25290
rect 27984 24488 28030 24500
rect 27984 24196 27990 24488
rect 28024 24196 28030 24488
rect 27984 24184 28030 24196
rect 29042 24488 29088 24500
rect 29042 24196 29048 24488
rect 29082 24196 29088 24488
rect 29042 24184 29088 24196
rect 30100 24488 30146 24500
rect 30100 24196 30106 24488
rect 30140 24196 30146 24488
rect 30100 24184 30146 24196
rect 31158 24488 31204 24500
rect 31158 24196 31164 24488
rect 31198 24196 31204 24488
rect 31158 24184 31204 24196
rect 32216 24488 32262 24500
rect 32216 24196 32222 24488
rect 32256 24196 32262 24488
rect 32216 24184 32262 24196
rect 33274 24488 33320 24500
rect 33274 24196 33280 24488
rect 33314 24196 33320 24488
rect 33274 24184 33320 24196
rect 33848 24180 34144 28370
rect 40304 28694 40358 29890
rect 40452 28694 40638 29890
rect 46836 29912 47170 34550
rect 53438 34564 53460 35760
rect 53554 34564 53776 35760
rect 59600 35834 60012 36084
rect 54086 35106 54132 35118
rect 54086 34814 54092 35106
rect 54126 34814 54132 35106
rect 54086 34802 54132 34814
rect 55144 35106 55190 35118
rect 55144 34814 55150 35106
rect 55184 34814 55190 35106
rect 55144 34802 55190 34814
rect 56202 35106 56248 35118
rect 56202 34814 56208 35106
rect 56242 34814 56248 35106
rect 56202 34802 56248 34814
rect 57260 35106 57306 35118
rect 57260 34814 57266 35106
rect 57300 34814 57306 35106
rect 57260 34802 57306 34814
rect 58318 35106 58364 35118
rect 58318 34814 58324 35106
rect 58358 34814 58364 35106
rect 58318 34802 58364 34814
rect 59376 35106 59422 35118
rect 59376 34814 59382 35106
rect 59416 34814 59422 35106
rect 59376 34802 59422 34814
rect 53438 34240 53776 34564
rect 47572 33998 47618 34010
rect 47572 33706 47578 33998
rect 47612 33706 47618 33998
rect 47572 33694 47618 33706
rect 48630 33998 48676 34010
rect 48630 33706 48636 33998
rect 48670 33706 48676 33998
rect 48630 33694 48676 33706
rect 49688 33998 49734 34010
rect 49688 33706 49694 33998
rect 49728 33706 49734 33998
rect 49688 33694 49734 33706
rect 50746 33998 50792 34010
rect 50746 33706 50752 33998
rect 50786 33706 50792 33998
rect 50746 33694 50792 33706
rect 51804 33998 51850 34010
rect 51804 33706 51810 33998
rect 51844 33706 51850 33998
rect 51804 33694 51850 33706
rect 52862 33998 52908 34010
rect 52862 33706 52868 33998
rect 52902 33706 52908 33998
rect 52862 33694 52908 33706
rect 47572 32904 47618 32916
rect 47572 32612 47578 32904
rect 47612 32612 47618 32904
rect 47572 32600 47618 32612
rect 48630 32904 48676 32916
rect 48630 32612 48636 32904
rect 48670 32612 48676 32904
rect 48630 32600 48676 32612
rect 49688 32904 49734 32916
rect 49688 32612 49694 32904
rect 49728 32612 49734 32904
rect 49688 32600 49734 32612
rect 50746 32904 50792 32916
rect 50746 32612 50752 32904
rect 50786 32612 50792 32904
rect 50746 32600 50792 32612
rect 51804 32904 51850 32916
rect 51804 32612 51810 32904
rect 51844 32612 51850 32904
rect 51804 32600 51850 32612
rect 52862 32904 52908 32916
rect 52862 32612 52868 32904
rect 52902 32612 52908 32904
rect 52862 32600 52908 32612
rect 47572 31446 47618 31458
rect 47572 31154 47578 31446
rect 47612 31154 47618 31446
rect 47572 31142 47618 31154
rect 48630 31446 48676 31458
rect 48630 31154 48636 31446
rect 48670 31154 48676 31446
rect 48630 31142 48676 31154
rect 49688 31446 49734 31458
rect 49688 31154 49694 31446
rect 49728 31154 49734 31446
rect 49688 31142 49734 31154
rect 50746 31446 50792 31458
rect 50746 31154 50752 31446
rect 50786 31154 50792 31446
rect 50746 31142 50792 31154
rect 51804 31446 51850 31458
rect 51804 31154 51810 31446
rect 51844 31154 51850 31446
rect 51804 31142 51850 31154
rect 52862 31446 52908 31458
rect 52862 31154 52868 31446
rect 52902 31154 52908 31446
rect 52862 31142 52908 31154
rect 47572 30352 47618 30364
rect 47572 30060 47578 30352
rect 47612 30060 47618 30352
rect 47572 30048 47618 30060
rect 48630 30352 48676 30364
rect 48630 30060 48636 30352
rect 48670 30060 48676 30352
rect 48630 30048 48676 30060
rect 49688 30352 49734 30364
rect 49688 30060 49694 30352
rect 49728 30060 49734 30352
rect 49688 30048 49734 30060
rect 50746 30352 50792 30364
rect 50746 30060 50752 30352
rect 50786 30060 50792 30352
rect 50746 30048 50792 30060
rect 51804 30352 51850 30364
rect 51804 30060 51810 30352
rect 51844 30060 51850 30352
rect 51804 30048 51850 30060
rect 52862 30352 52908 30364
rect 52862 30060 52868 30352
rect 52902 30060 52908 30352
rect 52862 30048 52908 30060
rect 53442 30052 53776 34240
rect 59600 34446 59684 35834
rect 59892 34446 60012 35834
rect 76634 38916 76978 39082
rect 76634 35694 76760 38916
rect 76908 35694 76978 38916
rect 77164 38922 77170 39094
rect 77204 38922 77210 39094
rect 77164 38910 77210 38922
rect 77822 39094 77868 39106
rect 77822 38922 77828 39094
rect 77862 38922 77868 39094
rect 77822 38910 77868 38922
rect 78480 39094 78526 39106
rect 78480 38922 78486 39094
rect 78520 38922 78526 39094
rect 78480 38910 78526 38922
rect 79138 39094 79184 39106
rect 79138 38922 79144 39094
rect 79178 38922 79184 39094
rect 79138 38910 79184 38922
rect 79796 39094 79842 39106
rect 79796 38922 79802 39094
rect 79836 38922 79842 39094
rect 80440 39100 80534 39410
rect 80846 39444 80908 39470
rect 81068 39444 81140 39522
rect 80846 39390 81140 39444
rect 85028 39516 85372 39542
rect 85028 39420 85084 39516
rect 85284 39420 85372 39516
rect 85028 39402 85372 39420
rect 80440 39088 80536 39100
rect 79796 38910 79842 38922
rect 79960 38910 80304 39076
rect 80440 39050 80496 39088
rect 77164 38400 77210 38412
rect 77164 38228 77170 38400
rect 77204 38228 77210 38400
rect 77164 38216 77210 38228
rect 77822 38400 77868 38412
rect 77822 38228 77828 38400
rect 77862 38228 77868 38400
rect 77822 38216 77868 38228
rect 78480 38400 78526 38412
rect 78480 38228 78486 38400
rect 78520 38228 78526 38400
rect 78480 38216 78526 38228
rect 79138 38400 79184 38412
rect 79138 38228 79144 38400
rect 79178 38228 79184 38400
rect 79138 38216 79184 38228
rect 79796 38400 79842 38412
rect 79796 38228 79802 38400
rect 79836 38228 79842 38400
rect 79796 38216 79842 38228
rect 77164 37706 77210 37718
rect 77164 37534 77170 37706
rect 77204 37534 77210 37706
rect 77164 37522 77210 37534
rect 77822 37706 77868 37718
rect 77822 37534 77828 37706
rect 77862 37534 77868 37706
rect 77822 37522 77868 37534
rect 78480 37706 78526 37718
rect 78480 37534 78486 37706
rect 78520 37534 78526 37706
rect 78480 37522 78526 37534
rect 79138 37706 79184 37718
rect 79138 37534 79144 37706
rect 79178 37534 79184 37706
rect 79138 37522 79184 37534
rect 79796 37706 79842 37718
rect 79796 37534 79802 37706
rect 79836 37534 79842 37706
rect 79796 37522 79842 37534
rect 77164 37012 77210 37024
rect 77164 36840 77170 37012
rect 77204 36840 77210 37012
rect 77164 36828 77210 36840
rect 77822 37012 77868 37024
rect 77822 36840 77828 37012
rect 77862 36840 77868 37012
rect 77822 36828 77868 36840
rect 78480 37012 78526 37024
rect 78480 36840 78486 37012
rect 78520 36840 78526 37012
rect 78480 36828 78526 36840
rect 79138 37012 79184 37024
rect 79138 36840 79144 37012
rect 79178 36840 79184 37012
rect 79138 36828 79184 36840
rect 79796 37012 79842 37024
rect 79796 36840 79802 37012
rect 79836 36840 79842 37012
rect 79796 36828 79842 36840
rect 77164 36318 77210 36330
rect 77164 36146 77170 36318
rect 77204 36146 77210 36318
rect 77164 36134 77210 36146
rect 77822 36318 77868 36330
rect 77822 36146 77828 36318
rect 77862 36146 77868 36318
rect 77822 36134 77868 36146
rect 78480 36318 78526 36330
rect 78480 36146 78486 36318
rect 78520 36146 78526 36318
rect 78480 36134 78526 36146
rect 79138 36318 79184 36330
rect 79138 36146 79144 36318
rect 79178 36146 79184 36318
rect 79138 36134 79184 36146
rect 79796 36318 79842 36330
rect 79796 36146 79802 36318
rect 79836 36146 79842 36318
rect 79796 36134 79842 36146
rect 76634 35530 76978 35694
rect 79960 35688 80086 38910
rect 80234 35688 80304 38910
rect 80490 38916 80496 39050
rect 80530 38916 80536 39088
rect 80490 38904 80536 38916
rect 81148 39088 81194 39100
rect 81148 38916 81154 39088
rect 81188 38916 81194 39088
rect 81148 38904 81194 38916
rect 81806 39088 81852 39100
rect 81806 38916 81812 39088
rect 81846 38916 81852 39088
rect 81806 38904 81852 38916
rect 82464 39088 82510 39100
rect 82464 38916 82470 39088
rect 82504 38916 82510 39088
rect 82464 38904 82510 38916
rect 83122 39088 83168 39100
rect 83122 38916 83128 39088
rect 83162 38916 83168 39088
rect 83800 39088 83846 39100
rect 83122 38904 83168 38916
rect 83270 38910 83614 39076
rect 80490 38394 80536 38406
rect 80490 38222 80496 38394
rect 80530 38222 80536 38394
rect 80490 38210 80536 38222
rect 81148 38394 81194 38406
rect 81148 38222 81154 38394
rect 81188 38222 81194 38394
rect 81148 38210 81194 38222
rect 81806 38394 81852 38406
rect 81806 38222 81812 38394
rect 81846 38222 81852 38394
rect 81806 38210 81852 38222
rect 82464 38394 82510 38406
rect 82464 38222 82470 38394
rect 82504 38222 82510 38394
rect 82464 38210 82510 38222
rect 83122 38394 83168 38406
rect 83122 38222 83128 38394
rect 83162 38222 83168 38394
rect 83122 38210 83168 38222
rect 80490 37700 80536 37712
rect 80490 37528 80496 37700
rect 80530 37528 80536 37700
rect 80490 37516 80536 37528
rect 81148 37700 81194 37712
rect 81148 37528 81154 37700
rect 81188 37528 81194 37700
rect 81148 37516 81194 37528
rect 81806 37700 81852 37712
rect 81806 37528 81812 37700
rect 81846 37528 81852 37700
rect 81806 37516 81852 37528
rect 82464 37700 82510 37712
rect 82464 37528 82470 37700
rect 82504 37528 82510 37700
rect 82464 37516 82510 37528
rect 83122 37700 83168 37712
rect 83122 37528 83128 37700
rect 83162 37528 83168 37700
rect 83122 37516 83168 37528
rect 80490 37006 80536 37018
rect 80490 36834 80496 37006
rect 80530 36834 80536 37006
rect 80490 36822 80536 36834
rect 81148 37006 81194 37018
rect 81148 36834 81154 37006
rect 81188 36834 81194 37006
rect 81148 36822 81194 36834
rect 81806 37006 81852 37018
rect 81806 36834 81812 37006
rect 81846 36834 81852 37006
rect 81806 36822 81852 36834
rect 82464 37006 82510 37018
rect 82464 36834 82470 37006
rect 82504 36834 82510 37006
rect 82464 36822 82510 36834
rect 83122 37006 83168 37018
rect 83122 36834 83128 37006
rect 83162 36834 83168 37006
rect 83122 36822 83168 36834
rect 80490 36312 80536 36324
rect 80490 36140 80496 36312
rect 80530 36140 80536 36312
rect 80490 36128 80536 36140
rect 81148 36312 81194 36324
rect 81148 36140 81154 36312
rect 81188 36140 81194 36312
rect 81148 36128 81194 36140
rect 81806 36312 81852 36324
rect 81806 36140 81812 36312
rect 81846 36140 81852 36312
rect 81806 36128 81852 36140
rect 82464 36312 82510 36324
rect 82464 36140 82470 36312
rect 82504 36140 82510 36312
rect 82464 36128 82510 36140
rect 83122 36312 83168 36324
rect 83122 36140 83128 36312
rect 83162 36140 83168 36312
rect 83122 36128 83168 36140
rect 77164 35624 77210 35636
rect 76680 34874 76932 35530
rect 77164 35452 77170 35624
rect 77204 35452 77210 35624
rect 77164 35440 77210 35452
rect 77822 35624 77868 35636
rect 77822 35452 77828 35624
rect 77862 35452 77868 35624
rect 77822 35440 77868 35452
rect 78480 35624 78526 35636
rect 78480 35452 78486 35624
rect 78520 35452 78526 35624
rect 78480 35440 78526 35452
rect 79138 35624 79184 35636
rect 79138 35452 79144 35624
rect 79178 35452 79184 35624
rect 79138 35440 79184 35452
rect 79796 35624 79842 35636
rect 79796 35452 79802 35624
rect 79836 35452 79842 35624
rect 79960 35524 80304 35688
rect 83270 35688 83396 38910
rect 83544 35688 83614 38910
rect 83800 38916 83806 39088
rect 83840 38916 83846 39088
rect 83800 38904 83846 38916
rect 84458 39088 84504 39100
rect 84458 38916 84464 39088
rect 84498 38916 84504 39088
rect 84458 38904 84504 38916
rect 85116 39088 85162 39100
rect 85116 38916 85122 39088
rect 85156 38916 85162 39088
rect 85116 38904 85162 38916
rect 85774 39088 85820 39100
rect 85774 38916 85780 39088
rect 85814 38916 85820 39088
rect 85774 38904 85820 38916
rect 86432 39088 86478 39100
rect 86432 38916 86438 39088
rect 86472 38916 86478 39088
rect 86432 38904 86478 38916
rect 86688 38988 87154 40396
rect 88846 40376 89414 40396
rect 86688 38762 86786 38988
rect 83800 38394 83846 38406
rect 83800 38222 83806 38394
rect 83840 38222 83846 38394
rect 83800 38210 83846 38222
rect 84458 38394 84504 38406
rect 84458 38222 84464 38394
rect 84498 38222 84504 38394
rect 84458 38210 84504 38222
rect 85116 38394 85162 38406
rect 85116 38222 85122 38394
rect 85156 38222 85162 38394
rect 85116 38210 85162 38222
rect 85774 38394 85820 38406
rect 85774 38222 85780 38394
rect 85814 38222 85820 38394
rect 85774 38210 85820 38222
rect 86432 38394 86478 38406
rect 86432 38222 86438 38394
rect 86472 38222 86478 38394
rect 86432 38210 86478 38222
rect 83800 37700 83846 37712
rect 83800 37528 83806 37700
rect 83840 37528 83846 37700
rect 83800 37516 83846 37528
rect 84458 37700 84504 37712
rect 84458 37528 84464 37700
rect 84498 37528 84504 37700
rect 84458 37516 84504 37528
rect 85116 37700 85162 37712
rect 85116 37528 85122 37700
rect 85156 37528 85162 37700
rect 85116 37516 85162 37528
rect 85774 37700 85820 37712
rect 85774 37528 85780 37700
rect 85814 37528 85820 37700
rect 85774 37516 85820 37528
rect 86432 37700 86478 37712
rect 86432 37528 86438 37700
rect 86472 37528 86478 37700
rect 86432 37516 86478 37528
rect 83800 37006 83846 37018
rect 83800 36834 83806 37006
rect 83840 36834 83846 37006
rect 83800 36822 83846 36834
rect 84458 37006 84504 37018
rect 84458 36834 84464 37006
rect 84498 36834 84504 37006
rect 84458 36822 84504 36834
rect 85116 37006 85162 37018
rect 85116 36834 85122 37006
rect 85156 36834 85162 37006
rect 85116 36822 85162 36834
rect 85774 37006 85820 37018
rect 85774 36834 85780 37006
rect 85814 36834 85820 37006
rect 85774 36822 85820 36834
rect 86432 37006 86478 37018
rect 86432 36834 86438 37006
rect 86472 36834 86478 37006
rect 86432 36822 86478 36834
rect 83800 36312 83846 36324
rect 83800 36140 83806 36312
rect 83840 36140 83846 36312
rect 83800 36128 83846 36140
rect 84458 36312 84504 36324
rect 84458 36140 84464 36312
rect 84498 36140 84504 36312
rect 84458 36128 84504 36140
rect 85116 36312 85162 36324
rect 85116 36140 85122 36312
rect 85156 36140 85162 36312
rect 85116 36128 85162 36140
rect 85774 36312 85820 36324
rect 85774 36140 85780 36312
rect 85814 36140 85820 36312
rect 85774 36128 85820 36140
rect 86432 36312 86478 36324
rect 86432 36140 86438 36312
rect 86472 36140 86478 36312
rect 86432 36128 86478 36140
rect 80490 35618 80536 35630
rect 79796 35440 79842 35452
rect 80016 34874 80268 35524
rect 80490 35446 80496 35618
rect 80530 35446 80536 35618
rect 81148 35618 81194 35630
rect 81148 35554 81154 35618
rect 80490 35434 80536 35446
rect 81094 35446 81154 35554
rect 81188 35554 81194 35618
rect 81806 35618 81852 35630
rect 81188 35446 81226 35554
rect 81094 34874 81226 35446
rect 81806 35446 81812 35618
rect 81846 35446 81852 35618
rect 81806 35434 81852 35446
rect 82464 35618 82510 35630
rect 82464 35446 82470 35618
rect 82504 35446 82510 35618
rect 82464 35434 82510 35446
rect 83122 35618 83168 35630
rect 83122 35446 83128 35618
rect 83162 35446 83168 35618
rect 83270 35524 83614 35688
rect 86696 35656 86786 38762
rect 86904 38762 87154 38988
rect 86904 35656 87008 38762
rect 83800 35618 83846 35630
rect 83122 35434 83168 35446
rect 83336 34874 83588 35524
rect 83800 35446 83806 35618
rect 83840 35446 83846 35618
rect 83800 35434 83846 35446
rect 84458 35618 84504 35630
rect 84458 35446 84464 35618
rect 84498 35446 84504 35618
rect 84458 35434 84504 35446
rect 85116 35618 85162 35630
rect 85116 35446 85122 35618
rect 85156 35446 85162 35618
rect 85116 35434 85162 35446
rect 85774 35618 85820 35630
rect 85774 35446 85780 35618
rect 85814 35446 85820 35618
rect 85774 35434 85820 35446
rect 86432 35618 86478 35630
rect 86432 35446 86438 35618
rect 86472 35446 86478 35618
rect 86432 35434 86478 35446
rect 86696 35242 87008 35656
rect 86710 34874 86962 35242
rect 76680 34670 86964 34874
rect 83336 34628 83588 34670
rect 59600 34156 60012 34446
rect 54086 34012 54132 34024
rect 54086 33720 54092 34012
rect 54126 33720 54132 34012
rect 54086 33708 54132 33720
rect 55144 34012 55190 34024
rect 55144 33720 55150 34012
rect 55184 33720 55190 34012
rect 55144 33708 55190 33720
rect 56202 34012 56248 34024
rect 56202 33720 56208 34012
rect 56242 33720 56248 34012
rect 56202 33708 56248 33720
rect 57260 34012 57306 34024
rect 57260 33720 57266 34012
rect 57300 33720 57306 34012
rect 57260 33708 57306 33720
rect 58318 34012 58364 34024
rect 58318 33720 58324 34012
rect 58358 33720 58364 34012
rect 58318 33708 58364 33720
rect 59376 34012 59422 34024
rect 59376 33720 59382 34012
rect 59416 33720 59422 34012
rect 59376 33708 59422 33720
rect 54086 32918 54132 32930
rect 54086 32626 54092 32918
rect 54126 32626 54132 32918
rect 54086 32614 54132 32626
rect 55144 32918 55190 32930
rect 55144 32626 55150 32918
rect 55184 32626 55190 32918
rect 55144 32614 55190 32626
rect 56202 32918 56248 32930
rect 56202 32626 56208 32918
rect 56242 32626 56248 32918
rect 56202 32614 56248 32626
rect 57260 32918 57306 32930
rect 57260 32626 57266 32918
rect 57300 32626 57306 32918
rect 57260 32614 57306 32626
rect 58318 32918 58364 32930
rect 58318 32626 58324 32918
rect 58358 32626 58364 32918
rect 58318 32614 58364 32626
rect 59376 32918 59422 32930
rect 59376 32626 59382 32918
rect 59416 32626 59422 32918
rect 59376 32614 59422 32626
rect 54086 31460 54132 31472
rect 54086 31168 54092 31460
rect 54126 31168 54132 31460
rect 54086 31156 54132 31168
rect 55144 31460 55190 31472
rect 55144 31168 55150 31460
rect 55184 31168 55190 31460
rect 55144 31156 55190 31168
rect 56202 31460 56248 31472
rect 56202 31168 56208 31460
rect 56242 31168 56248 31460
rect 56202 31156 56248 31168
rect 57260 31460 57306 31472
rect 57260 31168 57266 31460
rect 57300 31168 57306 31460
rect 57260 31156 57306 31168
rect 58318 31460 58364 31472
rect 58318 31168 58324 31460
rect 58358 31168 58364 31460
rect 58318 31156 58364 31168
rect 59376 31460 59422 31472
rect 59376 31168 59382 31460
rect 59416 31168 59422 31460
rect 59376 31156 59422 31168
rect 54086 30366 54132 30378
rect 54086 30074 54092 30366
rect 54126 30074 54132 30366
rect 54086 30062 54132 30074
rect 55144 30366 55190 30378
rect 55144 30074 55150 30366
rect 55184 30074 55190 30366
rect 55144 30062 55190 30074
rect 56202 30366 56248 30378
rect 56202 30074 56208 30366
rect 56242 30074 56248 30366
rect 56202 30062 56248 30074
rect 57260 30366 57306 30378
rect 57260 30074 57266 30366
rect 57300 30074 57306 30366
rect 57260 30062 57306 30074
rect 58318 30366 58364 30378
rect 58318 30074 58324 30366
rect 58358 30074 58364 30366
rect 58318 30062 58364 30074
rect 59376 30366 59422 30378
rect 59376 30074 59382 30366
rect 59416 30074 59422 30366
rect 59680 30090 60012 34156
rect 59376 30062 59422 30074
rect 40984 29236 41030 29248
rect 40984 28944 40990 29236
rect 41024 28944 41030 29236
rect 40984 28932 41030 28944
rect 42042 29236 42088 29248
rect 42042 28944 42048 29236
rect 42082 28944 42088 29236
rect 42042 28932 42088 28944
rect 43100 29236 43146 29248
rect 43100 28944 43106 29236
rect 43140 28944 43146 29236
rect 43100 28932 43146 28944
rect 44158 29236 44204 29248
rect 44158 28944 44164 29236
rect 44198 28944 44204 29236
rect 44158 28932 44204 28944
rect 45216 29236 45262 29248
rect 45216 28944 45222 29236
rect 45256 28944 45262 29236
rect 45216 28932 45262 28944
rect 46274 29236 46320 29248
rect 46274 28944 46280 29236
rect 46314 28944 46320 29236
rect 46274 28932 46320 28944
rect 34494 28142 34540 28154
rect 34494 27850 34500 28142
rect 34534 27850 34540 28142
rect 34494 27838 34540 27850
rect 35552 28142 35598 28154
rect 35552 27850 35558 28142
rect 35592 27850 35598 28142
rect 35552 27838 35598 27850
rect 36610 28142 36656 28154
rect 36610 27850 36616 28142
rect 36650 27850 36656 28142
rect 36610 27838 36656 27850
rect 37668 28142 37714 28154
rect 37668 27850 37674 28142
rect 37708 27850 37714 28142
rect 37668 27838 37714 27850
rect 38726 28142 38772 28154
rect 38726 27850 38732 28142
rect 38766 27850 38772 28142
rect 38726 27838 38772 27850
rect 39784 28142 39830 28154
rect 39784 27850 39790 28142
rect 39824 27850 39830 28142
rect 39784 27838 39830 27850
rect 34494 27048 34540 27060
rect 34494 26756 34500 27048
rect 34534 26756 34540 27048
rect 34494 26744 34540 26756
rect 35552 27048 35598 27060
rect 35552 26756 35558 27048
rect 35592 26756 35598 27048
rect 35552 26744 35598 26756
rect 36610 27048 36656 27060
rect 36610 26756 36616 27048
rect 36650 26756 36656 27048
rect 36610 26744 36656 26756
rect 37668 27048 37714 27060
rect 37668 26756 37674 27048
rect 37708 26756 37714 27048
rect 37668 26744 37714 26756
rect 38726 27048 38772 27060
rect 38726 26756 38732 27048
rect 38766 26756 38772 27048
rect 38726 26744 38772 26756
rect 39784 27048 39830 27060
rect 39784 26756 39790 27048
rect 39824 26756 39830 27048
rect 39784 26744 39830 26756
rect 34494 25588 34540 25600
rect 34494 25296 34500 25588
rect 34534 25296 34540 25588
rect 34494 25284 34540 25296
rect 35552 25588 35598 25600
rect 35552 25296 35558 25588
rect 35592 25296 35598 25588
rect 35552 25284 35598 25296
rect 36610 25588 36656 25600
rect 36610 25296 36616 25588
rect 36650 25296 36656 25588
rect 36610 25284 36656 25296
rect 37668 25588 37714 25600
rect 37668 25296 37674 25588
rect 37708 25296 37714 25588
rect 37668 25284 37714 25296
rect 38726 25588 38772 25600
rect 38726 25296 38732 25588
rect 38766 25296 38772 25588
rect 38726 25284 38772 25296
rect 39784 25588 39830 25600
rect 39784 25296 39790 25588
rect 39824 25296 39830 25588
rect 39784 25284 39830 25296
rect 34494 24494 34540 24506
rect 34494 24202 34500 24494
rect 34534 24202 34540 24494
rect 34494 24190 34540 24202
rect 35552 24494 35598 24506
rect 35552 24202 35558 24494
rect 35592 24202 35598 24494
rect 35552 24190 35598 24202
rect 36610 24494 36656 24506
rect 36610 24202 36616 24494
rect 36650 24202 36656 24494
rect 36610 24190 36656 24202
rect 37668 24494 37714 24506
rect 37668 24202 37674 24494
rect 37708 24202 37714 24494
rect 37668 24190 37714 24202
rect 38726 24494 38772 24506
rect 38726 24202 38732 24494
rect 38766 24202 38772 24494
rect 38726 24190 38772 24202
rect 39784 24494 39830 24506
rect 39784 24202 39790 24494
rect 39824 24202 39830 24494
rect 39784 24190 39830 24202
rect 21462 23378 21508 23390
rect 21462 23086 21468 23378
rect 21502 23086 21508 23378
rect 21462 23074 21508 23086
rect 22520 23378 22566 23390
rect 22520 23086 22526 23378
rect 22560 23086 22566 23378
rect 22520 23074 22566 23086
rect 23578 23378 23624 23390
rect 23578 23086 23584 23378
rect 23618 23086 23624 23378
rect 23578 23074 23624 23086
rect 24636 23378 24682 23390
rect 24636 23086 24642 23378
rect 24676 23086 24682 23378
rect 24636 23074 24682 23086
rect 25694 23378 25740 23390
rect 25694 23086 25700 23378
rect 25734 23086 25740 23378
rect 25694 23074 25740 23086
rect 26752 23378 26798 23390
rect 26752 23086 26758 23378
rect 26792 23086 26798 23378
rect 26752 23074 26798 23086
rect 14972 22300 15018 22312
rect 14972 22008 14978 22300
rect 15012 22008 15018 22300
rect 14972 21996 15018 22008
rect 16030 22300 16076 22312
rect 16030 22008 16036 22300
rect 16070 22008 16076 22300
rect 16030 21996 16076 22008
rect 17088 22300 17134 22312
rect 17088 22008 17094 22300
rect 17128 22008 17134 22300
rect 17088 21996 17134 22008
rect 18146 22300 18192 22312
rect 18146 22008 18152 22300
rect 18186 22008 18192 22300
rect 18146 21996 18192 22008
rect 19204 22300 19250 22312
rect 19204 22008 19210 22300
rect 19244 22008 19250 22300
rect 19204 21996 19250 22008
rect 20262 22300 20308 22312
rect 20262 22008 20268 22300
rect 20302 22008 20308 22300
rect 20262 21996 20308 22008
rect 14972 21206 15018 21218
rect 14972 20914 14978 21206
rect 15012 20914 15018 21206
rect 14972 20902 15018 20914
rect 16030 21206 16076 21218
rect 16030 20914 16036 21206
rect 16070 20914 16076 21206
rect 16030 20902 16076 20914
rect 17088 21206 17134 21218
rect 17088 20914 17094 21206
rect 17128 20914 17134 21206
rect 17088 20902 17134 20914
rect 18146 21206 18192 21218
rect 18146 20914 18152 21206
rect 18186 20914 18192 21206
rect 18146 20902 18192 20914
rect 19204 21206 19250 21218
rect 19204 20914 19210 21206
rect 19244 20914 19250 21206
rect 19204 20902 19250 20914
rect 20262 21206 20308 21218
rect 20262 20914 20268 21206
rect 20302 20914 20308 21206
rect 20262 20902 20308 20914
rect 14972 19718 15018 19730
rect 14972 19426 14978 19718
rect 15012 19426 15018 19718
rect 14972 19414 15018 19426
rect 16030 19718 16076 19730
rect 16030 19426 16036 19718
rect 16070 19426 16076 19718
rect 16030 19414 16076 19426
rect 17088 19718 17134 19730
rect 17088 19426 17094 19718
rect 17128 19426 17134 19718
rect 17088 19414 17134 19426
rect 18146 19718 18192 19730
rect 18146 19426 18152 19718
rect 18186 19426 18192 19718
rect 18146 19414 18192 19426
rect 19204 19718 19250 19730
rect 19204 19426 19210 19718
rect 19244 19426 19250 19718
rect 19204 19414 19250 19426
rect 20262 19718 20308 19730
rect 20262 19426 20268 19718
rect 20302 19426 20308 19718
rect 20262 19414 20308 19426
rect 14972 18624 15018 18636
rect 14972 18332 14978 18624
rect 15012 18332 15018 18624
rect 14972 18320 15018 18332
rect 16030 18624 16076 18636
rect 16030 18332 16036 18624
rect 16070 18332 16076 18624
rect 16030 18320 16076 18332
rect 17088 18624 17134 18636
rect 17088 18332 17094 18624
rect 17128 18332 17134 18624
rect 17088 18320 17134 18332
rect 18146 18624 18192 18636
rect 18146 18332 18152 18624
rect 18186 18332 18192 18624
rect 18146 18320 18192 18332
rect 19204 18624 19250 18636
rect 19204 18332 19210 18624
rect 19244 18332 19250 18624
rect 19204 18320 19250 18332
rect 20262 18624 20308 18636
rect 20262 18332 20268 18624
rect 20302 18332 20308 18624
rect 20262 18320 20308 18332
rect 8466 17522 8512 17534
rect 8466 17230 8472 17522
rect 8506 17230 8512 17522
rect 8466 17218 8512 17230
rect 9524 17522 9570 17534
rect 9524 17230 9530 17522
rect 9564 17230 9570 17522
rect 9524 17218 9570 17230
rect 10582 17522 10628 17534
rect 10582 17230 10588 17522
rect 10622 17230 10628 17522
rect 10582 17218 10628 17230
rect 11640 17522 11686 17534
rect 11640 17230 11646 17522
rect 11680 17230 11686 17522
rect 11640 17218 11686 17230
rect 12698 17522 12744 17534
rect 12698 17230 12704 17522
rect 12738 17230 12744 17522
rect 12698 17218 12744 17230
rect 13756 17522 13802 17534
rect 13756 17230 13762 17522
rect 13796 17230 13802 17522
rect 13756 17218 13802 17230
rect 1952 16420 1998 16432
rect 1952 16128 1958 16420
rect 1992 16128 1998 16420
rect 1952 16116 1998 16128
rect 3010 16420 3056 16432
rect 3010 16128 3016 16420
rect 3050 16128 3056 16420
rect 3010 16116 3056 16128
rect 4068 16420 4114 16432
rect 4068 16128 4074 16420
rect 4108 16128 4114 16420
rect 4068 16116 4114 16128
rect 5126 16420 5172 16432
rect 5126 16128 5132 16420
rect 5166 16128 5172 16420
rect 5126 16116 5172 16128
rect 6184 16420 6230 16432
rect 6184 16128 6190 16420
rect 6224 16128 6230 16420
rect 6184 16116 6230 16128
rect 7242 16420 7288 16432
rect 7242 16128 7248 16420
rect 7282 16128 7288 16420
rect 7242 16116 7288 16128
rect 1952 15326 1998 15338
rect 1952 15034 1958 15326
rect 1992 15034 1998 15326
rect 1952 15022 1998 15034
rect 3010 15326 3056 15338
rect 3010 15034 3016 15326
rect 3050 15034 3056 15326
rect 3010 15022 3056 15034
rect 4068 15326 4114 15338
rect 4068 15034 4074 15326
rect 4108 15034 4114 15326
rect 4068 15022 4114 15034
rect 5126 15326 5172 15338
rect 5126 15034 5132 15326
rect 5166 15034 5172 15326
rect 5126 15022 5172 15034
rect 6184 15326 6230 15338
rect 6184 15034 6190 15326
rect 6224 15034 6230 15326
rect 6184 15022 6230 15034
rect 7242 15326 7288 15338
rect 7242 15034 7248 15326
rect 7282 15034 7288 15326
rect 7242 15022 7288 15034
rect 1962 13846 2008 13858
rect 1962 13554 1968 13846
rect 2002 13554 2008 13846
rect 1962 13542 2008 13554
rect 3020 13846 3066 13858
rect 3020 13554 3026 13846
rect 3060 13554 3066 13846
rect 3020 13542 3066 13554
rect 4078 13846 4124 13858
rect 4078 13554 4084 13846
rect 4118 13554 4124 13846
rect 4078 13542 4124 13554
rect 5136 13846 5182 13858
rect 5136 13554 5142 13846
rect 5176 13554 5182 13846
rect 5136 13542 5182 13554
rect 6194 13846 6240 13858
rect 6194 13554 6200 13846
rect 6234 13554 6240 13846
rect 6194 13542 6240 13554
rect 7252 13846 7298 13858
rect 7252 13554 7258 13846
rect 7292 13554 7298 13846
rect 7252 13542 7298 13554
rect 1962 12752 2008 12764
rect 1962 12460 1968 12752
rect 2002 12460 2008 12752
rect 1962 12448 2008 12460
rect 3020 12752 3066 12764
rect 3020 12460 3026 12752
rect 3060 12460 3066 12752
rect 3020 12448 3066 12460
rect 4078 12752 4124 12764
rect 4078 12460 4084 12752
rect 4118 12460 4124 12752
rect 4078 12448 4124 12460
rect 5136 12752 5182 12764
rect 5136 12460 5142 12752
rect 5176 12460 5182 12752
rect 5136 12448 5182 12460
rect 6194 12752 6240 12764
rect 6194 12460 6200 12752
rect 6234 12460 6240 12752
rect 6194 12448 6240 12460
rect 7252 12752 7298 12764
rect 7252 12460 7258 12752
rect 7292 12460 7298 12752
rect 7252 12448 7298 12460
rect 1264 11116 1336 12312
rect 1430 11116 1560 12312
rect 7722 12320 8018 16980
rect 14216 16988 14346 18184
rect 14440 16988 14512 18184
rect 20748 18168 21044 22836
rect 27278 22852 27358 24048
rect 27452 22852 27574 24048
rect 33846 24054 34144 24180
rect 27984 23394 28030 23406
rect 27984 23102 27990 23394
rect 28024 23102 28030 23394
rect 27984 23090 28030 23102
rect 29042 23394 29088 23406
rect 29042 23102 29048 23394
rect 29082 23102 29088 23394
rect 29042 23090 29088 23102
rect 30100 23394 30146 23406
rect 30100 23102 30106 23394
rect 30140 23102 30146 23394
rect 30100 23090 30146 23102
rect 31158 23394 31204 23406
rect 31158 23102 31164 23394
rect 31198 23102 31204 23394
rect 31158 23090 31204 23102
rect 32216 23394 32262 23406
rect 32216 23102 32222 23394
rect 32256 23102 32262 23394
rect 32216 23090 32262 23102
rect 33274 23394 33320 23406
rect 33274 23102 33280 23394
rect 33314 23102 33320 23394
rect 33274 23090 33320 23102
rect 21462 22284 21508 22296
rect 21462 21992 21468 22284
rect 21502 21992 21508 22284
rect 21462 21980 21508 21992
rect 22520 22284 22566 22296
rect 22520 21992 22526 22284
rect 22560 21992 22566 22284
rect 22520 21980 22566 21992
rect 23578 22284 23624 22296
rect 23578 21992 23584 22284
rect 23618 21992 23624 22284
rect 23578 21980 23624 21992
rect 24636 22284 24682 22296
rect 24636 21992 24642 22284
rect 24676 21992 24682 22284
rect 24636 21980 24682 21992
rect 25694 22284 25740 22296
rect 25694 21992 25700 22284
rect 25734 21992 25740 22284
rect 25694 21980 25740 21992
rect 26752 22284 26798 22296
rect 26752 21992 26758 22284
rect 26792 21992 26798 22284
rect 26752 21980 26798 21992
rect 21462 21190 21508 21202
rect 21462 20898 21468 21190
rect 21502 20898 21508 21190
rect 21462 20886 21508 20898
rect 22520 21190 22566 21202
rect 22520 20898 22526 21190
rect 22560 20898 22566 21190
rect 22520 20886 22566 20898
rect 23578 21190 23624 21202
rect 23578 20898 23584 21190
rect 23618 20898 23624 21190
rect 23578 20886 23624 20898
rect 24636 21190 24682 21202
rect 24636 20898 24642 21190
rect 24676 20898 24682 21190
rect 24636 20886 24682 20898
rect 25694 21190 25740 21202
rect 25694 20898 25700 21190
rect 25734 20898 25740 21190
rect 25694 20886 25740 20898
rect 26752 21190 26798 21202
rect 26752 20898 26758 21190
rect 26792 20898 26798 21190
rect 26752 20886 26798 20898
rect 21462 19702 21508 19714
rect 21462 19410 21468 19702
rect 21502 19410 21508 19702
rect 21462 19398 21508 19410
rect 22520 19702 22566 19714
rect 22520 19410 22526 19702
rect 22560 19410 22566 19702
rect 22520 19398 22566 19410
rect 23578 19702 23624 19714
rect 23578 19410 23584 19702
rect 23618 19410 23624 19702
rect 23578 19398 23624 19410
rect 24636 19702 24682 19714
rect 24636 19410 24642 19702
rect 24676 19410 24682 19702
rect 24636 19398 24682 19410
rect 25694 19702 25740 19714
rect 25694 19410 25700 19702
rect 25734 19410 25740 19702
rect 25694 19398 25740 19410
rect 26752 19702 26798 19714
rect 26752 19410 26758 19702
rect 26792 19410 26798 19702
rect 26752 19398 26798 19410
rect 21462 18608 21508 18620
rect 21462 18316 21468 18608
rect 21502 18316 21508 18608
rect 21462 18304 21508 18316
rect 22520 18608 22566 18620
rect 22520 18316 22526 18608
rect 22560 18316 22566 18608
rect 22520 18304 22566 18316
rect 23578 18608 23624 18620
rect 23578 18316 23584 18608
rect 23618 18316 23624 18608
rect 23578 18304 23624 18316
rect 24636 18608 24682 18620
rect 24636 18316 24642 18608
rect 24676 18316 24682 18608
rect 24636 18304 24682 18316
rect 25694 18608 25740 18620
rect 25694 18316 25700 18608
rect 25734 18316 25740 18608
rect 25694 18304 25740 18316
rect 26752 18608 26798 18620
rect 26752 18316 26758 18608
rect 26792 18316 26798 18608
rect 26752 18304 26798 18316
rect 14972 17530 15018 17542
rect 14972 17238 14978 17530
rect 15012 17238 15018 17530
rect 14972 17226 15018 17238
rect 16030 17530 16076 17542
rect 16030 17238 16036 17530
rect 16070 17238 16076 17530
rect 16030 17226 16076 17238
rect 17088 17530 17134 17542
rect 17088 17238 17094 17530
rect 17128 17238 17134 17530
rect 17088 17226 17134 17238
rect 18146 17530 18192 17542
rect 18146 17238 18152 17530
rect 18186 17238 18192 17530
rect 18146 17226 18192 17238
rect 19204 17530 19250 17542
rect 19204 17238 19210 17530
rect 19244 17238 19250 17530
rect 19204 17226 19250 17238
rect 20262 17530 20308 17542
rect 20262 17238 20268 17530
rect 20302 17238 20308 17530
rect 20262 17226 20308 17238
rect 8466 16428 8512 16440
rect 8466 16136 8472 16428
rect 8506 16136 8512 16428
rect 8466 16124 8512 16136
rect 9524 16428 9570 16440
rect 9524 16136 9530 16428
rect 9564 16136 9570 16428
rect 9524 16124 9570 16136
rect 10582 16428 10628 16440
rect 10582 16136 10588 16428
rect 10622 16136 10628 16428
rect 10582 16124 10628 16136
rect 11640 16428 11686 16440
rect 11640 16136 11646 16428
rect 11680 16136 11686 16428
rect 11640 16124 11686 16136
rect 12698 16428 12744 16440
rect 12698 16136 12704 16428
rect 12738 16136 12744 16428
rect 12698 16124 12744 16136
rect 13756 16428 13802 16440
rect 13756 16136 13762 16428
rect 13796 16136 13802 16428
rect 13756 16124 13802 16136
rect 8466 15334 8512 15346
rect 8466 15042 8472 15334
rect 8506 15042 8512 15334
rect 8466 15030 8512 15042
rect 9524 15334 9570 15346
rect 9524 15042 9530 15334
rect 9564 15042 9570 15334
rect 9524 15030 9570 15042
rect 10582 15334 10628 15346
rect 10582 15042 10588 15334
rect 10622 15042 10628 15334
rect 10582 15030 10628 15042
rect 11640 15334 11686 15346
rect 11640 15042 11646 15334
rect 11680 15042 11686 15334
rect 11640 15030 11686 15042
rect 12698 15334 12744 15346
rect 12698 15042 12704 15334
rect 12738 15042 12744 15334
rect 12698 15030 12744 15042
rect 13756 15334 13802 15346
rect 13756 15042 13762 15334
rect 13796 15042 13802 15334
rect 13756 15030 13802 15042
rect 8476 13854 8522 13866
rect 8476 13562 8482 13854
rect 8516 13562 8522 13854
rect 8476 13550 8522 13562
rect 9534 13854 9580 13866
rect 9534 13562 9540 13854
rect 9574 13562 9580 13854
rect 9534 13550 9580 13562
rect 10592 13854 10638 13866
rect 10592 13562 10598 13854
rect 10632 13562 10638 13854
rect 10592 13550 10638 13562
rect 11650 13854 11696 13866
rect 11650 13562 11656 13854
rect 11690 13562 11696 13854
rect 11650 13550 11696 13562
rect 12708 13854 12754 13866
rect 12708 13562 12714 13854
rect 12748 13562 12754 13854
rect 12708 13550 12754 13562
rect 13766 13854 13812 13866
rect 13766 13562 13772 13854
rect 13806 13562 13812 13854
rect 13766 13550 13812 13562
rect 8476 12760 8522 12772
rect 8476 12468 8482 12760
rect 8516 12468 8522 12760
rect 8476 12456 8522 12468
rect 9534 12760 9580 12772
rect 9534 12468 9540 12760
rect 9574 12468 9580 12760
rect 9534 12456 9580 12468
rect 10592 12760 10638 12772
rect 10592 12468 10598 12760
rect 10632 12468 10638 12760
rect 10592 12456 10638 12468
rect 11650 12760 11696 12772
rect 11650 12468 11656 12760
rect 11690 12468 11696 12760
rect 11650 12456 11696 12468
rect 12708 12760 12754 12772
rect 12708 12468 12714 12760
rect 12748 12468 12754 12760
rect 12708 12456 12754 12468
rect 13766 12760 13812 12772
rect 13766 12468 13772 12760
rect 13806 12468 13812 12760
rect 13766 12456 13812 12468
rect 1962 11658 2008 11670
rect 1962 11366 1968 11658
rect 2002 11366 2008 11658
rect 1962 11354 2008 11366
rect 3020 11658 3066 11670
rect 3020 11366 3026 11658
rect 3060 11366 3066 11658
rect 3020 11354 3066 11366
rect 4078 11658 4124 11670
rect 4078 11366 4084 11658
rect 4118 11366 4124 11658
rect 4078 11354 4124 11366
rect 5136 11658 5182 11670
rect 5136 11366 5142 11658
rect 5176 11366 5182 11658
rect 5136 11354 5182 11366
rect 6194 11658 6240 11670
rect 6194 11366 6200 11658
rect 6234 11366 6240 11658
rect 6194 11354 6240 11366
rect 7252 11658 7298 11670
rect 7252 11366 7258 11658
rect 7292 11366 7298 11658
rect 7252 11354 7298 11366
rect 1264 6404 1560 11116
rect 7722 11124 7850 12320
rect 7944 11124 8018 12320
rect 14216 12328 14512 16988
rect 20748 16972 20836 18168
rect 20930 16972 21044 18168
rect 27278 18184 27574 22852
rect 33846 22858 33868 24054
rect 33962 22858 34144 24054
rect 40304 24054 40638 28694
rect 46836 28716 46946 29912
rect 47040 28716 47170 29912
rect 53438 29926 53776 30052
rect 47572 29258 47618 29270
rect 47572 28966 47578 29258
rect 47612 28966 47618 29258
rect 47572 28954 47618 28966
rect 48630 29258 48676 29270
rect 48630 28966 48636 29258
rect 48670 28966 48676 29258
rect 48630 28954 48676 28966
rect 49688 29258 49734 29270
rect 49688 28966 49694 29258
rect 49728 28966 49734 29258
rect 49688 28954 49734 28966
rect 50746 29258 50792 29270
rect 50746 28966 50752 29258
rect 50786 28966 50792 29258
rect 50746 28954 50792 28966
rect 51804 29258 51850 29270
rect 51804 28966 51810 29258
rect 51844 28966 51850 29258
rect 51804 28954 51850 28966
rect 52862 29258 52908 29270
rect 52862 28966 52868 29258
rect 52902 28966 52908 29258
rect 52862 28954 52908 28966
rect 40984 28142 41030 28154
rect 40984 27850 40990 28142
rect 41024 27850 41030 28142
rect 40984 27838 41030 27850
rect 42042 28142 42088 28154
rect 42042 27850 42048 28142
rect 42082 27850 42088 28142
rect 42042 27838 42088 27850
rect 43100 28142 43146 28154
rect 43100 27850 43106 28142
rect 43140 27850 43146 28142
rect 43100 27838 43146 27850
rect 44158 28142 44204 28154
rect 44158 27850 44164 28142
rect 44198 27850 44204 28142
rect 44158 27838 44204 27850
rect 45216 28142 45262 28154
rect 45216 27850 45222 28142
rect 45256 27850 45262 28142
rect 45216 27838 45262 27850
rect 46274 28142 46320 28154
rect 46274 27850 46280 28142
rect 46314 27850 46320 28142
rect 46274 27838 46320 27850
rect 40984 27048 41030 27060
rect 40984 26756 40990 27048
rect 41024 26756 41030 27048
rect 40984 26744 41030 26756
rect 42042 27048 42088 27060
rect 42042 26756 42048 27048
rect 42082 26756 42088 27048
rect 42042 26744 42088 26756
rect 43100 27048 43146 27060
rect 43100 26756 43106 27048
rect 43140 26756 43146 27048
rect 43100 26744 43146 26756
rect 44158 27048 44204 27060
rect 44158 26756 44164 27048
rect 44198 26756 44204 27048
rect 44158 26744 44204 26756
rect 45216 27048 45262 27060
rect 45216 26756 45222 27048
rect 45256 26756 45262 27048
rect 45216 26744 45262 26756
rect 46274 27048 46320 27060
rect 46274 26756 46280 27048
rect 46314 26756 46320 27048
rect 46274 26744 46320 26756
rect 40984 25588 41030 25600
rect 40984 25296 40990 25588
rect 41024 25296 41030 25588
rect 40984 25284 41030 25296
rect 42042 25588 42088 25600
rect 42042 25296 42048 25588
rect 42082 25296 42088 25588
rect 42042 25284 42088 25296
rect 43100 25588 43146 25600
rect 43100 25296 43106 25588
rect 43140 25296 43146 25588
rect 43100 25284 43146 25296
rect 44158 25588 44204 25600
rect 44158 25296 44164 25588
rect 44198 25296 44204 25588
rect 44158 25284 44204 25296
rect 45216 25588 45262 25600
rect 45216 25296 45222 25588
rect 45256 25296 45262 25588
rect 45216 25284 45262 25296
rect 46274 25588 46320 25600
rect 46274 25296 46280 25588
rect 46314 25296 46320 25588
rect 46274 25284 46320 25296
rect 40984 24494 41030 24506
rect 40984 24202 40990 24494
rect 41024 24202 41030 24494
rect 40984 24190 41030 24202
rect 42042 24494 42088 24506
rect 42042 24202 42048 24494
rect 42082 24202 42088 24494
rect 42042 24190 42088 24202
rect 43100 24494 43146 24506
rect 43100 24202 43106 24494
rect 43140 24202 43146 24494
rect 43100 24190 43146 24202
rect 44158 24494 44204 24506
rect 44158 24202 44164 24494
rect 44198 24202 44204 24494
rect 44158 24190 44204 24202
rect 45216 24494 45262 24506
rect 45216 24202 45222 24494
rect 45256 24202 45262 24494
rect 45216 24190 45262 24202
rect 46274 24494 46320 24506
rect 46274 24202 46280 24494
rect 46314 24202 46320 24494
rect 46274 24190 46320 24202
rect 34494 23400 34540 23412
rect 34494 23108 34500 23400
rect 34534 23108 34540 23400
rect 34494 23096 34540 23108
rect 35552 23400 35598 23412
rect 35552 23108 35558 23400
rect 35592 23108 35598 23400
rect 35552 23096 35598 23108
rect 36610 23400 36656 23412
rect 36610 23108 36616 23400
rect 36650 23108 36656 23400
rect 36610 23096 36656 23108
rect 37668 23400 37714 23412
rect 37668 23108 37674 23400
rect 37708 23108 37714 23400
rect 37668 23096 37714 23108
rect 38726 23400 38772 23412
rect 38726 23108 38732 23400
rect 38766 23108 38772 23400
rect 38726 23096 38772 23108
rect 39784 23400 39830 23412
rect 39784 23108 39790 23400
rect 39824 23108 39830 23400
rect 39784 23096 39830 23108
rect 33846 22534 34144 22858
rect 27984 22300 28030 22312
rect 27984 22008 27990 22300
rect 28024 22008 28030 22300
rect 27984 21996 28030 22008
rect 29042 22300 29088 22312
rect 29042 22008 29048 22300
rect 29082 22008 29088 22300
rect 29042 21996 29088 22008
rect 30100 22300 30146 22312
rect 30100 22008 30106 22300
rect 30140 22008 30146 22300
rect 30100 21996 30146 22008
rect 31158 22300 31204 22312
rect 31158 22008 31164 22300
rect 31198 22008 31204 22300
rect 31158 21996 31204 22008
rect 32216 22300 32262 22312
rect 32216 22008 32222 22300
rect 32256 22008 32262 22300
rect 32216 21996 32262 22008
rect 33274 22300 33320 22312
rect 33274 22008 33280 22300
rect 33314 22008 33320 22300
rect 33274 21996 33320 22008
rect 27984 21206 28030 21218
rect 27984 20914 27990 21206
rect 28024 20914 28030 21206
rect 27984 20902 28030 20914
rect 29042 21206 29088 21218
rect 29042 20914 29048 21206
rect 29082 20914 29088 21206
rect 29042 20902 29088 20914
rect 30100 21206 30146 21218
rect 30100 20914 30106 21206
rect 30140 20914 30146 21206
rect 30100 20902 30146 20914
rect 31158 21206 31204 21218
rect 31158 20914 31164 21206
rect 31198 20914 31204 21206
rect 31158 20902 31204 20914
rect 32216 21206 32262 21218
rect 32216 20914 32222 21206
rect 32256 20914 32262 21206
rect 32216 20902 32262 20914
rect 33274 21206 33320 21218
rect 33274 20914 33280 21206
rect 33314 20914 33320 21206
rect 33274 20902 33320 20914
rect 27984 19718 28030 19730
rect 27984 19426 27990 19718
rect 28024 19426 28030 19718
rect 27984 19414 28030 19426
rect 29042 19718 29088 19730
rect 29042 19426 29048 19718
rect 29082 19426 29088 19718
rect 29042 19414 29088 19426
rect 30100 19718 30146 19730
rect 30100 19426 30106 19718
rect 30140 19426 30146 19718
rect 30100 19414 30146 19426
rect 31158 19718 31204 19730
rect 31158 19426 31164 19718
rect 31198 19426 31204 19718
rect 31158 19414 31204 19426
rect 32216 19718 32262 19730
rect 32216 19426 32222 19718
rect 32256 19426 32262 19718
rect 32216 19414 32262 19426
rect 33274 19718 33320 19730
rect 33274 19426 33280 19718
rect 33314 19426 33320 19718
rect 33274 19414 33320 19426
rect 27984 18624 28030 18636
rect 27984 18332 27990 18624
rect 28024 18332 28030 18624
rect 27984 18320 28030 18332
rect 29042 18624 29088 18636
rect 29042 18332 29048 18624
rect 29082 18332 29088 18624
rect 29042 18320 29088 18332
rect 30100 18624 30146 18636
rect 30100 18332 30106 18624
rect 30140 18332 30146 18624
rect 30100 18320 30146 18332
rect 31158 18624 31204 18636
rect 31158 18332 31164 18624
rect 31198 18332 31204 18624
rect 31158 18320 31204 18332
rect 32216 18624 32262 18636
rect 32216 18332 32222 18624
rect 32256 18332 32262 18624
rect 32216 18320 32262 18332
rect 33274 18624 33320 18636
rect 33274 18332 33280 18624
rect 33314 18332 33320 18624
rect 33274 18320 33320 18332
rect 33848 18316 34144 22534
rect 40304 22858 40358 24054
rect 40452 22858 40638 24054
rect 46836 24076 47170 28716
rect 53438 28730 53460 29926
rect 53554 28730 53776 29926
rect 59586 29896 60030 30090
rect 54086 29272 54132 29284
rect 54086 28980 54092 29272
rect 54126 28980 54132 29272
rect 54086 28968 54132 28980
rect 55144 29272 55190 29284
rect 55144 28980 55150 29272
rect 55184 28980 55190 29272
rect 55144 28968 55190 28980
rect 56202 29272 56248 29284
rect 56202 28980 56208 29272
rect 56242 28980 56248 29272
rect 56202 28968 56248 28980
rect 57260 29272 57306 29284
rect 57260 28980 57266 29272
rect 57300 28980 57306 29272
rect 57260 28968 57306 28980
rect 58318 29272 58364 29284
rect 58318 28980 58324 29272
rect 58358 28980 58364 29272
rect 58318 28968 58364 28980
rect 59376 29272 59422 29284
rect 59376 28980 59382 29272
rect 59416 28980 59422 29272
rect 59376 28968 59422 28980
rect 53438 28406 53776 28730
rect 47572 28164 47618 28176
rect 47572 27872 47578 28164
rect 47612 27872 47618 28164
rect 47572 27860 47618 27872
rect 48630 28164 48676 28176
rect 48630 27872 48636 28164
rect 48670 27872 48676 28164
rect 48630 27860 48676 27872
rect 49688 28164 49734 28176
rect 49688 27872 49694 28164
rect 49728 27872 49734 28164
rect 49688 27860 49734 27872
rect 50746 28164 50792 28176
rect 50746 27872 50752 28164
rect 50786 27872 50792 28164
rect 50746 27860 50792 27872
rect 51804 28164 51850 28176
rect 51804 27872 51810 28164
rect 51844 27872 51850 28164
rect 51804 27860 51850 27872
rect 52862 28164 52908 28176
rect 52862 27872 52868 28164
rect 52902 27872 52908 28164
rect 52862 27860 52908 27872
rect 47572 27070 47618 27082
rect 47572 26778 47578 27070
rect 47612 26778 47618 27070
rect 47572 26766 47618 26778
rect 48630 27070 48676 27082
rect 48630 26778 48636 27070
rect 48670 26778 48676 27070
rect 48630 26766 48676 26778
rect 49688 27070 49734 27082
rect 49688 26778 49694 27070
rect 49728 26778 49734 27070
rect 49688 26766 49734 26778
rect 50746 27070 50792 27082
rect 50746 26778 50752 27070
rect 50786 26778 50792 27070
rect 50746 26766 50792 26778
rect 51804 27070 51850 27082
rect 51804 26778 51810 27070
rect 51844 26778 51850 27070
rect 51804 26766 51850 26778
rect 52862 27070 52908 27082
rect 52862 26778 52868 27070
rect 52902 26778 52908 27070
rect 52862 26766 52908 26778
rect 47572 25610 47618 25622
rect 47572 25318 47578 25610
rect 47612 25318 47618 25610
rect 47572 25306 47618 25318
rect 48630 25610 48676 25622
rect 48630 25318 48636 25610
rect 48670 25318 48676 25610
rect 48630 25306 48676 25318
rect 49688 25610 49734 25622
rect 49688 25318 49694 25610
rect 49728 25318 49734 25610
rect 49688 25306 49734 25318
rect 50746 25610 50792 25622
rect 50746 25318 50752 25610
rect 50786 25318 50792 25610
rect 50746 25306 50792 25318
rect 51804 25610 51850 25622
rect 51804 25318 51810 25610
rect 51844 25318 51850 25610
rect 51804 25306 51850 25318
rect 52862 25610 52908 25622
rect 52862 25318 52868 25610
rect 52902 25318 52908 25610
rect 52862 25306 52908 25318
rect 47572 24516 47618 24528
rect 47572 24224 47578 24516
rect 47612 24224 47618 24516
rect 47572 24212 47618 24224
rect 48630 24516 48676 24528
rect 48630 24224 48636 24516
rect 48670 24224 48676 24516
rect 48630 24212 48676 24224
rect 49688 24516 49734 24528
rect 49688 24224 49694 24516
rect 49728 24224 49734 24516
rect 49688 24212 49734 24224
rect 50746 24516 50792 24528
rect 50746 24224 50752 24516
rect 50786 24224 50792 24516
rect 50746 24212 50792 24224
rect 51804 24516 51850 24528
rect 51804 24224 51810 24516
rect 51844 24224 51850 24516
rect 51804 24212 51850 24224
rect 52862 24516 52908 24528
rect 52862 24224 52868 24516
rect 52902 24224 52908 24516
rect 52862 24212 52908 24224
rect 53442 24216 53776 28406
rect 59586 28426 59642 29896
rect 59974 28426 60030 29896
rect 54086 28178 54132 28190
rect 54086 27886 54092 28178
rect 54126 27886 54132 28178
rect 54086 27874 54132 27886
rect 55144 28178 55190 28190
rect 55144 27886 55150 28178
rect 55184 27886 55190 28178
rect 55144 27874 55190 27886
rect 56202 28178 56248 28190
rect 56202 27886 56208 28178
rect 56242 27886 56248 28178
rect 56202 27874 56248 27886
rect 57260 28178 57306 28190
rect 57260 27886 57266 28178
rect 57300 27886 57306 28178
rect 57260 27874 57306 27886
rect 58318 28178 58364 28190
rect 58318 27886 58324 28178
rect 58358 27886 58364 28178
rect 58318 27874 58364 27886
rect 59376 28178 59422 28190
rect 59376 27886 59382 28178
rect 59416 27886 59422 28178
rect 59586 28134 60030 28426
rect 59376 27874 59422 27886
rect 54086 27084 54132 27096
rect 54086 26792 54092 27084
rect 54126 26792 54132 27084
rect 54086 26780 54132 26792
rect 55144 27084 55190 27096
rect 55144 26792 55150 27084
rect 55184 26792 55190 27084
rect 55144 26780 55190 26792
rect 56202 27084 56248 27096
rect 56202 26792 56208 27084
rect 56242 26792 56248 27084
rect 56202 26780 56248 26792
rect 57260 27084 57306 27096
rect 57260 26792 57266 27084
rect 57300 26792 57306 27084
rect 57260 26780 57306 26792
rect 58318 27084 58364 27096
rect 58318 26792 58324 27084
rect 58358 26792 58364 27084
rect 58318 26780 58364 26792
rect 59376 27084 59422 27096
rect 59376 26792 59382 27084
rect 59416 26792 59422 27084
rect 59376 26780 59422 26792
rect 54086 25624 54132 25636
rect 54086 25332 54092 25624
rect 54126 25332 54132 25624
rect 54086 25320 54132 25332
rect 55144 25624 55190 25636
rect 55144 25332 55150 25624
rect 55184 25332 55190 25624
rect 55144 25320 55190 25332
rect 56202 25624 56248 25636
rect 56202 25332 56208 25624
rect 56242 25332 56248 25624
rect 56202 25320 56248 25332
rect 57260 25624 57306 25636
rect 57260 25332 57266 25624
rect 57300 25332 57306 25624
rect 57260 25320 57306 25332
rect 58318 25624 58364 25636
rect 58318 25332 58324 25624
rect 58358 25332 58364 25624
rect 58318 25320 58364 25332
rect 59376 25624 59422 25636
rect 59376 25332 59382 25624
rect 59416 25332 59422 25624
rect 59376 25320 59422 25332
rect 54086 24530 54132 24542
rect 54086 24238 54092 24530
rect 54126 24238 54132 24530
rect 54086 24226 54132 24238
rect 55144 24530 55190 24542
rect 55144 24238 55150 24530
rect 55184 24238 55190 24530
rect 55144 24226 55190 24238
rect 56202 24530 56248 24542
rect 56202 24238 56208 24530
rect 56242 24238 56248 24530
rect 56202 24226 56248 24238
rect 57260 24530 57306 24542
rect 57260 24238 57266 24530
rect 57300 24238 57306 24530
rect 57260 24226 57306 24238
rect 58318 24530 58364 24542
rect 58318 24238 58324 24530
rect 58358 24238 58364 24530
rect 58318 24226 58364 24238
rect 59376 24530 59422 24542
rect 59376 24238 59382 24530
rect 59416 24238 59422 24530
rect 59680 24514 60012 28134
rect 67546 26314 68312 26348
rect 67546 26216 67700 26314
rect 68180 26216 68312 26314
rect 67546 26160 68312 26216
rect 93948 26270 94478 26316
rect 93948 26190 94062 26270
rect 94392 26190 94478 26270
rect 93948 26134 94478 26190
rect 62106 25568 62152 25580
rect 62106 25276 62112 25568
rect 62146 25276 62152 25568
rect 62106 25264 62152 25276
rect 63164 25568 63210 25580
rect 63164 25276 63170 25568
rect 63204 25276 63210 25568
rect 63164 25264 63210 25276
rect 64222 25568 64268 25580
rect 64222 25276 64228 25568
rect 64262 25276 64268 25568
rect 64222 25264 64268 25276
rect 65280 25568 65326 25580
rect 65280 25276 65286 25568
rect 65320 25276 65326 25568
rect 65280 25264 65326 25276
rect 66338 25568 66384 25580
rect 66338 25276 66344 25568
rect 66378 25276 66384 25568
rect 66338 25264 66384 25276
rect 67396 25568 67442 25580
rect 67396 25276 67402 25568
rect 67436 25276 67442 25568
rect 67396 25264 67442 25276
rect 68568 25566 68614 25578
rect 68568 25274 68574 25566
rect 68608 25274 68614 25566
rect 68568 25262 68614 25274
rect 69626 25566 69672 25578
rect 69626 25274 69632 25566
rect 69666 25274 69672 25566
rect 69626 25262 69672 25274
rect 70684 25566 70730 25578
rect 70684 25274 70690 25566
rect 70724 25274 70730 25566
rect 70684 25262 70730 25274
rect 71742 25566 71788 25578
rect 71742 25274 71748 25566
rect 71782 25274 71788 25566
rect 71742 25262 71788 25274
rect 72800 25566 72846 25578
rect 72800 25274 72806 25566
rect 72840 25274 72846 25566
rect 72800 25262 72846 25274
rect 73858 25566 73904 25578
rect 73858 25274 73864 25566
rect 73898 25274 73904 25566
rect 73858 25262 73904 25274
rect 75262 25540 75308 25552
rect 75262 25248 75268 25540
rect 75302 25248 75308 25540
rect 75262 25236 75308 25248
rect 76320 25540 76366 25552
rect 76320 25248 76326 25540
rect 76360 25248 76366 25540
rect 76320 25236 76366 25248
rect 77378 25540 77424 25552
rect 77378 25248 77384 25540
rect 77418 25248 77424 25540
rect 77378 25236 77424 25248
rect 78436 25540 78482 25552
rect 78436 25248 78442 25540
rect 78476 25248 78482 25540
rect 78436 25236 78482 25248
rect 79494 25540 79540 25552
rect 79494 25248 79500 25540
rect 79534 25248 79540 25540
rect 79494 25236 79540 25248
rect 80552 25540 80598 25552
rect 80552 25248 80558 25540
rect 80592 25248 80598 25540
rect 80552 25236 80598 25248
rect 81724 25538 81770 25550
rect 81724 25246 81730 25538
rect 81764 25246 81770 25538
rect 81724 25234 81770 25246
rect 82782 25538 82828 25550
rect 82782 25246 82788 25538
rect 82822 25246 82828 25538
rect 82782 25234 82828 25246
rect 83840 25538 83886 25550
rect 83840 25246 83846 25538
rect 83880 25246 83886 25538
rect 83840 25234 83886 25246
rect 84898 25538 84944 25550
rect 84898 25246 84904 25538
rect 84938 25246 84944 25538
rect 84898 25234 84944 25246
rect 85956 25538 86002 25550
rect 85956 25246 85962 25538
rect 85996 25246 86002 25538
rect 85956 25234 86002 25246
rect 87014 25538 87060 25550
rect 87014 25246 87020 25538
rect 87054 25246 87060 25538
rect 87014 25234 87060 25246
rect 88496 25532 88542 25544
rect 88496 25240 88502 25532
rect 88536 25240 88542 25532
rect 88496 25228 88542 25240
rect 89554 25532 89600 25544
rect 89554 25240 89560 25532
rect 89594 25240 89600 25532
rect 89554 25228 89600 25240
rect 90612 25532 90658 25544
rect 90612 25240 90618 25532
rect 90652 25240 90658 25532
rect 90612 25228 90658 25240
rect 91670 25532 91716 25544
rect 91670 25240 91676 25532
rect 91710 25240 91716 25532
rect 91670 25228 91716 25240
rect 92728 25532 92774 25544
rect 92728 25240 92734 25532
rect 92768 25240 92774 25532
rect 92728 25228 92774 25240
rect 93786 25532 93832 25544
rect 93786 25240 93792 25532
rect 93826 25240 93832 25532
rect 93786 25228 93832 25240
rect 94958 25530 95004 25542
rect 94958 25238 94964 25530
rect 94998 25238 95004 25530
rect 94958 25226 95004 25238
rect 96016 25530 96062 25542
rect 96016 25238 96022 25530
rect 96056 25238 96062 25530
rect 96016 25226 96062 25238
rect 97074 25530 97120 25542
rect 97074 25238 97080 25530
rect 97114 25238 97120 25530
rect 97074 25226 97120 25238
rect 98132 25530 98178 25542
rect 98132 25238 98138 25530
rect 98172 25238 98178 25530
rect 98132 25226 98178 25238
rect 99190 25530 99236 25542
rect 99190 25238 99196 25530
rect 99230 25238 99236 25530
rect 99190 25226 99236 25238
rect 100248 25530 100294 25542
rect 100248 25238 100254 25530
rect 100288 25238 100294 25530
rect 100248 25226 100294 25238
rect 59376 24226 59422 24238
rect 59572 24250 60012 24514
rect 100676 25032 101320 25566
rect 40984 23400 41030 23412
rect 40984 23108 40990 23400
rect 41024 23108 41030 23400
rect 40984 23096 41030 23108
rect 42042 23400 42088 23412
rect 42042 23108 42048 23400
rect 42082 23108 42088 23400
rect 42042 23096 42088 23108
rect 43100 23400 43146 23412
rect 43100 23108 43106 23400
rect 43140 23108 43146 23400
rect 43100 23096 43146 23108
rect 44158 23400 44204 23412
rect 44158 23108 44164 23400
rect 44198 23108 44204 23400
rect 44158 23096 44204 23108
rect 45216 23400 45262 23412
rect 45216 23108 45222 23400
rect 45256 23108 45262 23400
rect 45216 23096 45262 23108
rect 46274 23400 46320 23412
rect 46274 23108 46280 23400
rect 46314 23108 46320 23400
rect 46274 23096 46320 23108
rect 34494 22306 34540 22318
rect 34494 22014 34500 22306
rect 34534 22014 34540 22306
rect 34494 22002 34540 22014
rect 35552 22306 35598 22318
rect 35552 22014 35558 22306
rect 35592 22014 35598 22306
rect 35552 22002 35598 22014
rect 36610 22306 36656 22318
rect 36610 22014 36616 22306
rect 36650 22014 36656 22306
rect 36610 22002 36656 22014
rect 37668 22306 37714 22318
rect 37668 22014 37674 22306
rect 37708 22014 37714 22306
rect 37668 22002 37714 22014
rect 38726 22306 38772 22318
rect 38726 22014 38732 22306
rect 38766 22014 38772 22306
rect 38726 22002 38772 22014
rect 39784 22306 39830 22318
rect 39784 22014 39790 22306
rect 39824 22014 39830 22306
rect 39784 22002 39830 22014
rect 34494 21212 34540 21224
rect 34494 20920 34500 21212
rect 34534 20920 34540 21212
rect 34494 20908 34540 20920
rect 35552 21212 35598 21224
rect 35552 20920 35558 21212
rect 35592 20920 35598 21212
rect 35552 20908 35598 20920
rect 36610 21212 36656 21224
rect 36610 20920 36616 21212
rect 36650 20920 36656 21212
rect 36610 20908 36656 20920
rect 37668 21212 37714 21224
rect 37668 20920 37674 21212
rect 37708 20920 37714 21212
rect 37668 20908 37714 20920
rect 38726 21212 38772 21224
rect 38726 20920 38732 21212
rect 38766 20920 38772 21212
rect 38726 20908 38772 20920
rect 39784 21212 39830 21224
rect 39784 20920 39790 21212
rect 39824 20920 39830 21212
rect 39784 20908 39830 20920
rect 34494 19724 34540 19736
rect 34494 19432 34500 19724
rect 34534 19432 34540 19724
rect 34494 19420 34540 19432
rect 35552 19724 35598 19736
rect 35552 19432 35558 19724
rect 35592 19432 35598 19724
rect 35552 19420 35598 19432
rect 36610 19724 36656 19736
rect 36610 19432 36616 19724
rect 36650 19432 36656 19724
rect 36610 19420 36656 19432
rect 37668 19724 37714 19736
rect 37668 19432 37674 19724
rect 37708 19432 37714 19724
rect 37668 19420 37714 19432
rect 38726 19724 38772 19736
rect 38726 19432 38732 19724
rect 38766 19432 38772 19724
rect 38726 19420 38772 19432
rect 39784 19724 39830 19736
rect 39784 19432 39790 19724
rect 39824 19432 39830 19724
rect 39784 19420 39830 19432
rect 34494 18630 34540 18642
rect 34494 18338 34500 18630
rect 34534 18338 34540 18630
rect 34494 18326 34540 18338
rect 35552 18630 35598 18642
rect 35552 18338 35558 18630
rect 35592 18338 35598 18630
rect 35552 18326 35598 18338
rect 36610 18630 36656 18642
rect 36610 18338 36616 18630
rect 36650 18338 36656 18630
rect 36610 18326 36656 18338
rect 37668 18630 37714 18642
rect 37668 18338 37674 18630
rect 37708 18338 37714 18630
rect 37668 18326 37714 18338
rect 38726 18630 38772 18642
rect 38726 18338 38732 18630
rect 38766 18338 38772 18630
rect 38726 18326 38772 18338
rect 39784 18630 39830 18642
rect 39784 18338 39790 18630
rect 39824 18338 39830 18630
rect 39784 18326 39830 18338
rect 21462 17514 21508 17526
rect 21462 17222 21468 17514
rect 21502 17222 21508 17514
rect 21462 17210 21508 17222
rect 22520 17514 22566 17526
rect 22520 17222 22526 17514
rect 22560 17222 22566 17514
rect 22520 17210 22566 17222
rect 23578 17514 23624 17526
rect 23578 17222 23584 17514
rect 23618 17222 23624 17514
rect 23578 17210 23624 17222
rect 24636 17514 24682 17526
rect 24636 17222 24642 17514
rect 24676 17222 24682 17514
rect 24636 17210 24682 17222
rect 25694 17514 25740 17526
rect 25694 17222 25700 17514
rect 25734 17222 25740 17514
rect 25694 17210 25740 17222
rect 26752 17514 26798 17526
rect 26752 17222 26758 17514
rect 26792 17222 26798 17514
rect 26752 17210 26798 17222
rect 14972 16436 15018 16448
rect 14972 16144 14978 16436
rect 15012 16144 15018 16436
rect 14972 16132 15018 16144
rect 16030 16436 16076 16448
rect 16030 16144 16036 16436
rect 16070 16144 16076 16436
rect 16030 16132 16076 16144
rect 17088 16436 17134 16448
rect 17088 16144 17094 16436
rect 17128 16144 17134 16436
rect 17088 16132 17134 16144
rect 18146 16436 18192 16448
rect 18146 16144 18152 16436
rect 18186 16144 18192 16436
rect 18146 16132 18192 16144
rect 19204 16436 19250 16448
rect 19204 16144 19210 16436
rect 19244 16144 19250 16436
rect 19204 16132 19250 16144
rect 20262 16436 20308 16448
rect 20262 16144 20268 16436
rect 20302 16144 20308 16436
rect 20262 16132 20308 16144
rect 14972 15342 15018 15354
rect 14972 15050 14978 15342
rect 15012 15050 15018 15342
rect 14972 15038 15018 15050
rect 16030 15342 16076 15354
rect 16030 15050 16036 15342
rect 16070 15050 16076 15342
rect 16030 15038 16076 15050
rect 17088 15342 17134 15354
rect 17088 15050 17094 15342
rect 17128 15050 17134 15342
rect 17088 15038 17134 15050
rect 18146 15342 18192 15354
rect 18146 15050 18152 15342
rect 18186 15050 18192 15342
rect 18146 15038 18192 15050
rect 19204 15342 19250 15354
rect 19204 15050 19210 15342
rect 19244 15050 19250 15342
rect 19204 15038 19250 15050
rect 20262 15342 20308 15354
rect 20262 15050 20268 15342
rect 20302 15050 20308 15342
rect 20262 15038 20308 15050
rect 14982 13862 15028 13874
rect 14982 13570 14988 13862
rect 15022 13570 15028 13862
rect 14982 13558 15028 13570
rect 16040 13862 16086 13874
rect 16040 13570 16046 13862
rect 16080 13570 16086 13862
rect 16040 13558 16086 13570
rect 17098 13862 17144 13874
rect 17098 13570 17104 13862
rect 17138 13570 17144 13862
rect 17098 13558 17144 13570
rect 18156 13862 18202 13874
rect 18156 13570 18162 13862
rect 18196 13570 18202 13862
rect 18156 13558 18202 13570
rect 19214 13862 19260 13874
rect 19214 13570 19220 13862
rect 19254 13570 19260 13862
rect 19214 13558 19260 13570
rect 20272 13862 20318 13874
rect 20272 13570 20278 13862
rect 20312 13570 20318 13862
rect 20272 13558 20318 13570
rect 14982 12768 15028 12780
rect 14982 12476 14988 12768
rect 15022 12476 15028 12768
rect 14982 12464 15028 12476
rect 16040 12768 16086 12780
rect 16040 12476 16046 12768
rect 16080 12476 16086 12768
rect 16040 12464 16086 12476
rect 17098 12768 17144 12780
rect 17098 12476 17104 12768
rect 17138 12476 17144 12768
rect 17098 12464 17144 12476
rect 18156 12768 18202 12780
rect 18156 12476 18162 12768
rect 18196 12476 18202 12768
rect 18156 12464 18202 12476
rect 19214 12768 19260 12780
rect 19214 12476 19220 12768
rect 19254 12476 19260 12768
rect 19214 12464 19260 12476
rect 20272 12768 20318 12780
rect 20272 12476 20278 12768
rect 20312 12476 20318 12768
rect 20272 12464 20318 12476
rect 8476 11666 8522 11678
rect 8476 11374 8482 11666
rect 8516 11374 8522 11666
rect 8476 11362 8522 11374
rect 9534 11666 9580 11678
rect 9534 11374 9540 11666
rect 9574 11374 9580 11666
rect 9534 11362 9580 11374
rect 10592 11666 10638 11678
rect 10592 11374 10598 11666
rect 10632 11374 10638 11666
rect 10592 11362 10638 11374
rect 11650 11666 11696 11678
rect 11650 11374 11656 11666
rect 11690 11374 11696 11666
rect 11650 11362 11696 11374
rect 12708 11666 12754 11678
rect 12708 11374 12714 11666
rect 12748 11374 12754 11666
rect 12708 11362 12754 11374
rect 13766 11666 13812 11678
rect 13766 11374 13772 11666
rect 13806 11374 13812 11666
rect 13766 11362 13812 11374
rect 1962 10564 2008 10576
rect 1962 10272 1968 10564
rect 2002 10272 2008 10564
rect 1962 10260 2008 10272
rect 3020 10564 3066 10576
rect 3020 10272 3026 10564
rect 3060 10272 3066 10564
rect 3020 10260 3066 10272
rect 4078 10564 4124 10576
rect 4078 10272 4084 10564
rect 4118 10272 4124 10564
rect 4078 10260 4124 10272
rect 5136 10564 5182 10576
rect 5136 10272 5142 10564
rect 5176 10272 5182 10564
rect 5136 10260 5182 10272
rect 6194 10564 6240 10576
rect 6194 10272 6200 10564
rect 6234 10272 6240 10564
rect 6194 10260 6240 10272
rect 7252 10564 7298 10576
rect 7252 10272 7258 10564
rect 7292 10272 7298 10564
rect 7252 10260 7298 10272
rect 1962 9470 2008 9482
rect 1962 9178 1968 9470
rect 2002 9178 2008 9470
rect 1962 9166 2008 9178
rect 3020 9470 3066 9482
rect 3020 9178 3026 9470
rect 3060 9178 3066 9470
rect 3020 9166 3066 9178
rect 4078 9470 4124 9482
rect 4078 9178 4084 9470
rect 4118 9178 4124 9470
rect 4078 9166 4124 9178
rect 5136 9470 5182 9482
rect 5136 9178 5142 9470
rect 5176 9178 5182 9470
rect 5136 9166 5182 9178
rect 6194 9470 6240 9482
rect 6194 9178 6200 9470
rect 6234 9178 6240 9470
rect 6194 9166 6240 9178
rect 7252 9470 7298 9482
rect 7252 9178 7258 9470
rect 7292 9178 7298 9470
rect 7252 9166 7298 9178
rect 1980 7938 2026 7950
rect 1980 7646 1986 7938
rect 2020 7646 2026 7938
rect 1980 7634 2026 7646
rect 3038 7938 3084 7950
rect 3038 7646 3044 7938
rect 3078 7646 3084 7938
rect 3038 7634 3084 7646
rect 4096 7938 4142 7950
rect 4096 7646 4102 7938
rect 4136 7646 4142 7938
rect 4096 7634 4142 7646
rect 5154 7938 5200 7950
rect 5154 7646 5160 7938
rect 5194 7646 5200 7938
rect 5154 7634 5200 7646
rect 6212 7938 6258 7950
rect 6212 7646 6218 7938
rect 6252 7646 6258 7938
rect 6212 7634 6258 7646
rect 7270 7938 7316 7950
rect 7270 7646 7276 7938
rect 7310 7646 7316 7938
rect 7270 7634 7316 7646
rect 1980 6844 2026 6856
rect 1980 6552 1986 6844
rect 2020 6552 2026 6844
rect 1980 6540 2026 6552
rect 3038 6844 3084 6856
rect 3038 6552 3044 6844
rect 3078 6552 3084 6844
rect 3038 6540 3084 6552
rect 4096 6844 4142 6856
rect 4096 6552 4102 6844
rect 4136 6552 4142 6844
rect 4096 6540 4142 6552
rect 5154 6844 5200 6856
rect 5154 6552 5160 6844
rect 5194 6552 5200 6844
rect 5154 6540 5200 6552
rect 6212 6844 6258 6856
rect 6212 6552 6218 6844
rect 6252 6552 6258 6844
rect 6212 6540 6258 6552
rect 7270 6844 7316 6856
rect 7270 6552 7276 6844
rect 7310 6552 7316 6844
rect 7270 6540 7316 6552
rect 1264 5208 1354 6404
rect 1448 5208 1560 6404
rect 7722 6412 8018 11124
rect 14216 11132 14356 12328
rect 14450 11132 14512 12328
rect 20748 12312 21044 16972
rect 27278 16988 27358 18184
rect 27452 16988 27574 18184
rect 33846 18190 34144 18316
rect 27984 17530 28030 17542
rect 27984 17238 27990 17530
rect 28024 17238 28030 17530
rect 27984 17226 28030 17238
rect 29042 17530 29088 17542
rect 29042 17238 29048 17530
rect 29082 17238 29088 17530
rect 29042 17226 29088 17238
rect 30100 17530 30146 17542
rect 30100 17238 30106 17530
rect 30140 17238 30146 17530
rect 30100 17226 30146 17238
rect 31158 17530 31204 17542
rect 31158 17238 31164 17530
rect 31198 17238 31204 17530
rect 31158 17226 31204 17238
rect 32216 17530 32262 17542
rect 32216 17238 32222 17530
rect 32256 17238 32262 17530
rect 32216 17226 32262 17238
rect 33274 17530 33320 17542
rect 33274 17238 33280 17530
rect 33314 17238 33320 17530
rect 33274 17226 33320 17238
rect 21462 16420 21508 16432
rect 21462 16128 21468 16420
rect 21502 16128 21508 16420
rect 21462 16116 21508 16128
rect 22520 16420 22566 16432
rect 22520 16128 22526 16420
rect 22560 16128 22566 16420
rect 22520 16116 22566 16128
rect 23578 16420 23624 16432
rect 23578 16128 23584 16420
rect 23618 16128 23624 16420
rect 23578 16116 23624 16128
rect 24636 16420 24682 16432
rect 24636 16128 24642 16420
rect 24676 16128 24682 16420
rect 24636 16116 24682 16128
rect 25694 16420 25740 16432
rect 25694 16128 25700 16420
rect 25734 16128 25740 16420
rect 25694 16116 25740 16128
rect 26752 16420 26798 16432
rect 26752 16128 26758 16420
rect 26792 16128 26798 16420
rect 26752 16116 26798 16128
rect 21462 15326 21508 15338
rect 21462 15034 21468 15326
rect 21502 15034 21508 15326
rect 21462 15022 21508 15034
rect 22520 15326 22566 15338
rect 22520 15034 22526 15326
rect 22560 15034 22566 15326
rect 22520 15022 22566 15034
rect 23578 15326 23624 15338
rect 23578 15034 23584 15326
rect 23618 15034 23624 15326
rect 23578 15022 23624 15034
rect 24636 15326 24682 15338
rect 24636 15034 24642 15326
rect 24676 15034 24682 15326
rect 24636 15022 24682 15034
rect 25694 15326 25740 15338
rect 25694 15034 25700 15326
rect 25734 15034 25740 15326
rect 25694 15022 25740 15034
rect 26752 15326 26798 15338
rect 26752 15034 26758 15326
rect 26792 15034 26798 15326
rect 26752 15022 26798 15034
rect 21472 13846 21518 13858
rect 21472 13554 21478 13846
rect 21512 13554 21518 13846
rect 21472 13542 21518 13554
rect 22530 13846 22576 13858
rect 22530 13554 22536 13846
rect 22570 13554 22576 13846
rect 22530 13542 22576 13554
rect 23588 13846 23634 13858
rect 23588 13554 23594 13846
rect 23628 13554 23634 13846
rect 23588 13542 23634 13554
rect 24646 13846 24692 13858
rect 24646 13554 24652 13846
rect 24686 13554 24692 13846
rect 24646 13542 24692 13554
rect 25704 13846 25750 13858
rect 25704 13554 25710 13846
rect 25744 13554 25750 13846
rect 25704 13542 25750 13554
rect 26762 13846 26808 13858
rect 26762 13554 26768 13846
rect 26802 13554 26808 13846
rect 26762 13542 26808 13554
rect 21472 12752 21518 12764
rect 21472 12460 21478 12752
rect 21512 12460 21518 12752
rect 21472 12448 21518 12460
rect 22530 12752 22576 12764
rect 22530 12460 22536 12752
rect 22570 12460 22576 12752
rect 22530 12448 22576 12460
rect 23588 12752 23634 12764
rect 23588 12460 23594 12752
rect 23628 12460 23634 12752
rect 23588 12448 23634 12460
rect 24646 12752 24692 12764
rect 24646 12460 24652 12752
rect 24686 12460 24692 12752
rect 24646 12448 24692 12460
rect 25704 12752 25750 12764
rect 25704 12460 25710 12752
rect 25744 12460 25750 12752
rect 25704 12448 25750 12460
rect 26762 12752 26808 12764
rect 26762 12460 26768 12752
rect 26802 12460 26808 12752
rect 26762 12448 26808 12460
rect 14982 11674 15028 11686
rect 14982 11382 14988 11674
rect 15022 11382 15028 11674
rect 14982 11370 15028 11382
rect 16040 11674 16086 11686
rect 16040 11382 16046 11674
rect 16080 11382 16086 11674
rect 16040 11370 16086 11382
rect 17098 11674 17144 11686
rect 17098 11382 17104 11674
rect 17138 11382 17144 11674
rect 17098 11370 17144 11382
rect 18156 11674 18202 11686
rect 18156 11382 18162 11674
rect 18196 11382 18202 11674
rect 18156 11370 18202 11382
rect 19214 11674 19260 11686
rect 19214 11382 19220 11674
rect 19254 11382 19260 11674
rect 19214 11370 19260 11382
rect 20272 11674 20318 11686
rect 20272 11382 20278 11674
rect 20312 11382 20318 11674
rect 20272 11370 20318 11382
rect 8476 10572 8522 10584
rect 8476 10280 8482 10572
rect 8516 10280 8522 10572
rect 8476 10268 8522 10280
rect 9534 10572 9580 10584
rect 9534 10280 9540 10572
rect 9574 10280 9580 10572
rect 9534 10268 9580 10280
rect 10592 10572 10638 10584
rect 10592 10280 10598 10572
rect 10632 10280 10638 10572
rect 10592 10268 10638 10280
rect 11650 10572 11696 10584
rect 11650 10280 11656 10572
rect 11690 10280 11696 10572
rect 11650 10268 11696 10280
rect 12708 10572 12754 10584
rect 12708 10280 12714 10572
rect 12748 10280 12754 10572
rect 12708 10268 12754 10280
rect 13766 10572 13812 10584
rect 13766 10280 13772 10572
rect 13806 10280 13812 10572
rect 13766 10268 13812 10280
rect 8476 9478 8522 9490
rect 8476 9186 8482 9478
rect 8516 9186 8522 9478
rect 8476 9174 8522 9186
rect 9534 9478 9580 9490
rect 9534 9186 9540 9478
rect 9574 9186 9580 9478
rect 9534 9174 9580 9186
rect 10592 9478 10638 9490
rect 10592 9186 10598 9478
rect 10632 9186 10638 9478
rect 10592 9174 10638 9186
rect 11650 9478 11696 9490
rect 11650 9186 11656 9478
rect 11690 9186 11696 9478
rect 11650 9174 11696 9186
rect 12708 9478 12754 9490
rect 12708 9186 12714 9478
rect 12748 9186 12754 9478
rect 12708 9174 12754 9186
rect 13766 9478 13812 9490
rect 13766 9186 13772 9478
rect 13806 9186 13812 9478
rect 13766 9174 13812 9186
rect 8494 7946 8540 7958
rect 8494 7654 8500 7946
rect 8534 7654 8540 7946
rect 8494 7642 8540 7654
rect 9552 7946 9598 7958
rect 9552 7654 9558 7946
rect 9592 7654 9598 7946
rect 9552 7642 9598 7654
rect 10610 7946 10656 7958
rect 10610 7654 10616 7946
rect 10650 7654 10656 7946
rect 10610 7642 10656 7654
rect 11668 7946 11714 7958
rect 11668 7654 11674 7946
rect 11708 7654 11714 7946
rect 11668 7642 11714 7654
rect 12726 7946 12772 7958
rect 12726 7654 12732 7946
rect 12766 7654 12772 7946
rect 12726 7642 12772 7654
rect 13784 7946 13830 7958
rect 13784 7654 13790 7946
rect 13824 7654 13830 7946
rect 13784 7642 13830 7654
rect 8494 6852 8540 6864
rect 8494 6560 8500 6852
rect 8534 6560 8540 6852
rect 8494 6548 8540 6560
rect 9552 6852 9598 6864
rect 9552 6560 9558 6852
rect 9592 6560 9598 6852
rect 9552 6548 9598 6560
rect 10610 6852 10656 6864
rect 10610 6560 10616 6852
rect 10650 6560 10656 6852
rect 10610 6548 10656 6560
rect 11668 6852 11714 6864
rect 11668 6560 11674 6852
rect 11708 6560 11714 6852
rect 11668 6548 11714 6560
rect 12726 6852 12772 6864
rect 12726 6560 12732 6852
rect 12766 6560 12772 6852
rect 12726 6548 12772 6560
rect 13784 6852 13830 6864
rect 13784 6560 13790 6852
rect 13824 6560 13830 6852
rect 13784 6548 13830 6560
rect 1980 5750 2026 5762
rect 1980 5458 1986 5750
rect 2020 5458 2026 5750
rect 1980 5446 2026 5458
rect 3038 5750 3084 5762
rect 3038 5458 3044 5750
rect 3078 5458 3084 5750
rect 3038 5446 3084 5458
rect 4096 5750 4142 5762
rect 4096 5458 4102 5750
rect 4136 5458 4142 5750
rect 4096 5446 4142 5458
rect 5154 5750 5200 5762
rect 5154 5458 5160 5750
rect 5194 5458 5200 5750
rect 5154 5446 5200 5458
rect 6212 5750 6258 5762
rect 6212 5458 6218 5750
rect 6252 5458 6258 5750
rect 6212 5446 6258 5458
rect 7270 5750 7316 5762
rect 7270 5458 7276 5750
rect 7310 5458 7316 5750
rect 7270 5446 7316 5458
rect 1264 -3192 1560 5208
rect 7722 5216 7868 6412
rect 7962 5216 8018 6412
rect 14216 6420 14512 11132
rect 20748 11116 20846 12312
rect 20940 11116 21044 12312
rect 27278 12328 27574 16988
rect 33846 16994 33868 18190
rect 33962 16994 34144 18190
rect 40304 18190 40638 22858
rect 46836 22880 46946 24076
rect 47040 22880 47170 24076
rect 53438 24090 53776 24216
rect 47572 23422 47618 23434
rect 47572 23130 47578 23422
rect 47612 23130 47618 23422
rect 47572 23118 47618 23130
rect 48630 23422 48676 23434
rect 48630 23130 48636 23422
rect 48670 23130 48676 23422
rect 48630 23118 48676 23130
rect 49688 23422 49734 23434
rect 49688 23130 49694 23422
rect 49728 23130 49734 23422
rect 49688 23118 49734 23130
rect 50746 23422 50792 23434
rect 50746 23130 50752 23422
rect 50786 23130 50792 23422
rect 50746 23118 50792 23130
rect 51804 23422 51850 23434
rect 51804 23130 51810 23422
rect 51844 23130 51850 23422
rect 51804 23118 51850 23130
rect 52862 23422 52908 23434
rect 52862 23130 52868 23422
rect 52902 23130 52908 23422
rect 52862 23118 52908 23130
rect 40984 22306 41030 22318
rect 40984 22014 40990 22306
rect 41024 22014 41030 22306
rect 40984 22002 41030 22014
rect 42042 22306 42088 22318
rect 42042 22014 42048 22306
rect 42082 22014 42088 22306
rect 42042 22002 42088 22014
rect 43100 22306 43146 22318
rect 43100 22014 43106 22306
rect 43140 22014 43146 22306
rect 43100 22002 43146 22014
rect 44158 22306 44204 22318
rect 44158 22014 44164 22306
rect 44198 22014 44204 22306
rect 44158 22002 44204 22014
rect 45216 22306 45262 22318
rect 45216 22014 45222 22306
rect 45256 22014 45262 22306
rect 45216 22002 45262 22014
rect 46274 22306 46320 22318
rect 46274 22014 46280 22306
rect 46314 22014 46320 22306
rect 46274 22002 46320 22014
rect 40984 21212 41030 21224
rect 40984 20920 40990 21212
rect 41024 20920 41030 21212
rect 40984 20908 41030 20920
rect 42042 21212 42088 21224
rect 42042 20920 42048 21212
rect 42082 20920 42088 21212
rect 42042 20908 42088 20920
rect 43100 21212 43146 21224
rect 43100 20920 43106 21212
rect 43140 20920 43146 21212
rect 43100 20908 43146 20920
rect 44158 21212 44204 21224
rect 44158 20920 44164 21212
rect 44198 20920 44204 21212
rect 44158 20908 44204 20920
rect 45216 21212 45262 21224
rect 45216 20920 45222 21212
rect 45256 20920 45262 21212
rect 45216 20908 45262 20920
rect 46274 21212 46320 21224
rect 46274 20920 46280 21212
rect 46314 20920 46320 21212
rect 46274 20908 46320 20920
rect 40984 19724 41030 19736
rect 40984 19432 40990 19724
rect 41024 19432 41030 19724
rect 40984 19420 41030 19432
rect 42042 19724 42088 19736
rect 42042 19432 42048 19724
rect 42082 19432 42088 19724
rect 42042 19420 42088 19432
rect 43100 19724 43146 19736
rect 43100 19432 43106 19724
rect 43140 19432 43146 19724
rect 43100 19420 43146 19432
rect 44158 19724 44204 19736
rect 44158 19432 44164 19724
rect 44198 19432 44204 19724
rect 44158 19420 44204 19432
rect 45216 19724 45262 19736
rect 45216 19432 45222 19724
rect 45256 19432 45262 19724
rect 45216 19420 45262 19432
rect 46274 19724 46320 19736
rect 46274 19432 46280 19724
rect 46314 19432 46320 19724
rect 46274 19420 46320 19432
rect 40984 18630 41030 18642
rect 40984 18338 40990 18630
rect 41024 18338 41030 18630
rect 40984 18326 41030 18338
rect 42042 18630 42088 18642
rect 42042 18338 42048 18630
rect 42082 18338 42088 18630
rect 42042 18326 42088 18338
rect 43100 18630 43146 18642
rect 43100 18338 43106 18630
rect 43140 18338 43146 18630
rect 43100 18326 43146 18338
rect 44158 18630 44204 18642
rect 44158 18338 44164 18630
rect 44198 18338 44204 18630
rect 44158 18326 44204 18338
rect 45216 18630 45262 18642
rect 45216 18338 45222 18630
rect 45256 18338 45262 18630
rect 45216 18326 45262 18338
rect 46274 18630 46320 18642
rect 46274 18338 46280 18630
rect 46314 18338 46320 18630
rect 46274 18326 46320 18338
rect 34494 17536 34540 17548
rect 34494 17244 34500 17536
rect 34534 17244 34540 17536
rect 34494 17232 34540 17244
rect 35552 17536 35598 17548
rect 35552 17244 35558 17536
rect 35592 17244 35598 17536
rect 35552 17232 35598 17244
rect 36610 17536 36656 17548
rect 36610 17244 36616 17536
rect 36650 17244 36656 17536
rect 36610 17232 36656 17244
rect 37668 17536 37714 17548
rect 37668 17244 37674 17536
rect 37708 17244 37714 17536
rect 37668 17232 37714 17244
rect 38726 17536 38772 17548
rect 38726 17244 38732 17536
rect 38766 17244 38772 17536
rect 38726 17232 38772 17244
rect 39784 17536 39830 17548
rect 39784 17244 39790 17536
rect 39824 17244 39830 17536
rect 39784 17232 39830 17244
rect 33846 16670 34144 16994
rect 27984 16436 28030 16448
rect 27984 16144 27990 16436
rect 28024 16144 28030 16436
rect 27984 16132 28030 16144
rect 29042 16436 29088 16448
rect 29042 16144 29048 16436
rect 29082 16144 29088 16436
rect 29042 16132 29088 16144
rect 30100 16436 30146 16448
rect 30100 16144 30106 16436
rect 30140 16144 30146 16436
rect 30100 16132 30146 16144
rect 31158 16436 31204 16448
rect 31158 16144 31164 16436
rect 31198 16144 31204 16436
rect 31158 16132 31204 16144
rect 32216 16436 32262 16448
rect 32216 16144 32222 16436
rect 32256 16144 32262 16436
rect 32216 16132 32262 16144
rect 33274 16436 33320 16448
rect 33274 16144 33280 16436
rect 33314 16144 33320 16436
rect 33274 16132 33320 16144
rect 27984 15342 28030 15354
rect 27984 15050 27990 15342
rect 28024 15050 28030 15342
rect 27984 15038 28030 15050
rect 29042 15342 29088 15354
rect 29042 15050 29048 15342
rect 29082 15050 29088 15342
rect 29042 15038 29088 15050
rect 30100 15342 30146 15354
rect 30100 15050 30106 15342
rect 30140 15050 30146 15342
rect 30100 15038 30146 15050
rect 31158 15342 31204 15354
rect 31158 15050 31164 15342
rect 31198 15050 31204 15342
rect 31158 15038 31204 15050
rect 32216 15342 32262 15354
rect 32216 15050 32222 15342
rect 32256 15050 32262 15342
rect 32216 15038 32262 15050
rect 33274 15342 33320 15354
rect 33274 15050 33280 15342
rect 33314 15050 33320 15342
rect 33274 15038 33320 15050
rect 27994 13862 28040 13874
rect 27994 13570 28000 13862
rect 28034 13570 28040 13862
rect 27994 13558 28040 13570
rect 29052 13862 29098 13874
rect 29052 13570 29058 13862
rect 29092 13570 29098 13862
rect 29052 13558 29098 13570
rect 30110 13862 30156 13874
rect 30110 13570 30116 13862
rect 30150 13570 30156 13862
rect 30110 13558 30156 13570
rect 31168 13862 31214 13874
rect 31168 13570 31174 13862
rect 31208 13570 31214 13862
rect 31168 13558 31214 13570
rect 32226 13862 32272 13874
rect 32226 13570 32232 13862
rect 32266 13570 32272 13862
rect 32226 13558 32272 13570
rect 33284 13862 33330 13874
rect 33284 13570 33290 13862
rect 33324 13570 33330 13862
rect 33284 13558 33330 13570
rect 27994 12768 28040 12780
rect 27994 12476 28000 12768
rect 28034 12476 28040 12768
rect 27994 12464 28040 12476
rect 29052 12768 29098 12780
rect 29052 12476 29058 12768
rect 29092 12476 29098 12768
rect 29052 12464 29098 12476
rect 30110 12768 30156 12780
rect 30110 12476 30116 12768
rect 30150 12476 30156 12768
rect 30110 12464 30156 12476
rect 31168 12768 31214 12780
rect 31168 12476 31174 12768
rect 31208 12476 31214 12768
rect 31168 12464 31214 12476
rect 32226 12768 32272 12780
rect 32226 12476 32232 12768
rect 32266 12476 32272 12768
rect 32226 12464 32272 12476
rect 33284 12768 33330 12780
rect 33284 12476 33290 12768
rect 33324 12476 33330 12768
rect 33284 12464 33330 12476
rect 21472 11658 21518 11670
rect 21472 11366 21478 11658
rect 21512 11366 21518 11658
rect 21472 11354 21518 11366
rect 22530 11658 22576 11670
rect 22530 11366 22536 11658
rect 22570 11366 22576 11658
rect 22530 11354 22576 11366
rect 23588 11658 23634 11670
rect 23588 11366 23594 11658
rect 23628 11366 23634 11658
rect 23588 11354 23634 11366
rect 24646 11658 24692 11670
rect 24646 11366 24652 11658
rect 24686 11366 24692 11658
rect 24646 11354 24692 11366
rect 25704 11658 25750 11670
rect 25704 11366 25710 11658
rect 25744 11366 25750 11658
rect 25704 11354 25750 11366
rect 26762 11658 26808 11670
rect 26762 11366 26768 11658
rect 26802 11366 26808 11658
rect 26762 11354 26808 11366
rect 14982 10580 15028 10592
rect 14982 10288 14988 10580
rect 15022 10288 15028 10580
rect 14982 10276 15028 10288
rect 16040 10580 16086 10592
rect 16040 10288 16046 10580
rect 16080 10288 16086 10580
rect 16040 10276 16086 10288
rect 17098 10580 17144 10592
rect 17098 10288 17104 10580
rect 17138 10288 17144 10580
rect 17098 10276 17144 10288
rect 18156 10580 18202 10592
rect 18156 10288 18162 10580
rect 18196 10288 18202 10580
rect 18156 10276 18202 10288
rect 19214 10580 19260 10592
rect 19214 10288 19220 10580
rect 19254 10288 19260 10580
rect 19214 10276 19260 10288
rect 20272 10580 20318 10592
rect 20272 10288 20278 10580
rect 20312 10288 20318 10580
rect 20272 10276 20318 10288
rect 14982 9486 15028 9498
rect 14982 9194 14988 9486
rect 15022 9194 15028 9486
rect 14982 9182 15028 9194
rect 16040 9486 16086 9498
rect 16040 9194 16046 9486
rect 16080 9194 16086 9486
rect 16040 9182 16086 9194
rect 17098 9486 17144 9498
rect 17098 9194 17104 9486
rect 17138 9194 17144 9486
rect 17098 9182 17144 9194
rect 18156 9486 18202 9498
rect 18156 9194 18162 9486
rect 18196 9194 18202 9486
rect 18156 9182 18202 9194
rect 19214 9486 19260 9498
rect 19214 9194 19220 9486
rect 19254 9194 19260 9486
rect 19214 9182 19260 9194
rect 20272 9486 20318 9498
rect 20272 9194 20278 9486
rect 20312 9194 20318 9486
rect 20272 9182 20318 9194
rect 15000 7954 15046 7966
rect 15000 7662 15006 7954
rect 15040 7662 15046 7954
rect 15000 7650 15046 7662
rect 16058 7954 16104 7966
rect 16058 7662 16064 7954
rect 16098 7662 16104 7954
rect 16058 7650 16104 7662
rect 17116 7954 17162 7966
rect 17116 7662 17122 7954
rect 17156 7662 17162 7954
rect 17116 7650 17162 7662
rect 18174 7954 18220 7966
rect 18174 7662 18180 7954
rect 18214 7662 18220 7954
rect 18174 7650 18220 7662
rect 19232 7954 19278 7966
rect 19232 7662 19238 7954
rect 19272 7662 19278 7954
rect 19232 7650 19278 7662
rect 20290 7954 20336 7966
rect 20290 7662 20296 7954
rect 20330 7662 20336 7954
rect 20290 7650 20336 7662
rect 15000 6860 15046 6872
rect 15000 6568 15006 6860
rect 15040 6568 15046 6860
rect 15000 6556 15046 6568
rect 16058 6860 16104 6872
rect 16058 6568 16064 6860
rect 16098 6568 16104 6860
rect 16058 6556 16104 6568
rect 17116 6860 17162 6872
rect 17116 6568 17122 6860
rect 17156 6568 17162 6860
rect 17116 6556 17162 6568
rect 18174 6860 18220 6872
rect 18174 6568 18180 6860
rect 18214 6568 18220 6860
rect 18174 6556 18220 6568
rect 19232 6860 19278 6872
rect 19232 6568 19238 6860
rect 19272 6568 19278 6860
rect 19232 6556 19278 6568
rect 20290 6860 20336 6872
rect 20290 6568 20296 6860
rect 20330 6568 20336 6860
rect 20290 6556 20336 6568
rect 8494 5758 8540 5770
rect 8494 5466 8500 5758
rect 8534 5466 8540 5758
rect 8494 5454 8540 5466
rect 9552 5758 9598 5770
rect 9552 5466 9558 5758
rect 9592 5466 9598 5758
rect 9552 5454 9598 5466
rect 10610 5758 10656 5770
rect 10610 5466 10616 5758
rect 10650 5466 10656 5758
rect 10610 5454 10656 5466
rect 11668 5758 11714 5770
rect 11668 5466 11674 5758
rect 11708 5466 11714 5758
rect 11668 5454 11714 5466
rect 12726 5758 12772 5770
rect 12726 5466 12732 5758
rect 12766 5466 12772 5758
rect 12726 5454 12772 5466
rect 13784 5758 13830 5770
rect 13784 5466 13790 5758
rect 13824 5466 13830 5758
rect 13784 5454 13830 5466
rect 1980 4656 2026 4668
rect 1980 4364 1986 4656
rect 2020 4364 2026 4656
rect 1980 4352 2026 4364
rect 3038 4656 3084 4668
rect 3038 4364 3044 4656
rect 3078 4364 3084 4656
rect 3038 4352 3084 4364
rect 4096 4656 4142 4668
rect 4096 4364 4102 4656
rect 4136 4364 4142 4656
rect 4096 4352 4142 4364
rect 5154 4656 5200 4668
rect 5154 4364 5160 4656
rect 5194 4364 5200 4656
rect 5154 4352 5200 4364
rect 6212 4656 6258 4668
rect 6212 4364 6218 4656
rect 6252 4364 6258 4656
rect 6212 4352 6258 4364
rect 7270 4656 7316 4668
rect 7270 4364 7276 4656
rect 7310 4364 7316 4656
rect 7270 4352 7316 4364
rect 1980 3562 2026 3574
rect 1980 3270 1986 3562
rect 2020 3270 2026 3562
rect 1980 3258 2026 3270
rect 3038 3562 3084 3574
rect 3038 3270 3044 3562
rect 3078 3270 3084 3562
rect 3038 3258 3084 3270
rect 4096 3562 4142 3574
rect 4096 3270 4102 3562
rect 4136 3270 4142 3562
rect 4096 3258 4142 3270
rect 5154 3562 5200 3574
rect 5154 3270 5160 3562
rect 5194 3270 5200 3562
rect 5154 3258 5200 3270
rect 6212 3562 6258 3574
rect 6212 3270 6218 3562
rect 6252 3270 6258 3562
rect 6212 3258 6258 3270
rect 7270 3562 7316 3574
rect 7270 3270 7276 3562
rect 7310 3270 7316 3562
rect 7270 3258 7316 3270
rect 7722 -3192 8018 5216
rect 14216 5224 14374 6420
rect 14468 5224 14512 6420
rect 20748 6404 21044 11116
rect 27278 11132 27368 12328
rect 27462 11132 27574 12328
rect 33848 12334 34144 16670
rect 40304 16994 40358 18190
rect 40452 16994 40638 18190
rect 46836 18212 47170 22880
rect 53438 22894 53460 24090
rect 53554 22894 53776 24090
rect 54086 23436 54132 23448
rect 54086 23144 54092 23436
rect 54126 23144 54132 23436
rect 54086 23132 54132 23144
rect 55144 23436 55190 23448
rect 55144 23144 55150 23436
rect 55184 23144 55190 23436
rect 55144 23132 55190 23144
rect 56202 23436 56248 23448
rect 56202 23144 56208 23436
rect 56242 23144 56248 23436
rect 56202 23132 56248 23144
rect 57260 23436 57306 23448
rect 57260 23144 57266 23436
rect 57300 23144 57306 23436
rect 57260 23132 57306 23144
rect 58318 23436 58364 23448
rect 58318 23144 58324 23436
rect 58358 23144 58364 23436
rect 58318 23132 58364 23144
rect 59376 23436 59422 23448
rect 59376 23144 59382 23436
rect 59416 23144 59422 23436
rect 59376 23132 59422 23144
rect 53438 22570 53776 22894
rect 47572 22328 47618 22340
rect 47572 22036 47578 22328
rect 47612 22036 47618 22328
rect 47572 22024 47618 22036
rect 48630 22328 48676 22340
rect 48630 22036 48636 22328
rect 48670 22036 48676 22328
rect 48630 22024 48676 22036
rect 49688 22328 49734 22340
rect 49688 22036 49694 22328
rect 49728 22036 49734 22328
rect 49688 22024 49734 22036
rect 50746 22328 50792 22340
rect 50746 22036 50752 22328
rect 50786 22036 50792 22328
rect 50746 22024 50792 22036
rect 51804 22328 51850 22340
rect 51804 22036 51810 22328
rect 51844 22036 51850 22328
rect 51804 22024 51850 22036
rect 52862 22328 52908 22340
rect 52862 22036 52868 22328
rect 52902 22036 52908 22328
rect 52862 22024 52908 22036
rect 47572 21234 47618 21246
rect 47572 20942 47578 21234
rect 47612 20942 47618 21234
rect 47572 20930 47618 20942
rect 48630 21234 48676 21246
rect 48630 20942 48636 21234
rect 48670 20942 48676 21234
rect 48630 20930 48676 20942
rect 49688 21234 49734 21246
rect 49688 20942 49694 21234
rect 49728 20942 49734 21234
rect 49688 20930 49734 20942
rect 50746 21234 50792 21246
rect 50746 20942 50752 21234
rect 50786 20942 50792 21234
rect 50746 20930 50792 20942
rect 51804 21234 51850 21246
rect 51804 20942 51810 21234
rect 51844 20942 51850 21234
rect 51804 20930 51850 20942
rect 52862 21234 52908 21246
rect 52862 20942 52868 21234
rect 52902 20942 52908 21234
rect 52862 20930 52908 20942
rect 47572 19746 47618 19758
rect 47572 19454 47578 19746
rect 47612 19454 47618 19746
rect 47572 19442 47618 19454
rect 48630 19746 48676 19758
rect 48630 19454 48636 19746
rect 48670 19454 48676 19746
rect 48630 19442 48676 19454
rect 49688 19746 49734 19758
rect 49688 19454 49694 19746
rect 49728 19454 49734 19746
rect 49688 19442 49734 19454
rect 50746 19746 50792 19758
rect 50746 19454 50752 19746
rect 50786 19454 50792 19746
rect 50746 19442 50792 19454
rect 51804 19746 51850 19758
rect 51804 19454 51810 19746
rect 51844 19454 51850 19746
rect 51804 19442 51850 19454
rect 52862 19746 52908 19758
rect 52862 19454 52868 19746
rect 52902 19454 52908 19746
rect 52862 19442 52908 19454
rect 47572 18652 47618 18664
rect 47572 18360 47578 18652
rect 47612 18360 47618 18652
rect 47572 18348 47618 18360
rect 48630 18652 48676 18664
rect 48630 18360 48636 18652
rect 48670 18360 48676 18652
rect 48630 18348 48676 18360
rect 49688 18652 49734 18664
rect 49688 18360 49694 18652
rect 49728 18360 49734 18652
rect 49688 18348 49734 18360
rect 50746 18652 50792 18664
rect 50746 18360 50752 18652
rect 50786 18360 50792 18652
rect 50746 18348 50792 18360
rect 51804 18652 51850 18664
rect 51804 18360 51810 18652
rect 51844 18360 51850 18652
rect 51804 18348 51850 18360
rect 52862 18652 52908 18664
rect 52862 18360 52868 18652
rect 52902 18360 52908 18652
rect 52862 18348 52908 18360
rect 53442 18352 53776 22570
rect 59572 22696 59614 24250
rect 59864 22696 60012 24250
rect 62106 24474 62152 24486
rect 62106 24182 62112 24474
rect 62146 24182 62152 24474
rect 62106 24170 62152 24182
rect 63164 24474 63210 24486
rect 63164 24182 63170 24474
rect 63204 24182 63210 24474
rect 63164 24170 63210 24182
rect 64222 24474 64268 24486
rect 64222 24182 64228 24474
rect 64262 24182 64268 24474
rect 64222 24170 64268 24182
rect 65280 24474 65326 24486
rect 65280 24182 65286 24474
rect 65320 24182 65326 24474
rect 65280 24170 65326 24182
rect 66338 24474 66384 24486
rect 66338 24182 66344 24474
rect 66378 24182 66384 24474
rect 66338 24170 66384 24182
rect 67396 24474 67442 24486
rect 67396 24182 67402 24474
rect 67436 24182 67442 24474
rect 67396 24170 67442 24182
rect 68568 24472 68614 24484
rect 68568 24180 68574 24472
rect 68608 24180 68614 24472
rect 68568 24168 68614 24180
rect 69626 24472 69672 24484
rect 69626 24180 69632 24472
rect 69666 24180 69672 24472
rect 69626 24168 69672 24180
rect 70684 24472 70730 24484
rect 70684 24180 70690 24472
rect 70724 24180 70730 24472
rect 70684 24168 70730 24180
rect 71742 24472 71788 24484
rect 71742 24180 71748 24472
rect 71782 24180 71788 24472
rect 71742 24168 71788 24180
rect 72800 24472 72846 24484
rect 72800 24180 72806 24472
rect 72840 24180 72846 24472
rect 72800 24168 72846 24180
rect 73858 24472 73904 24484
rect 73858 24180 73864 24472
rect 73898 24180 73904 24472
rect 73858 24168 73904 24180
rect 75262 24446 75308 24458
rect 59572 22418 60012 22696
rect 61458 24034 61608 24160
rect 61458 22838 61480 24034
rect 61574 23280 61608 24034
rect 67920 24032 68070 24158
rect 75262 24154 75268 24446
rect 75302 24154 75308 24446
rect 75262 24142 75308 24154
rect 76320 24446 76366 24458
rect 76320 24154 76326 24446
rect 76360 24154 76366 24446
rect 76320 24142 76366 24154
rect 77378 24446 77424 24458
rect 77378 24154 77384 24446
rect 77418 24154 77424 24446
rect 77378 24142 77424 24154
rect 78436 24446 78482 24458
rect 78436 24154 78442 24446
rect 78476 24154 78482 24446
rect 78436 24142 78482 24154
rect 79494 24446 79540 24458
rect 79494 24154 79500 24446
rect 79534 24154 79540 24446
rect 79494 24142 79540 24154
rect 80552 24446 80598 24458
rect 80552 24154 80558 24446
rect 80592 24154 80598 24446
rect 80552 24142 80598 24154
rect 81724 24444 81770 24456
rect 81724 24152 81730 24444
rect 81764 24152 81770 24444
rect 81724 24140 81770 24152
rect 82782 24444 82828 24456
rect 82782 24152 82788 24444
rect 82822 24152 82828 24444
rect 82782 24140 82828 24152
rect 83840 24444 83886 24456
rect 83840 24152 83846 24444
rect 83880 24152 83886 24444
rect 83840 24140 83886 24152
rect 84898 24444 84944 24456
rect 84898 24152 84904 24444
rect 84938 24152 84944 24444
rect 84898 24140 84944 24152
rect 85956 24444 86002 24456
rect 85956 24152 85962 24444
rect 85996 24152 86002 24444
rect 85956 24140 86002 24152
rect 87014 24444 87060 24456
rect 87014 24152 87020 24444
rect 87054 24152 87060 24444
rect 87014 24140 87060 24152
rect 88496 24438 88542 24450
rect 88496 24146 88502 24438
rect 88536 24146 88542 24438
rect 88496 24134 88542 24146
rect 89554 24438 89600 24450
rect 89554 24146 89560 24438
rect 89594 24146 89600 24438
rect 89554 24134 89600 24146
rect 90612 24438 90658 24450
rect 90612 24146 90618 24438
rect 90652 24146 90658 24438
rect 90612 24134 90658 24146
rect 91670 24438 91716 24450
rect 91670 24146 91676 24438
rect 91710 24146 91716 24438
rect 91670 24134 91716 24146
rect 92728 24438 92774 24450
rect 92728 24146 92734 24438
rect 92768 24146 92774 24438
rect 92728 24134 92774 24146
rect 93786 24438 93832 24450
rect 93786 24146 93792 24438
rect 93826 24146 93832 24438
rect 93786 24134 93832 24146
rect 94958 24436 95004 24448
rect 94958 24144 94964 24436
rect 94998 24144 95004 24436
rect 94958 24132 95004 24144
rect 96016 24436 96062 24448
rect 96016 24144 96022 24436
rect 96056 24144 96062 24436
rect 96016 24132 96062 24144
rect 97074 24436 97120 24448
rect 97074 24144 97080 24436
rect 97114 24144 97120 24436
rect 97074 24132 97120 24144
rect 98132 24436 98178 24448
rect 98132 24144 98138 24436
rect 98172 24144 98178 24436
rect 98132 24132 98178 24144
rect 99190 24436 99236 24448
rect 99190 24144 99196 24436
rect 99230 24144 99236 24436
rect 100248 24436 100294 24448
rect 100248 24350 100254 24436
rect 100232 24224 100254 24350
rect 99190 24132 99236 24144
rect 100248 24144 100254 24224
rect 100288 24350 100294 24436
rect 100676 24350 100786 25032
rect 100288 24224 100786 24350
rect 100288 24144 100294 24224
rect 100248 24132 100294 24144
rect 67920 23790 67942 24032
rect 62106 23380 62152 23392
rect 62106 23280 62112 23380
rect 61574 23154 62112 23280
rect 61574 22838 61608 23154
rect 62106 23088 62112 23154
rect 62146 23088 62152 23380
rect 62106 23076 62152 23088
rect 63164 23380 63210 23392
rect 63164 23088 63170 23380
rect 63204 23088 63210 23380
rect 63164 23076 63210 23088
rect 64222 23380 64268 23392
rect 64222 23088 64228 23380
rect 64262 23088 64268 23380
rect 64222 23076 64268 23088
rect 65280 23380 65326 23392
rect 65280 23088 65286 23380
rect 65320 23088 65326 23380
rect 65280 23076 65326 23088
rect 66338 23380 66384 23392
rect 66338 23088 66344 23380
rect 66378 23088 66384 23380
rect 66338 23076 66384 23088
rect 67396 23380 67442 23392
rect 67396 23088 67402 23380
rect 67436 23088 67442 23380
rect 67396 23076 67442 23088
rect 61458 22514 61608 22838
rect 67596 22836 67942 23790
rect 68036 23790 68070 24032
rect 74614 24006 74764 24132
rect 68036 22836 68186 23790
rect 74614 23606 74636 24006
rect 68568 23378 68614 23390
rect 68568 23086 68574 23378
rect 68608 23086 68614 23378
rect 68568 23074 68614 23086
rect 69626 23378 69672 23390
rect 69626 23086 69632 23378
rect 69666 23086 69672 23378
rect 69626 23074 69672 23086
rect 70684 23378 70730 23390
rect 70684 23086 70690 23378
rect 70724 23086 70730 23378
rect 70684 23074 70730 23086
rect 71742 23378 71788 23390
rect 71742 23086 71748 23378
rect 71782 23086 71788 23378
rect 71742 23074 71788 23086
rect 72800 23378 72846 23390
rect 72800 23086 72806 23378
rect 72840 23086 72846 23378
rect 72800 23074 72846 23086
rect 73858 23378 73904 23390
rect 73858 23086 73864 23378
rect 73898 23086 73904 23378
rect 73858 23074 73904 23086
rect 54086 22342 54132 22354
rect 54086 22050 54092 22342
rect 54126 22050 54132 22342
rect 54086 22038 54132 22050
rect 55144 22342 55190 22354
rect 55144 22050 55150 22342
rect 55184 22050 55190 22342
rect 55144 22038 55190 22050
rect 56202 22342 56248 22354
rect 56202 22050 56208 22342
rect 56242 22050 56248 22342
rect 56202 22038 56248 22050
rect 57260 22342 57306 22354
rect 57260 22050 57266 22342
rect 57300 22050 57306 22342
rect 57260 22038 57306 22050
rect 58318 22342 58364 22354
rect 58318 22050 58324 22342
rect 58358 22050 58364 22342
rect 58318 22038 58364 22050
rect 59376 22342 59422 22354
rect 59376 22050 59382 22342
rect 59416 22050 59422 22342
rect 59376 22038 59422 22050
rect 54086 21248 54132 21260
rect 54086 20956 54092 21248
rect 54126 20956 54132 21248
rect 54086 20944 54132 20956
rect 55144 21248 55190 21260
rect 55144 20956 55150 21248
rect 55184 20956 55190 21248
rect 55144 20944 55190 20956
rect 56202 21248 56248 21260
rect 56202 20956 56208 21248
rect 56242 20956 56248 21248
rect 56202 20944 56248 20956
rect 57260 21248 57306 21260
rect 57260 20956 57266 21248
rect 57300 20956 57306 21248
rect 57260 20944 57306 20956
rect 58318 21248 58364 21260
rect 58318 20956 58324 21248
rect 58358 20956 58364 21248
rect 58318 20944 58364 20956
rect 59376 21248 59422 21260
rect 59376 20956 59382 21248
rect 59416 20956 59422 21248
rect 59376 20944 59422 20956
rect 54086 19760 54132 19772
rect 54086 19468 54092 19760
rect 54126 19468 54132 19760
rect 54086 19456 54132 19468
rect 55144 19760 55190 19772
rect 55144 19468 55150 19760
rect 55184 19468 55190 19760
rect 55144 19456 55190 19468
rect 56202 19760 56248 19772
rect 56202 19468 56208 19760
rect 56242 19468 56248 19760
rect 56202 19456 56248 19468
rect 57260 19760 57306 19772
rect 57260 19468 57266 19760
rect 57300 19468 57306 19760
rect 57260 19456 57306 19468
rect 58318 19760 58364 19772
rect 58318 19468 58324 19760
rect 58358 19468 58364 19760
rect 58318 19456 58364 19468
rect 59376 19760 59422 19772
rect 59376 19468 59382 19760
rect 59416 19468 59422 19760
rect 59376 19456 59422 19468
rect 59680 18686 60012 22418
rect 62106 22286 62152 22298
rect 62106 21994 62112 22286
rect 62146 21994 62152 22286
rect 62106 21982 62152 21994
rect 63164 22286 63210 22298
rect 63164 21994 63170 22286
rect 63204 21994 63210 22286
rect 63164 21982 63210 21994
rect 64222 22286 64268 22298
rect 64222 21994 64228 22286
rect 64262 21994 64268 22286
rect 64222 21982 64268 21994
rect 65280 22286 65326 22298
rect 65280 21994 65286 22286
rect 65320 21994 65326 22286
rect 65280 21982 65326 21994
rect 66338 22286 66384 22298
rect 66338 21994 66344 22286
rect 66378 21994 66384 22286
rect 66338 21982 66384 21994
rect 67396 22286 67442 22298
rect 67396 21994 67402 22286
rect 67436 21994 67442 22286
rect 67396 21982 67442 21994
rect 62106 21192 62152 21204
rect 62106 21012 62112 21192
rect 62080 20900 62112 21012
rect 62146 21012 62152 21192
rect 63164 21192 63210 21204
rect 62146 20900 62180 21012
rect 62080 19730 62180 20900
rect 63164 20900 63170 21192
rect 63204 20900 63210 21192
rect 63164 20888 63210 20900
rect 64222 21192 64268 21204
rect 64222 20900 64228 21192
rect 64262 20900 64268 21192
rect 64222 20888 64268 20900
rect 65280 21192 65326 21204
rect 65280 20900 65286 21192
rect 65320 20900 65326 21192
rect 65280 20888 65326 20900
rect 66338 21192 66384 21204
rect 66338 20900 66344 21192
rect 66378 20900 66384 21192
rect 67396 21192 67442 21204
rect 67396 21044 67402 21192
rect 66338 20888 66384 20900
rect 67374 20900 67402 21044
rect 67436 21044 67442 21192
rect 67436 20900 67474 21044
rect 62080 19560 62118 19730
rect 62112 19438 62118 19560
rect 62152 19560 62180 19730
rect 63170 19730 63216 19742
rect 62152 19438 62158 19560
rect 62112 19426 62158 19438
rect 63170 19438 63176 19730
rect 63210 19438 63216 19730
rect 63170 19426 63216 19438
rect 64228 19730 64274 19742
rect 64228 19438 64234 19730
rect 64268 19438 64274 19730
rect 64228 19426 64274 19438
rect 65286 19730 65332 19742
rect 65286 19438 65292 19730
rect 65326 19438 65332 19730
rect 65286 19426 65332 19438
rect 66344 19730 66390 19742
rect 66344 19438 66350 19730
rect 66384 19438 66390 19730
rect 67374 19730 67474 20900
rect 67374 19592 67408 19730
rect 66344 19426 66390 19438
rect 67402 19438 67408 19592
rect 67442 19592 67474 19730
rect 67442 19438 67448 19592
rect 67402 19426 67448 19438
rect 54086 18666 54132 18678
rect 54086 18374 54092 18666
rect 54126 18374 54132 18666
rect 54086 18362 54132 18374
rect 55144 18666 55190 18678
rect 55144 18374 55150 18666
rect 55184 18374 55190 18666
rect 55144 18362 55190 18374
rect 56202 18666 56248 18678
rect 56202 18374 56208 18666
rect 56242 18374 56248 18666
rect 56202 18362 56248 18374
rect 57260 18666 57306 18678
rect 57260 18374 57266 18666
rect 57300 18374 57306 18666
rect 57260 18362 57306 18374
rect 58318 18666 58364 18678
rect 58318 18374 58324 18666
rect 58358 18374 58364 18666
rect 58318 18362 58364 18374
rect 59376 18666 59422 18678
rect 59376 18374 59382 18666
rect 59416 18374 59422 18666
rect 59376 18362 59422 18374
rect 59628 18464 60012 18686
rect 40984 17536 41030 17548
rect 40984 17244 40990 17536
rect 41024 17244 41030 17536
rect 40984 17232 41030 17244
rect 42042 17536 42088 17548
rect 42042 17244 42048 17536
rect 42082 17244 42088 17536
rect 42042 17232 42088 17244
rect 43100 17536 43146 17548
rect 43100 17244 43106 17536
rect 43140 17244 43146 17536
rect 43100 17232 43146 17244
rect 44158 17536 44204 17548
rect 44158 17244 44164 17536
rect 44198 17244 44204 17536
rect 44158 17232 44204 17244
rect 45216 17536 45262 17548
rect 45216 17244 45222 17536
rect 45256 17244 45262 17536
rect 45216 17232 45262 17244
rect 46274 17536 46320 17548
rect 46274 17244 46280 17536
rect 46314 17244 46320 17536
rect 46274 17232 46320 17244
rect 34494 16442 34540 16454
rect 34494 16150 34500 16442
rect 34534 16150 34540 16442
rect 34494 16138 34540 16150
rect 35552 16442 35598 16454
rect 35552 16150 35558 16442
rect 35592 16150 35598 16442
rect 35552 16138 35598 16150
rect 36610 16442 36656 16454
rect 36610 16150 36616 16442
rect 36650 16150 36656 16442
rect 36610 16138 36656 16150
rect 37668 16442 37714 16454
rect 37668 16150 37674 16442
rect 37708 16150 37714 16442
rect 37668 16138 37714 16150
rect 38726 16442 38772 16454
rect 38726 16150 38732 16442
rect 38766 16150 38772 16442
rect 38726 16138 38772 16150
rect 39784 16442 39830 16454
rect 39784 16150 39790 16442
rect 39824 16150 39830 16442
rect 39784 16138 39830 16150
rect 34494 15348 34540 15360
rect 34494 15056 34500 15348
rect 34534 15056 34540 15348
rect 34494 15044 34540 15056
rect 35552 15348 35598 15360
rect 35552 15056 35558 15348
rect 35592 15056 35598 15348
rect 35552 15044 35598 15056
rect 36610 15348 36656 15360
rect 36610 15056 36616 15348
rect 36650 15056 36656 15348
rect 36610 15044 36656 15056
rect 37668 15348 37714 15360
rect 37668 15056 37674 15348
rect 37708 15056 37714 15348
rect 37668 15044 37714 15056
rect 38726 15348 38772 15360
rect 38726 15056 38732 15348
rect 38766 15056 38772 15348
rect 38726 15044 38772 15056
rect 39784 15348 39830 15360
rect 39784 15056 39790 15348
rect 39824 15056 39830 15348
rect 39784 15044 39830 15056
rect 34504 13868 34550 13880
rect 34504 13576 34510 13868
rect 34544 13576 34550 13868
rect 34504 13564 34550 13576
rect 35562 13868 35608 13880
rect 35562 13576 35568 13868
rect 35602 13576 35608 13868
rect 35562 13564 35608 13576
rect 36620 13868 36666 13880
rect 36620 13576 36626 13868
rect 36660 13576 36666 13868
rect 36620 13564 36666 13576
rect 37678 13868 37724 13880
rect 37678 13576 37684 13868
rect 37718 13576 37724 13868
rect 37678 13564 37724 13576
rect 38736 13868 38782 13880
rect 38736 13576 38742 13868
rect 38776 13576 38782 13868
rect 38736 13564 38782 13576
rect 39794 13868 39840 13880
rect 39794 13576 39800 13868
rect 39834 13576 39840 13868
rect 39794 13564 39840 13576
rect 34504 12774 34550 12786
rect 34504 12482 34510 12774
rect 34544 12482 34550 12774
rect 34504 12470 34550 12482
rect 35562 12774 35608 12786
rect 35562 12482 35568 12774
rect 35602 12482 35608 12774
rect 35562 12470 35608 12482
rect 36620 12774 36666 12786
rect 36620 12482 36626 12774
rect 36660 12482 36666 12774
rect 36620 12470 36666 12482
rect 37678 12774 37724 12786
rect 37678 12482 37684 12774
rect 37718 12482 37724 12774
rect 37678 12470 37724 12482
rect 38736 12774 38782 12786
rect 38736 12482 38742 12774
rect 38776 12482 38782 12774
rect 38736 12470 38782 12482
rect 39794 12774 39840 12786
rect 39794 12482 39800 12774
rect 39834 12482 39840 12774
rect 39794 12470 39840 12482
rect 27994 11674 28040 11686
rect 27994 11382 28000 11674
rect 28034 11382 28040 11674
rect 27994 11370 28040 11382
rect 29052 11674 29098 11686
rect 29052 11382 29058 11674
rect 29092 11382 29098 11674
rect 29052 11370 29098 11382
rect 30110 11674 30156 11686
rect 30110 11382 30116 11674
rect 30150 11382 30156 11674
rect 30110 11370 30156 11382
rect 31168 11674 31214 11686
rect 31168 11382 31174 11674
rect 31208 11382 31214 11674
rect 31168 11370 31214 11382
rect 32226 11674 32272 11686
rect 32226 11382 32232 11674
rect 32266 11382 32272 11674
rect 32226 11370 32272 11382
rect 33284 11674 33330 11686
rect 33284 11382 33290 11674
rect 33324 11382 33330 11674
rect 33284 11370 33330 11382
rect 21472 10564 21518 10576
rect 21472 10272 21478 10564
rect 21512 10272 21518 10564
rect 21472 10260 21518 10272
rect 22530 10564 22576 10576
rect 22530 10272 22536 10564
rect 22570 10272 22576 10564
rect 22530 10260 22576 10272
rect 23588 10564 23634 10576
rect 23588 10272 23594 10564
rect 23628 10272 23634 10564
rect 23588 10260 23634 10272
rect 24646 10564 24692 10576
rect 24646 10272 24652 10564
rect 24686 10272 24692 10564
rect 24646 10260 24692 10272
rect 25704 10564 25750 10576
rect 25704 10272 25710 10564
rect 25744 10272 25750 10564
rect 25704 10260 25750 10272
rect 26762 10564 26808 10576
rect 26762 10272 26768 10564
rect 26802 10272 26808 10564
rect 26762 10260 26808 10272
rect 21472 9470 21518 9482
rect 21472 9178 21478 9470
rect 21512 9178 21518 9470
rect 21472 9166 21518 9178
rect 22530 9470 22576 9482
rect 22530 9178 22536 9470
rect 22570 9178 22576 9470
rect 22530 9166 22576 9178
rect 23588 9470 23634 9482
rect 23588 9178 23594 9470
rect 23628 9178 23634 9470
rect 23588 9166 23634 9178
rect 24646 9470 24692 9482
rect 24646 9178 24652 9470
rect 24686 9178 24692 9470
rect 24646 9166 24692 9178
rect 25704 9470 25750 9482
rect 25704 9178 25710 9470
rect 25744 9178 25750 9470
rect 25704 9166 25750 9178
rect 26762 9470 26808 9482
rect 26762 9178 26768 9470
rect 26802 9178 26808 9470
rect 26762 9166 26808 9178
rect 21490 7938 21536 7950
rect 21490 7646 21496 7938
rect 21530 7646 21536 7938
rect 21490 7634 21536 7646
rect 22548 7938 22594 7950
rect 22548 7646 22554 7938
rect 22588 7646 22594 7938
rect 22548 7634 22594 7646
rect 23606 7938 23652 7950
rect 23606 7646 23612 7938
rect 23646 7646 23652 7938
rect 23606 7634 23652 7646
rect 24664 7938 24710 7950
rect 24664 7646 24670 7938
rect 24704 7646 24710 7938
rect 24664 7634 24710 7646
rect 25722 7938 25768 7950
rect 25722 7646 25728 7938
rect 25762 7646 25768 7938
rect 25722 7634 25768 7646
rect 26780 7938 26826 7950
rect 26780 7646 26786 7938
rect 26820 7646 26826 7938
rect 26780 7634 26826 7646
rect 21490 6844 21536 6856
rect 21490 6552 21496 6844
rect 21530 6552 21536 6844
rect 21490 6540 21536 6552
rect 22548 6844 22594 6856
rect 22548 6552 22554 6844
rect 22588 6552 22594 6844
rect 22548 6540 22594 6552
rect 23606 6844 23652 6856
rect 23606 6552 23612 6844
rect 23646 6552 23652 6844
rect 23606 6540 23652 6552
rect 24664 6844 24710 6856
rect 24664 6552 24670 6844
rect 24704 6552 24710 6844
rect 24664 6540 24710 6552
rect 25722 6844 25768 6856
rect 25722 6552 25728 6844
rect 25762 6552 25768 6844
rect 25722 6540 25768 6552
rect 26780 6844 26826 6856
rect 26780 6552 26786 6844
rect 26820 6552 26826 6844
rect 26780 6540 26826 6552
rect 15000 5766 15046 5778
rect 15000 5474 15006 5766
rect 15040 5474 15046 5766
rect 15000 5462 15046 5474
rect 16058 5766 16104 5778
rect 16058 5474 16064 5766
rect 16098 5474 16104 5766
rect 16058 5462 16104 5474
rect 17116 5766 17162 5778
rect 17116 5474 17122 5766
rect 17156 5474 17162 5766
rect 17116 5462 17162 5474
rect 18174 5766 18220 5778
rect 18174 5474 18180 5766
rect 18214 5474 18220 5766
rect 18174 5462 18220 5474
rect 19232 5766 19278 5778
rect 19232 5474 19238 5766
rect 19272 5474 19278 5766
rect 19232 5462 19278 5474
rect 20290 5766 20336 5778
rect 20290 5474 20296 5766
rect 20330 5474 20336 5766
rect 20290 5462 20336 5474
rect 8494 4664 8540 4676
rect 8494 4372 8500 4664
rect 8534 4372 8540 4664
rect 8494 4360 8540 4372
rect 9552 4664 9598 4676
rect 9552 4372 9558 4664
rect 9592 4372 9598 4664
rect 9552 4360 9598 4372
rect 10610 4664 10656 4676
rect 10610 4372 10616 4664
rect 10650 4372 10656 4664
rect 10610 4360 10656 4372
rect 11668 4664 11714 4676
rect 11668 4372 11674 4664
rect 11708 4372 11714 4664
rect 11668 4360 11714 4372
rect 12726 4664 12772 4676
rect 12726 4372 12732 4664
rect 12766 4372 12772 4664
rect 12726 4360 12772 4372
rect 13784 4664 13830 4676
rect 13784 4372 13790 4664
rect 13824 4372 13830 4664
rect 13784 4360 13830 4372
rect 8494 3570 8540 3582
rect 8494 3278 8500 3570
rect 8534 3278 8540 3570
rect 8494 3266 8540 3278
rect 9552 3570 9598 3582
rect 9552 3278 9558 3570
rect 9592 3278 9598 3570
rect 9552 3266 9598 3278
rect 10610 3570 10656 3582
rect 10610 3278 10616 3570
rect 10650 3278 10656 3570
rect 10610 3266 10656 3278
rect 11668 3570 11714 3582
rect 11668 3278 11674 3570
rect 11708 3278 11714 3570
rect 11668 3266 11714 3278
rect 12726 3570 12772 3582
rect 12726 3278 12732 3570
rect 12766 3278 12772 3570
rect 12726 3266 12772 3278
rect 13784 3570 13830 3582
rect 13784 3278 13790 3570
rect 13824 3278 13830 3570
rect 13784 3266 13830 3278
rect 14216 -3192 14512 5224
rect 20748 5208 20864 6404
rect 20958 5208 21044 6404
rect 27278 6420 27574 11132
rect 33848 11138 33878 12334
rect 33972 11138 34144 12334
rect 40304 12334 40638 16994
rect 46836 17016 46946 18212
rect 47040 17016 47170 18212
rect 53438 18226 53776 18352
rect 47572 17558 47618 17570
rect 47572 17266 47578 17558
rect 47612 17266 47618 17558
rect 47572 17254 47618 17266
rect 48630 17558 48676 17570
rect 48630 17266 48636 17558
rect 48670 17266 48676 17558
rect 48630 17254 48676 17266
rect 49688 17558 49734 17570
rect 49688 17266 49694 17558
rect 49728 17266 49734 17558
rect 49688 17254 49734 17266
rect 50746 17558 50792 17570
rect 50746 17266 50752 17558
rect 50786 17266 50792 17558
rect 50746 17254 50792 17266
rect 51804 17558 51850 17570
rect 51804 17266 51810 17558
rect 51844 17266 51850 17558
rect 51804 17254 51850 17266
rect 52862 17558 52908 17570
rect 52862 17266 52868 17558
rect 52902 17266 52908 17558
rect 52862 17254 52908 17266
rect 40984 16442 41030 16454
rect 40984 16150 40990 16442
rect 41024 16150 41030 16442
rect 40984 16138 41030 16150
rect 42042 16442 42088 16454
rect 42042 16150 42048 16442
rect 42082 16150 42088 16442
rect 42042 16138 42088 16150
rect 43100 16442 43146 16454
rect 43100 16150 43106 16442
rect 43140 16150 43146 16442
rect 43100 16138 43146 16150
rect 44158 16442 44204 16454
rect 44158 16150 44164 16442
rect 44198 16150 44204 16442
rect 44158 16138 44204 16150
rect 45216 16442 45262 16454
rect 45216 16150 45222 16442
rect 45256 16150 45262 16442
rect 45216 16138 45262 16150
rect 46274 16442 46320 16454
rect 46274 16150 46280 16442
rect 46314 16150 46320 16442
rect 46274 16138 46320 16150
rect 40984 15348 41030 15360
rect 40984 15056 40990 15348
rect 41024 15056 41030 15348
rect 40984 15044 41030 15056
rect 42042 15348 42088 15360
rect 42042 15056 42048 15348
rect 42082 15056 42088 15348
rect 42042 15044 42088 15056
rect 43100 15348 43146 15360
rect 43100 15056 43106 15348
rect 43140 15056 43146 15348
rect 43100 15044 43146 15056
rect 44158 15348 44204 15360
rect 44158 15056 44164 15348
rect 44198 15056 44204 15348
rect 44158 15044 44204 15056
rect 45216 15348 45262 15360
rect 45216 15056 45222 15348
rect 45256 15056 45262 15348
rect 45216 15044 45262 15056
rect 46274 15348 46320 15360
rect 46274 15056 46280 15348
rect 46314 15056 46320 15348
rect 46274 15044 46320 15056
rect 40994 13868 41040 13880
rect 40994 13576 41000 13868
rect 41034 13576 41040 13868
rect 40994 13564 41040 13576
rect 42052 13868 42098 13880
rect 42052 13576 42058 13868
rect 42092 13576 42098 13868
rect 42052 13564 42098 13576
rect 43110 13868 43156 13880
rect 43110 13576 43116 13868
rect 43150 13576 43156 13868
rect 43110 13564 43156 13576
rect 44168 13868 44214 13880
rect 44168 13576 44174 13868
rect 44208 13576 44214 13868
rect 44168 13564 44214 13576
rect 45226 13868 45272 13880
rect 45226 13576 45232 13868
rect 45266 13576 45272 13868
rect 45226 13564 45272 13576
rect 46284 13868 46330 13880
rect 46284 13576 46290 13868
rect 46324 13576 46330 13868
rect 46284 13564 46330 13576
rect 40994 12774 41040 12786
rect 40994 12482 41000 12774
rect 41034 12482 41040 12774
rect 40994 12470 41040 12482
rect 42052 12774 42098 12786
rect 42052 12482 42058 12774
rect 42092 12482 42098 12774
rect 42052 12470 42098 12482
rect 43110 12774 43156 12786
rect 43110 12482 43116 12774
rect 43150 12482 43156 12774
rect 43110 12470 43156 12482
rect 44168 12774 44214 12786
rect 44168 12482 44174 12774
rect 44208 12482 44214 12774
rect 44168 12470 44214 12482
rect 45226 12774 45272 12786
rect 45226 12482 45232 12774
rect 45266 12482 45272 12774
rect 45226 12470 45272 12482
rect 46284 12774 46330 12786
rect 46284 12482 46290 12774
rect 46324 12482 46330 12774
rect 46284 12470 46330 12482
rect 34504 11680 34550 11692
rect 34504 11388 34510 11680
rect 34544 11388 34550 11680
rect 34504 11376 34550 11388
rect 35562 11680 35608 11692
rect 35562 11388 35568 11680
rect 35602 11388 35608 11680
rect 35562 11376 35608 11388
rect 36620 11680 36666 11692
rect 36620 11388 36626 11680
rect 36660 11388 36666 11680
rect 36620 11376 36666 11388
rect 37678 11680 37724 11692
rect 37678 11388 37684 11680
rect 37718 11388 37724 11680
rect 37678 11376 37724 11388
rect 38736 11680 38782 11692
rect 38736 11388 38742 11680
rect 38776 11388 38782 11680
rect 38736 11376 38782 11388
rect 39794 11680 39840 11692
rect 39794 11388 39800 11680
rect 39834 11388 39840 11680
rect 39794 11376 39840 11388
rect 27994 10580 28040 10592
rect 27994 10288 28000 10580
rect 28034 10288 28040 10580
rect 27994 10276 28040 10288
rect 29052 10580 29098 10592
rect 29052 10288 29058 10580
rect 29092 10288 29098 10580
rect 29052 10276 29098 10288
rect 30110 10580 30156 10592
rect 30110 10288 30116 10580
rect 30150 10288 30156 10580
rect 30110 10276 30156 10288
rect 31168 10580 31214 10592
rect 31168 10288 31174 10580
rect 31208 10288 31214 10580
rect 31168 10276 31214 10288
rect 32226 10580 32272 10592
rect 32226 10288 32232 10580
rect 32266 10288 32272 10580
rect 32226 10276 32272 10288
rect 33284 10580 33330 10592
rect 33284 10288 33290 10580
rect 33324 10288 33330 10580
rect 33284 10276 33330 10288
rect 27994 9486 28040 9498
rect 27994 9194 28000 9486
rect 28034 9194 28040 9486
rect 27994 9182 28040 9194
rect 29052 9486 29098 9498
rect 29052 9194 29058 9486
rect 29092 9194 29098 9486
rect 29052 9182 29098 9194
rect 30110 9486 30156 9498
rect 30110 9194 30116 9486
rect 30150 9194 30156 9486
rect 30110 9182 30156 9194
rect 31168 9486 31214 9498
rect 31168 9194 31174 9486
rect 31208 9194 31214 9486
rect 31168 9182 31214 9194
rect 32226 9486 32272 9498
rect 32226 9194 32232 9486
rect 32266 9194 32272 9486
rect 32226 9182 32272 9194
rect 33284 9486 33330 9498
rect 33284 9194 33290 9486
rect 33324 9194 33330 9486
rect 33284 9182 33330 9194
rect 28012 7954 28058 7966
rect 28012 7662 28018 7954
rect 28052 7662 28058 7954
rect 28012 7650 28058 7662
rect 29070 7954 29116 7966
rect 29070 7662 29076 7954
rect 29110 7662 29116 7954
rect 29070 7650 29116 7662
rect 30128 7954 30174 7966
rect 30128 7662 30134 7954
rect 30168 7662 30174 7954
rect 30128 7650 30174 7662
rect 31186 7954 31232 7966
rect 31186 7662 31192 7954
rect 31226 7662 31232 7954
rect 31186 7650 31232 7662
rect 32244 7954 32290 7966
rect 32244 7662 32250 7954
rect 32284 7662 32290 7954
rect 32244 7650 32290 7662
rect 33302 7954 33348 7966
rect 33302 7662 33308 7954
rect 33342 7662 33348 7954
rect 33302 7650 33348 7662
rect 28012 6860 28058 6872
rect 28012 6568 28018 6860
rect 28052 6568 28058 6860
rect 28012 6556 28058 6568
rect 29070 6860 29116 6872
rect 29070 6568 29076 6860
rect 29110 6568 29116 6860
rect 29070 6556 29116 6568
rect 30128 6860 30174 6872
rect 30128 6568 30134 6860
rect 30168 6568 30174 6860
rect 30128 6556 30174 6568
rect 31186 6860 31232 6872
rect 31186 6568 31192 6860
rect 31226 6568 31232 6860
rect 31186 6556 31232 6568
rect 32244 6860 32290 6872
rect 32244 6568 32250 6860
rect 32284 6568 32290 6860
rect 32244 6556 32290 6568
rect 33302 6860 33348 6872
rect 33302 6568 33308 6860
rect 33342 6568 33348 6860
rect 33302 6556 33348 6568
rect 21490 5750 21536 5762
rect 21490 5458 21496 5750
rect 21530 5458 21536 5750
rect 21490 5446 21536 5458
rect 22548 5750 22594 5762
rect 22548 5458 22554 5750
rect 22588 5458 22594 5750
rect 22548 5446 22594 5458
rect 23606 5750 23652 5762
rect 23606 5458 23612 5750
rect 23646 5458 23652 5750
rect 23606 5446 23652 5458
rect 24664 5750 24710 5762
rect 24664 5458 24670 5750
rect 24704 5458 24710 5750
rect 24664 5446 24710 5458
rect 25722 5750 25768 5762
rect 25722 5458 25728 5750
rect 25762 5458 25768 5750
rect 25722 5446 25768 5458
rect 26780 5750 26826 5762
rect 26780 5458 26786 5750
rect 26820 5458 26826 5750
rect 26780 5446 26826 5458
rect 15000 4672 15046 4684
rect 15000 4380 15006 4672
rect 15040 4380 15046 4672
rect 15000 4368 15046 4380
rect 16058 4672 16104 4684
rect 16058 4380 16064 4672
rect 16098 4380 16104 4672
rect 16058 4368 16104 4380
rect 17116 4672 17162 4684
rect 17116 4380 17122 4672
rect 17156 4380 17162 4672
rect 17116 4368 17162 4380
rect 18174 4672 18220 4684
rect 18174 4380 18180 4672
rect 18214 4380 18220 4672
rect 18174 4368 18220 4380
rect 19232 4672 19278 4684
rect 19232 4380 19238 4672
rect 19272 4380 19278 4672
rect 19232 4368 19278 4380
rect 20290 4672 20336 4684
rect 20290 4380 20296 4672
rect 20330 4380 20336 4672
rect 20290 4368 20336 4380
rect 15000 3578 15046 3590
rect 15000 3286 15006 3578
rect 15040 3286 15046 3578
rect 15000 3274 15046 3286
rect 16058 3578 16104 3590
rect 16058 3286 16064 3578
rect 16098 3286 16104 3578
rect 16058 3274 16104 3286
rect 17116 3578 17162 3590
rect 17116 3286 17122 3578
rect 17156 3286 17162 3578
rect 17116 3274 17162 3286
rect 18174 3578 18220 3590
rect 18174 3286 18180 3578
rect 18214 3286 18220 3578
rect 18174 3274 18220 3286
rect 19232 3578 19278 3590
rect 19232 3286 19238 3578
rect 19272 3286 19278 3578
rect 19232 3274 19278 3286
rect 20290 3578 20336 3590
rect 20290 3286 20296 3578
rect 20330 3286 20336 3578
rect 20290 3274 20336 3286
rect 20748 -3192 21044 5208
rect 27278 5224 27386 6420
rect 27480 5224 27574 6420
rect 33848 6426 34144 11138
rect 40304 11138 40368 12334
rect 40462 11138 40638 12334
rect 46836 12356 47170 17016
rect 53438 17030 53460 18226
rect 53554 17030 53776 18226
rect 54086 17572 54132 17584
rect 54086 17280 54092 17572
rect 54126 17280 54132 17572
rect 54086 17268 54132 17280
rect 55144 17572 55190 17584
rect 55144 17280 55150 17572
rect 55184 17280 55190 17572
rect 55144 17268 55190 17280
rect 56202 17572 56248 17584
rect 56202 17280 56208 17572
rect 56242 17280 56248 17572
rect 56202 17268 56248 17280
rect 57260 17572 57306 17584
rect 57260 17280 57266 17572
rect 57300 17280 57306 17572
rect 57260 17268 57306 17280
rect 58318 17572 58364 17584
rect 58318 17280 58324 17572
rect 58358 17280 58364 17572
rect 58318 17268 58364 17280
rect 59376 17572 59422 17584
rect 59376 17280 59382 17572
rect 59416 17280 59422 17572
rect 59376 17268 59422 17280
rect 53438 16706 53776 17030
rect 47572 16464 47618 16476
rect 47572 16172 47578 16464
rect 47612 16172 47618 16464
rect 47572 16160 47618 16172
rect 48630 16464 48676 16476
rect 48630 16172 48636 16464
rect 48670 16172 48676 16464
rect 48630 16160 48676 16172
rect 49688 16464 49734 16476
rect 49688 16172 49694 16464
rect 49728 16172 49734 16464
rect 49688 16160 49734 16172
rect 50746 16464 50792 16476
rect 50746 16172 50752 16464
rect 50786 16172 50792 16464
rect 50746 16160 50792 16172
rect 51804 16464 51850 16476
rect 51804 16172 51810 16464
rect 51844 16172 51850 16464
rect 51804 16160 51850 16172
rect 52862 16464 52908 16476
rect 52862 16172 52868 16464
rect 52902 16172 52908 16464
rect 52862 16160 52908 16172
rect 47572 15370 47618 15382
rect 47572 15078 47578 15370
rect 47612 15078 47618 15370
rect 47572 15066 47618 15078
rect 48630 15370 48676 15382
rect 48630 15078 48636 15370
rect 48670 15078 48676 15370
rect 48630 15066 48676 15078
rect 49688 15370 49734 15382
rect 49688 15078 49694 15370
rect 49728 15078 49734 15370
rect 49688 15066 49734 15078
rect 50746 15370 50792 15382
rect 50746 15078 50752 15370
rect 50786 15078 50792 15370
rect 50746 15066 50792 15078
rect 51804 15370 51850 15382
rect 51804 15078 51810 15370
rect 51844 15078 51850 15370
rect 51804 15066 51850 15078
rect 52862 15370 52908 15382
rect 52862 15078 52868 15370
rect 52902 15078 52908 15370
rect 52862 15066 52908 15078
rect 47582 13890 47628 13902
rect 47582 13598 47588 13890
rect 47622 13598 47628 13890
rect 47582 13586 47628 13598
rect 48640 13890 48686 13902
rect 48640 13598 48646 13890
rect 48680 13598 48686 13890
rect 48640 13586 48686 13598
rect 49698 13890 49744 13902
rect 49698 13598 49704 13890
rect 49738 13598 49744 13890
rect 49698 13586 49744 13598
rect 50756 13890 50802 13902
rect 50756 13598 50762 13890
rect 50796 13598 50802 13890
rect 50756 13586 50802 13598
rect 51814 13890 51860 13902
rect 51814 13598 51820 13890
rect 51854 13598 51860 13890
rect 51814 13586 51860 13598
rect 52872 13890 52918 13902
rect 52872 13598 52878 13890
rect 52912 13598 52918 13890
rect 52872 13586 52918 13598
rect 47582 12796 47628 12808
rect 47582 12504 47588 12796
rect 47622 12504 47628 12796
rect 47582 12492 47628 12504
rect 48640 12796 48686 12808
rect 48640 12504 48646 12796
rect 48680 12504 48686 12796
rect 48640 12492 48686 12504
rect 49698 12796 49744 12808
rect 49698 12504 49704 12796
rect 49738 12504 49744 12796
rect 49698 12492 49744 12504
rect 50756 12796 50802 12808
rect 50756 12504 50762 12796
rect 50796 12504 50802 12796
rect 50756 12492 50802 12504
rect 51814 12796 51860 12808
rect 51814 12504 51820 12796
rect 51854 12504 51860 12796
rect 51814 12492 51860 12504
rect 52872 12796 52918 12808
rect 52872 12504 52878 12796
rect 52912 12504 52918 12796
rect 52872 12492 52918 12504
rect 40994 11680 41040 11692
rect 40994 11388 41000 11680
rect 41034 11388 41040 11680
rect 40994 11376 41040 11388
rect 42052 11680 42098 11692
rect 42052 11388 42058 11680
rect 42092 11388 42098 11680
rect 42052 11376 42098 11388
rect 43110 11680 43156 11692
rect 43110 11388 43116 11680
rect 43150 11388 43156 11680
rect 43110 11376 43156 11388
rect 44168 11680 44214 11692
rect 44168 11388 44174 11680
rect 44208 11388 44214 11680
rect 44168 11376 44214 11388
rect 45226 11680 45272 11692
rect 45226 11388 45232 11680
rect 45266 11388 45272 11680
rect 45226 11376 45272 11388
rect 46284 11680 46330 11692
rect 46284 11388 46290 11680
rect 46324 11388 46330 11680
rect 46284 11376 46330 11388
rect 34504 10586 34550 10598
rect 34504 10294 34510 10586
rect 34544 10294 34550 10586
rect 34504 10282 34550 10294
rect 35562 10586 35608 10598
rect 35562 10294 35568 10586
rect 35602 10294 35608 10586
rect 35562 10282 35608 10294
rect 36620 10586 36666 10598
rect 36620 10294 36626 10586
rect 36660 10294 36666 10586
rect 36620 10282 36666 10294
rect 37678 10586 37724 10598
rect 37678 10294 37684 10586
rect 37718 10294 37724 10586
rect 37678 10282 37724 10294
rect 38736 10586 38782 10598
rect 38736 10294 38742 10586
rect 38776 10294 38782 10586
rect 38736 10282 38782 10294
rect 39794 10586 39840 10598
rect 39794 10294 39800 10586
rect 39834 10294 39840 10586
rect 39794 10282 39840 10294
rect 34504 9492 34550 9504
rect 34504 9200 34510 9492
rect 34544 9200 34550 9492
rect 34504 9188 34550 9200
rect 35562 9492 35608 9504
rect 35562 9200 35568 9492
rect 35602 9200 35608 9492
rect 35562 9188 35608 9200
rect 36620 9492 36666 9504
rect 36620 9200 36626 9492
rect 36660 9200 36666 9492
rect 36620 9188 36666 9200
rect 37678 9492 37724 9504
rect 37678 9200 37684 9492
rect 37718 9200 37724 9492
rect 37678 9188 37724 9200
rect 38736 9492 38782 9504
rect 38736 9200 38742 9492
rect 38776 9200 38782 9492
rect 38736 9188 38782 9200
rect 39794 9492 39840 9504
rect 39794 9200 39800 9492
rect 39834 9200 39840 9492
rect 39794 9188 39840 9200
rect 34522 7960 34568 7972
rect 34522 7668 34528 7960
rect 34562 7668 34568 7960
rect 34522 7656 34568 7668
rect 35580 7960 35626 7972
rect 35580 7668 35586 7960
rect 35620 7668 35626 7960
rect 35580 7656 35626 7668
rect 36638 7960 36684 7972
rect 36638 7668 36644 7960
rect 36678 7668 36684 7960
rect 36638 7656 36684 7668
rect 37696 7960 37742 7972
rect 37696 7668 37702 7960
rect 37736 7668 37742 7960
rect 37696 7656 37742 7668
rect 38754 7960 38800 7972
rect 38754 7668 38760 7960
rect 38794 7668 38800 7960
rect 38754 7656 38800 7668
rect 39812 7960 39858 7972
rect 39812 7668 39818 7960
rect 39852 7668 39858 7960
rect 39812 7656 39858 7668
rect 34522 6866 34568 6878
rect 34522 6574 34528 6866
rect 34562 6574 34568 6866
rect 34522 6562 34568 6574
rect 35580 6866 35626 6878
rect 35580 6574 35586 6866
rect 35620 6574 35626 6866
rect 35580 6562 35626 6574
rect 36638 6866 36684 6878
rect 36638 6574 36644 6866
rect 36678 6574 36684 6866
rect 36638 6562 36684 6574
rect 37696 6866 37742 6878
rect 37696 6574 37702 6866
rect 37736 6574 37742 6866
rect 37696 6562 37742 6574
rect 38754 6866 38800 6878
rect 38754 6574 38760 6866
rect 38794 6574 38800 6866
rect 38754 6562 38800 6574
rect 39812 6866 39858 6878
rect 39812 6574 39818 6866
rect 39852 6574 39858 6866
rect 39812 6562 39858 6574
rect 28012 5766 28058 5778
rect 28012 5474 28018 5766
rect 28052 5474 28058 5766
rect 28012 5462 28058 5474
rect 29070 5766 29116 5778
rect 29070 5474 29076 5766
rect 29110 5474 29116 5766
rect 29070 5462 29116 5474
rect 30128 5766 30174 5778
rect 30128 5474 30134 5766
rect 30168 5474 30174 5766
rect 30128 5462 30174 5474
rect 31186 5766 31232 5778
rect 31186 5474 31192 5766
rect 31226 5474 31232 5766
rect 31186 5462 31232 5474
rect 32244 5766 32290 5778
rect 32244 5474 32250 5766
rect 32284 5474 32290 5766
rect 32244 5462 32290 5474
rect 33302 5766 33348 5778
rect 33302 5474 33308 5766
rect 33342 5474 33348 5766
rect 33302 5462 33348 5474
rect 21490 4656 21536 4668
rect 21490 4364 21496 4656
rect 21530 4364 21536 4656
rect 21490 4352 21536 4364
rect 22548 4656 22594 4668
rect 22548 4364 22554 4656
rect 22588 4364 22594 4656
rect 22548 4352 22594 4364
rect 23606 4656 23652 4668
rect 23606 4364 23612 4656
rect 23646 4364 23652 4656
rect 23606 4352 23652 4364
rect 24664 4656 24710 4668
rect 24664 4364 24670 4656
rect 24704 4364 24710 4656
rect 24664 4352 24710 4364
rect 25722 4656 25768 4668
rect 25722 4364 25728 4656
rect 25762 4364 25768 4656
rect 25722 4352 25768 4364
rect 26780 4656 26826 4668
rect 26780 4364 26786 4656
rect 26820 4364 26826 4656
rect 26780 4352 26826 4364
rect 21490 3562 21536 3574
rect 21490 3270 21496 3562
rect 21530 3270 21536 3562
rect 21490 3258 21536 3270
rect 22548 3562 22594 3574
rect 22548 3270 22554 3562
rect 22588 3270 22594 3562
rect 22548 3258 22594 3270
rect 23606 3562 23652 3574
rect 23606 3270 23612 3562
rect 23646 3270 23652 3562
rect 23606 3258 23652 3270
rect 24664 3562 24710 3574
rect 24664 3270 24670 3562
rect 24704 3270 24710 3562
rect 24664 3258 24710 3270
rect 25722 3562 25768 3574
rect 25722 3270 25728 3562
rect 25762 3270 25768 3562
rect 25722 3258 25768 3270
rect 26780 3562 26826 3574
rect 26780 3270 26786 3562
rect 26820 3270 26826 3562
rect 26780 3258 26826 3270
rect 27278 -3192 27574 5224
rect 33848 5230 33896 6426
rect 33990 5230 34144 6426
rect 40304 6426 40638 11138
rect 46836 11160 46956 12356
rect 47050 11160 47170 12356
rect 53442 12370 53776 16706
rect 59628 16980 59698 18464
rect 59892 16980 60012 18464
rect 62112 18636 62158 18648
rect 62112 18344 62118 18636
rect 62152 18344 62158 18636
rect 62112 18332 62158 18344
rect 63170 18636 63216 18648
rect 63170 18344 63176 18636
rect 63210 18344 63216 18636
rect 63170 18332 63216 18344
rect 64228 18636 64274 18648
rect 64228 18344 64234 18636
rect 64268 18344 64274 18636
rect 64228 18332 64274 18344
rect 65286 18636 65332 18648
rect 65286 18344 65292 18636
rect 65326 18344 65332 18636
rect 65286 18332 65332 18344
rect 66344 18636 66390 18648
rect 66344 18344 66350 18636
rect 66384 18344 66390 18636
rect 66344 18332 66390 18344
rect 67402 18636 67448 18648
rect 67402 18344 67408 18636
rect 67442 18344 67448 18636
rect 67402 18332 67448 18344
rect 59628 16702 60012 16980
rect 54086 16478 54132 16490
rect 54086 16186 54092 16478
rect 54126 16186 54132 16478
rect 54086 16174 54132 16186
rect 55144 16478 55190 16490
rect 55144 16186 55150 16478
rect 55184 16186 55190 16478
rect 55144 16174 55190 16186
rect 56202 16478 56248 16490
rect 56202 16186 56208 16478
rect 56242 16186 56248 16478
rect 56202 16174 56248 16186
rect 57260 16478 57306 16490
rect 57260 16186 57266 16478
rect 57300 16186 57306 16478
rect 57260 16174 57306 16186
rect 58318 16478 58364 16490
rect 58318 16186 58324 16478
rect 58358 16186 58364 16478
rect 58318 16174 58364 16186
rect 59376 16478 59422 16490
rect 59376 16186 59382 16478
rect 59416 16186 59422 16478
rect 59376 16174 59422 16186
rect 54086 15384 54132 15396
rect 54086 15092 54092 15384
rect 54126 15092 54132 15384
rect 54086 15080 54132 15092
rect 55144 15384 55190 15396
rect 55144 15092 55150 15384
rect 55184 15092 55190 15384
rect 55144 15080 55190 15092
rect 56202 15384 56248 15396
rect 56202 15092 56208 15384
rect 56242 15092 56248 15384
rect 56202 15080 56248 15092
rect 57260 15384 57306 15396
rect 57260 15092 57266 15384
rect 57300 15092 57306 15384
rect 57260 15080 57306 15092
rect 58318 15384 58364 15396
rect 58318 15092 58324 15384
rect 58358 15092 58364 15384
rect 58318 15080 58364 15092
rect 59376 15384 59422 15396
rect 59376 15092 59382 15384
rect 59416 15092 59422 15384
rect 59376 15080 59422 15092
rect 54096 13904 54142 13916
rect 54096 13612 54102 13904
rect 54136 13612 54142 13904
rect 54096 13600 54142 13612
rect 55154 13904 55200 13916
rect 55154 13612 55160 13904
rect 55194 13612 55200 13904
rect 55154 13600 55200 13612
rect 56212 13904 56258 13916
rect 56212 13612 56218 13904
rect 56252 13612 56258 13904
rect 56212 13600 56258 13612
rect 57270 13904 57316 13916
rect 57270 13612 57276 13904
rect 57310 13612 57316 13904
rect 57270 13600 57316 13612
rect 58328 13904 58374 13916
rect 58328 13612 58334 13904
rect 58368 13612 58374 13904
rect 58328 13600 58374 13612
rect 59386 13904 59432 13916
rect 59386 13612 59392 13904
rect 59426 13612 59432 13904
rect 59386 13600 59432 13612
rect 54096 12810 54142 12822
rect 54096 12518 54102 12810
rect 54136 12518 54142 12810
rect 54096 12506 54142 12518
rect 55154 12810 55200 12822
rect 55154 12518 55160 12810
rect 55194 12518 55200 12810
rect 55154 12506 55200 12518
rect 56212 12810 56258 12822
rect 56212 12518 56218 12810
rect 56252 12518 56258 12810
rect 56212 12506 56258 12518
rect 57270 12810 57316 12822
rect 57270 12518 57276 12810
rect 57310 12518 57316 12810
rect 57270 12506 57316 12518
rect 58328 12810 58374 12822
rect 58328 12518 58334 12810
rect 58368 12518 58374 12810
rect 58328 12506 58374 12518
rect 59386 12810 59432 12822
rect 59386 12518 59392 12810
rect 59426 12518 59432 12810
rect 59680 12694 60012 16702
rect 61464 18196 61614 18322
rect 61464 17000 61486 18196
rect 61580 17000 61614 18196
rect 67596 18208 68186 22836
rect 74374 22810 74636 23606
rect 74730 23606 74764 24006
rect 81076 24004 81226 24130
rect 81076 23754 81098 24004
rect 74730 22810 74964 23606
rect 75262 23352 75308 23364
rect 75262 23060 75268 23352
rect 75302 23060 75308 23352
rect 75262 23048 75308 23060
rect 76320 23352 76366 23364
rect 76320 23060 76326 23352
rect 76360 23060 76366 23352
rect 76320 23048 76366 23060
rect 77378 23352 77424 23364
rect 77378 23060 77384 23352
rect 77418 23060 77424 23352
rect 77378 23048 77424 23060
rect 78436 23352 78482 23364
rect 78436 23060 78442 23352
rect 78476 23060 78482 23352
rect 78436 23048 78482 23060
rect 79494 23352 79540 23364
rect 79494 23060 79500 23352
rect 79534 23060 79540 23352
rect 79494 23048 79540 23060
rect 80552 23352 80598 23364
rect 80552 23060 80558 23352
rect 80592 23060 80598 23352
rect 80552 23048 80598 23060
rect 68568 22284 68614 22296
rect 68568 21992 68574 22284
rect 68608 21992 68614 22284
rect 68568 21980 68614 21992
rect 69626 22284 69672 22296
rect 69626 21992 69632 22284
rect 69666 21992 69672 22284
rect 69626 21980 69672 21992
rect 70684 22284 70730 22296
rect 70684 21992 70690 22284
rect 70724 21992 70730 22284
rect 70684 21980 70730 21992
rect 71742 22284 71788 22296
rect 71742 21992 71748 22284
rect 71782 21992 71788 22284
rect 71742 21980 71788 21992
rect 72800 22284 72846 22296
rect 72800 21992 72806 22284
rect 72840 21992 72846 22284
rect 72800 21980 72846 21992
rect 73858 22284 73904 22296
rect 73858 21992 73864 22284
rect 73898 21992 73904 22284
rect 73858 21980 73904 21992
rect 68568 21190 68614 21202
rect 68568 21066 68574 21190
rect 68562 20898 68574 21066
rect 68608 21066 68614 21190
rect 69626 21190 69672 21202
rect 68608 20898 68662 21066
rect 68562 19742 68662 20898
rect 69626 20898 69632 21190
rect 69666 20898 69672 21190
rect 69626 20886 69672 20898
rect 70684 21190 70730 21202
rect 70684 20898 70690 21190
rect 70724 20898 70730 21190
rect 70684 20886 70730 20898
rect 71742 21190 71788 21202
rect 71742 20898 71748 21190
rect 71782 20898 71788 21190
rect 71742 20886 71788 20898
rect 72800 21190 72846 21202
rect 72800 20898 72806 21190
rect 72840 20898 72846 21190
rect 73858 21190 73904 21202
rect 73858 21132 73864 21190
rect 72800 20886 72846 20898
rect 73822 20898 73864 21132
rect 73898 21132 73904 21190
rect 73898 20898 73954 21132
rect 68562 19614 68582 19742
rect 68576 19450 68582 19614
rect 68616 19614 68662 19742
rect 69634 19742 69680 19754
rect 68616 19450 68622 19614
rect 68576 19438 68622 19450
rect 69634 19450 69640 19742
rect 69674 19450 69680 19742
rect 69634 19438 69680 19450
rect 70692 19742 70738 19754
rect 70692 19450 70698 19742
rect 70732 19450 70738 19742
rect 70692 19438 70738 19450
rect 71750 19742 71796 19754
rect 71750 19450 71756 19742
rect 71790 19450 71796 19742
rect 71750 19438 71796 19450
rect 72808 19742 72854 19754
rect 72808 19450 72814 19742
rect 72848 19450 72854 19742
rect 73822 19742 73954 20898
rect 73822 19636 73872 19742
rect 72808 19438 72854 19450
rect 73866 19450 73872 19636
rect 73906 19636 73954 19742
rect 73906 19450 73912 19636
rect 73866 19438 73912 19450
rect 68576 18648 68622 18660
rect 68576 18356 68582 18648
rect 68616 18356 68622 18648
rect 68576 18344 68622 18356
rect 69634 18648 69680 18660
rect 69634 18356 69640 18648
rect 69674 18356 69680 18648
rect 69634 18344 69680 18356
rect 70692 18648 70738 18660
rect 70692 18356 70698 18648
rect 70732 18356 70738 18648
rect 70692 18344 70738 18356
rect 71750 18648 71796 18660
rect 71750 18356 71756 18648
rect 71790 18356 71796 18648
rect 71750 18344 71796 18356
rect 72808 18648 72854 18660
rect 72808 18356 72814 18648
rect 72848 18356 72854 18648
rect 72808 18344 72854 18356
rect 73866 18648 73912 18660
rect 73866 18356 73872 18648
rect 73906 18356 73912 18648
rect 73866 18344 73912 18356
rect 62112 17542 62158 17554
rect 62112 17250 62118 17542
rect 62152 17250 62158 17542
rect 62112 17238 62158 17250
rect 63170 17542 63216 17554
rect 63170 17250 63176 17542
rect 63210 17250 63216 17542
rect 63170 17238 63216 17250
rect 64228 17542 64274 17554
rect 64228 17250 64234 17542
rect 64268 17250 64274 17542
rect 64228 17238 64274 17250
rect 65286 17542 65332 17554
rect 65286 17250 65292 17542
rect 65326 17250 65332 17542
rect 65286 17238 65332 17250
rect 66344 17542 66390 17554
rect 66344 17250 66350 17542
rect 66384 17250 66390 17542
rect 66344 17238 66390 17250
rect 67402 17542 67448 17554
rect 67402 17250 67408 17542
rect 67442 17250 67448 17542
rect 67402 17238 67448 17250
rect 61464 16676 61614 17000
rect 67596 17012 67950 18208
rect 68044 17012 68186 18208
rect 74374 18168 74964 22810
rect 80820 22808 81098 23754
rect 81192 23754 81226 24004
rect 87848 23998 87998 24124
rect 81192 22808 81372 23754
rect 87848 23606 87870 23998
rect 81724 23350 81770 23362
rect 81724 23058 81730 23350
rect 81764 23058 81770 23350
rect 81724 23046 81770 23058
rect 82782 23350 82828 23362
rect 82782 23058 82788 23350
rect 82822 23058 82828 23350
rect 82782 23046 82828 23058
rect 83840 23350 83886 23362
rect 83840 23058 83846 23350
rect 83880 23058 83886 23350
rect 83840 23046 83886 23058
rect 84898 23350 84944 23362
rect 84898 23058 84904 23350
rect 84938 23058 84944 23350
rect 84898 23046 84944 23058
rect 85956 23350 86002 23362
rect 85956 23058 85962 23350
rect 85996 23058 86002 23350
rect 85956 23046 86002 23058
rect 87014 23350 87060 23362
rect 87014 23058 87020 23350
rect 87054 23058 87060 23350
rect 87014 23046 87060 23058
rect 75262 22258 75308 22270
rect 75262 21966 75268 22258
rect 75302 21966 75308 22258
rect 75262 21954 75308 21966
rect 76320 22258 76366 22270
rect 76320 21966 76326 22258
rect 76360 21966 76366 22258
rect 76320 21954 76366 21966
rect 77378 22258 77424 22270
rect 77378 21966 77384 22258
rect 77418 21966 77424 22258
rect 77378 21954 77424 21966
rect 78436 22258 78482 22270
rect 78436 21966 78442 22258
rect 78476 21966 78482 22258
rect 78436 21954 78482 21966
rect 79494 22258 79540 22270
rect 79494 21966 79500 22258
rect 79534 21966 79540 22258
rect 79494 21954 79540 21966
rect 80552 22258 80598 22270
rect 80552 21966 80558 22258
rect 80592 21966 80598 22258
rect 80552 21954 80598 21966
rect 75262 21164 75308 21176
rect 75262 20984 75268 21164
rect 75236 20872 75268 20984
rect 75302 20984 75308 21164
rect 76320 21164 76366 21176
rect 75302 20872 75336 20984
rect 75236 19702 75336 20872
rect 76320 20872 76326 21164
rect 76360 20872 76366 21164
rect 76320 20860 76366 20872
rect 77378 21164 77424 21176
rect 77378 20872 77384 21164
rect 77418 20872 77424 21164
rect 77378 20860 77424 20872
rect 78436 21164 78482 21176
rect 78436 20872 78442 21164
rect 78476 20872 78482 21164
rect 78436 20860 78482 20872
rect 79494 21164 79540 21176
rect 79494 20872 79500 21164
rect 79534 20872 79540 21164
rect 80552 21164 80598 21176
rect 80552 21016 80558 21164
rect 79494 20860 79540 20872
rect 80530 20872 80558 21016
rect 80592 21016 80598 21164
rect 80592 20872 80630 21016
rect 75236 19532 75274 19702
rect 75268 19410 75274 19532
rect 75308 19532 75336 19702
rect 76326 19702 76372 19714
rect 75308 19410 75314 19532
rect 75268 19398 75314 19410
rect 76326 19410 76332 19702
rect 76366 19410 76372 19702
rect 76326 19398 76372 19410
rect 77384 19702 77430 19714
rect 77384 19410 77390 19702
rect 77424 19410 77430 19702
rect 77384 19398 77430 19410
rect 78442 19702 78488 19714
rect 78442 19410 78448 19702
rect 78482 19410 78488 19702
rect 78442 19398 78488 19410
rect 79500 19702 79546 19714
rect 79500 19410 79506 19702
rect 79540 19410 79546 19702
rect 80530 19702 80630 20872
rect 80530 19564 80564 19702
rect 79500 19398 79546 19410
rect 80558 19410 80564 19564
rect 80598 19564 80630 19702
rect 80598 19410 80604 19564
rect 80558 19398 80604 19410
rect 75268 18608 75314 18620
rect 75268 18316 75274 18608
rect 75308 18316 75314 18608
rect 75268 18304 75314 18316
rect 76326 18608 76372 18620
rect 76326 18316 76332 18608
rect 76366 18316 76372 18608
rect 76326 18304 76372 18316
rect 77384 18608 77430 18620
rect 77384 18316 77390 18608
rect 77424 18316 77430 18608
rect 77384 18304 77430 18316
rect 78442 18608 78488 18620
rect 78442 18316 78448 18608
rect 78482 18316 78488 18608
rect 78442 18304 78488 18316
rect 79500 18608 79546 18620
rect 79500 18316 79506 18608
rect 79540 18316 79546 18608
rect 79500 18304 79546 18316
rect 80558 18608 80604 18620
rect 80558 18316 80564 18608
rect 80598 18316 80604 18608
rect 80558 18304 80604 18316
rect 68576 17554 68622 17566
rect 68576 17262 68582 17554
rect 68616 17262 68622 17554
rect 68576 17250 68622 17262
rect 69634 17554 69680 17566
rect 69634 17262 69640 17554
rect 69674 17262 69680 17554
rect 69634 17250 69680 17262
rect 70692 17554 70738 17566
rect 70692 17262 70698 17554
rect 70732 17262 70738 17554
rect 70692 17250 70738 17262
rect 71750 17554 71796 17566
rect 71750 17262 71756 17554
rect 71790 17262 71796 17554
rect 71750 17250 71796 17262
rect 72808 17554 72854 17566
rect 72808 17262 72814 17554
rect 72848 17262 72854 17554
rect 72808 17250 72854 17262
rect 73866 17554 73912 17566
rect 73866 17262 73872 17554
rect 73906 17262 73912 17554
rect 73866 17250 73912 17262
rect 62112 16448 62158 16460
rect 62112 16156 62118 16448
rect 62152 16156 62158 16448
rect 62112 16144 62158 16156
rect 63170 16448 63216 16460
rect 63170 16156 63176 16448
rect 63210 16156 63216 16448
rect 63170 16144 63216 16156
rect 64228 16448 64274 16460
rect 64228 16156 64234 16448
rect 64268 16156 64274 16448
rect 64228 16144 64274 16156
rect 65286 16448 65332 16460
rect 65286 16156 65292 16448
rect 65326 16156 65332 16448
rect 65286 16144 65332 16156
rect 66344 16448 66390 16460
rect 66344 16156 66350 16448
rect 66384 16156 66390 16448
rect 66344 16144 66390 16156
rect 67402 16448 67448 16460
rect 67402 16156 67408 16448
rect 67442 16156 67448 16448
rect 67402 16144 67448 16156
rect 62112 15354 62158 15366
rect 62112 15146 62118 15354
rect 62080 15062 62118 15146
rect 62152 15146 62158 15354
rect 63170 15354 63216 15366
rect 62152 15062 62180 15146
rect 62080 13872 62180 15062
rect 63170 15062 63176 15354
rect 63210 15062 63216 15354
rect 63170 15050 63216 15062
rect 64228 15354 64274 15366
rect 64228 15062 64234 15354
rect 64268 15062 64274 15354
rect 64228 15050 64274 15062
rect 65286 15354 65332 15366
rect 65286 15062 65292 15354
rect 65326 15062 65332 15354
rect 65286 15050 65332 15062
rect 66344 15354 66390 15366
rect 66344 15062 66350 15354
rect 66384 15062 66390 15354
rect 67402 15354 67448 15366
rect 67402 15212 67408 15354
rect 66344 15050 66390 15062
rect 67374 15062 67408 15212
rect 67442 15212 67448 15354
rect 67442 15062 67474 15212
rect 62080 13694 62118 13872
rect 62112 13580 62118 13694
rect 62152 13694 62180 13872
rect 63170 13872 63216 13884
rect 62152 13580 62158 13694
rect 62112 13568 62158 13580
rect 63170 13580 63176 13872
rect 63210 13580 63216 13872
rect 63170 13568 63216 13580
rect 64228 13872 64274 13884
rect 64228 13580 64234 13872
rect 64268 13580 64274 13872
rect 64228 13568 64274 13580
rect 65286 13872 65332 13884
rect 65286 13580 65292 13872
rect 65326 13580 65332 13872
rect 65286 13568 65332 13580
rect 66344 13872 66390 13884
rect 66344 13580 66350 13872
rect 66384 13580 66390 13872
rect 67374 13872 67474 15062
rect 67374 13760 67408 13872
rect 66344 13568 66390 13580
rect 67402 13580 67408 13760
rect 67442 13760 67474 13872
rect 67442 13580 67448 13760
rect 67402 13568 67448 13580
rect 59386 12506 59432 12518
rect 59642 12542 60012 12694
rect 47582 11702 47628 11714
rect 47582 11410 47588 11702
rect 47622 11410 47628 11702
rect 47582 11398 47628 11410
rect 48640 11702 48686 11714
rect 48640 11410 48646 11702
rect 48680 11410 48686 11702
rect 48640 11398 48686 11410
rect 49698 11702 49744 11714
rect 49698 11410 49704 11702
rect 49738 11410 49744 11702
rect 49698 11398 49744 11410
rect 50756 11702 50802 11714
rect 50756 11410 50762 11702
rect 50796 11410 50802 11702
rect 50756 11398 50802 11410
rect 51814 11702 51860 11714
rect 51814 11410 51820 11702
rect 51854 11410 51860 11702
rect 51814 11398 51860 11410
rect 52872 11702 52918 11714
rect 52872 11410 52878 11702
rect 52912 11410 52918 11702
rect 52872 11398 52918 11410
rect 40994 10586 41040 10598
rect 40994 10294 41000 10586
rect 41034 10294 41040 10586
rect 40994 10282 41040 10294
rect 42052 10586 42098 10598
rect 42052 10294 42058 10586
rect 42092 10294 42098 10586
rect 42052 10282 42098 10294
rect 43110 10586 43156 10598
rect 43110 10294 43116 10586
rect 43150 10294 43156 10586
rect 43110 10282 43156 10294
rect 44168 10586 44214 10598
rect 44168 10294 44174 10586
rect 44208 10294 44214 10586
rect 44168 10282 44214 10294
rect 45226 10586 45272 10598
rect 45226 10294 45232 10586
rect 45266 10294 45272 10586
rect 45226 10282 45272 10294
rect 46284 10586 46330 10598
rect 46284 10294 46290 10586
rect 46324 10294 46330 10586
rect 46284 10282 46330 10294
rect 40994 9492 41040 9504
rect 40994 9200 41000 9492
rect 41034 9200 41040 9492
rect 40994 9188 41040 9200
rect 42052 9492 42098 9504
rect 42052 9200 42058 9492
rect 42092 9200 42098 9492
rect 42052 9188 42098 9200
rect 43110 9492 43156 9504
rect 43110 9200 43116 9492
rect 43150 9200 43156 9492
rect 43110 9188 43156 9200
rect 44168 9492 44214 9504
rect 44168 9200 44174 9492
rect 44208 9200 44214 9492
rect 44168 9188 44214 9200
rect 45226 9492 45272 9504
rect 45226 9200 45232 9492
rect 45266 9200 45272 9492
rect 45226 9188 45272 9200
rect 46284 9492 46330 9504
rect 46284 9200 46290 9492
rect 46324 9200 46330 9492
rect 46284 9188 46330 9200
rect 41012 7960 41058 7972
rect 41012 7668 41018 7960
rect 41052 7668 41058 7960
rect 41012 7656 41058 7668
rect 42070 7960 42116 7972
rect 42070 7668 42076 7960
rect 42110 7668 42116 7960
rect 42070 7656 42116 7668
rect 43128 7960 43174 7972
rect 43128 7668 43134 7960
rect 43168 7668 43174 7960
rect 43128 7656 43174 7668
rect 44186 7960 44232 7972
rect 44186 7668 44192 7960
rect 44226 7668 44232 7960
rect 44186 7656 44232 7668
rect 45244 7960 45290 7972
rect 45244 7668 45250 7960
rect 45284 7668 45290 7960
rect 45244 7656 45290 7668
rect 46302 7960 46348 7972
rect 46302 7668 46308 7960
rect 46342 7668 46348 7960
rect 46302 7656 46348 7668
rect 41012 6866 41058 6878
rect 41012 6574 41018 6866
rect 41052 6574 41058 6866
rect 41012 6562 41058 6574
rect 42070 6866 42116 6878
rect 42070 6574 42076 6866
rect 42110 6574 42116 6866
rect 42070 6562 42116 6574
rect 43128 6866 43174 6878
rect 43128 6574 43134 6866
rect 43168 6574 43174 6866
rect 43128 6562 43174 6574
rect 44186 6866 44232 6878
rect 44186 6574 44192 6866
rect 44226 6574 44232 6866
rect 44186 6562 44232 6574
rect 45244 6866 45290 6878
rect 45244 6574 45250 6866
rect 45284 6574 45290 6866
rect 45244 6562 45290 6574
rect 46302 6866 46348 6878
rect 46302 6574 46308 6866
rect 46342 6574 46348 6866
rect 46302 6562 46348 6574
rect 34522 5772 34568 5784
rect 34522 5480 34528 5772
rect 34562 5480 34568 5772
rect 34522 5468 34568 5480
rect 35580 5772 35626 5784
rect 35580 5480 35586 5772
rect 35620 5480 35626 5772
rect 35580 5468 35626 5480
rect 36638 5772 36684 5784
rect 36638 5480 36644 5772
rect 36678 5480 36684 5772
rect 36638 5468 36684 5480
rect 37696 5772 37742 5784
rect 37696 5480 37702 5772
rect 37736 5480 37742 5772
rect 37696 5468 37742 5480
rect 38754 5772 38800 5784
rect 38754 5480 38760 5772
rect 38794 5480 38800 5772
rect 38754 5468 38800 5480
rect 39812 5772 39858 5784
rect 39812 5480 39818 5772
rect 39852 5480 39858 5772
rect 40304 5642 40386 6426
rect 39812 5468 39858 5480
rect 28012 4672 28058 4684
rect 28012 4380 28018 4672
rect 28052 4380 28058 4672
rect 28012 4368 28058 4380
rect 29070 4672 29116 4684
rect 29070 4380 29076 4672
rect 29110 4380 29116 4672
rect 29070 4368 29116 4380
rect 30128 4672 30174 4684
rect 30128 4380 30134 4672
rect 30168 4380 30174 4672
rect 30128 4368 30174 4380
rect 31186 4672 31232 4684
rect 31186 4380 31192 4672
rect 31226 4380 31232 4672
rect 31186 4368 31232 4380
rect 32244 4672 32290 4684
rect 32244 4380 32250 4672
rect 32284 4380 32290 4672
rect 32244 4368 32290 4380
rect 33302 4672 33348 4684
rect 33302 4380 33308 4672
rect 33342 4380 33348 4672
rect 33302 4368 33348 4380
rect 28012 3578 28058 3590
rect 28012 3286 28018 3578
rect 28052 3286 28058 3578
rect 28012 3274 28058 3286
rect 29070 3578 29116 3590
rect 29070 3286 29076 3578
rect 29110 3286 29116 3578
rect 29070 3274 29116 3286
rect 30128 3578 30174 3590
rect 30128 3286 30134 3578
rect 30168 3286 30174 3578
rect 30128 3274 30174 3286
rect 31186 3578 31232 3590
rect 31186 3286 31192 3578
rect 31226 3286 31232 3578
rect 31186 3274 31232 3286
rect 32244 3578 32290 3590
rect 32244 3286 32250 3578
rect 32284 3286 32290 3578
rect 32244 3274 32290 3286
rect 33302 3578 33348 3590
rect 33302 3286 33308 3578
rect 33342 3286 33348 3578
rect 33302 3274 33348 3286
rect 33848 -3192 34144 5230
rect 40364 5230 40386 5642
rect 40480 5642 40638 6426
rect 46836 6448 47170 11160
rect 53442 11174 53470 12370
rect 53564 11174 53776 12370
rect 54096 11716 54142 11728
rect 54096 11424 54102 11716
rect 54136 11424 54142 11716
rect 54096 11412 54142 11424
rect 55154 11716 55200 11728
rect 55154 11424 55160 11716
rect 55194 11424 55200 11716
rect 55154 11412 55200 11424
rect 56212 11716 56258 11728
rect 56212 11424 56218 11716
rect 56252 11424 56258 11716
rect 56212 11412 56258 11424
rect 57270 11716 57316 11728
rect 57270 11424 57276 11716
rect 57310 11424 57316 11716
rect 57270 11412 57316 11424
rect 58328 11716 58374 11728
rect 58328 11424 58334 11716
rect 58368 11424 58374 11716
rect 58328 11412 58374 11424
rect 59386 11716 59432 11728
rect 59386 11424 59392 11716
rect 59426 11424 59432 11716
rect 59386 11412 59432 11424
rect 47582 10608 47628 10620
rect 47582 10316 47588 10608
rect 47622 10316 47628 10608
rect 47582 10304 47628 10316
rect 48640 10608 48686 10620
rect 48640 10316 48646 10608
rect 48680 10316 48686 10608
rect 48640 10304 48686 10316
rect 49698 10608 49744 10620
rect 49698 10316 49704 10608
rect 49738 10316 49744 10608
rect 49698 10304 49744 10316
rect 50756 10608 50802 10620
rect 50756 10316 50762 10608
rect 50796 10316 50802 10608
rect 50756 10304 50802 10316
rect 51814 10608 51860 10620
rect 51814 10316 51820 10608
rect 51854 10316 51860 10608
rect 51814 10304 51860 10316
rect 52872 10608 52918 10620
rect 52872 10316 52878 10608
rect 52912 10316 52918 10608
rect 52872 10304 52918 10316
rect 47582 9514 47628 9526
rect 47582 9222 47588 9514
rect 47622 9222 47628 9514
rect 47582 9210 47628 9222
rect 48640 9514 48686 9526
rect 48640 9222 48646 9514
rect 48680 9222 48686 9514
rect 48640 9210 48686 9222
rect 49698 9514 49744 9526
rect 49698 9222 49704 9514
rect 49738 9222 49744 9514
rect 49698 9210 49744 9222
rect 50756 9514 50802 9526
rect 50756 9222 50762 9514
rect 50796 9222 50802 9514
rect 50756 9210 50802 9222
rect 51814 9514 51860 9526
rect 51814 9222 51820 9514
rect 51854 9222 51860 9514
rect 51814 9210 51860 9222
rect 52872 9514 52918 9526
rect 52872 9222 52878 9514
rect 52912 9222 52918 9514
rect 52872 9210 52918 9222
rect 47600 7982 47646 7994
rect 47600 7690 47606 7982
rect 47640 7690 47646 7982
rect 47600 7678 47646 7690
rect 48658 7982 48704 7994
rect 48658 7690 48664 7982
rect 48698 7690 48704 7982
rect 48658 7678 48704 7690
rect 49716 7982 49762 7994
rect 49716 7690 49722 7982
rect 49756 7690 49762 7982
rect 49716 7678 49762 7690
rect 50774 7982 50820 7994
rect 50774 7690 50780 7982
rect 50814 7690 50820 7982
rect 50774 7678 50820 7690
rect 51832 7982 51878 7994
rect 51832 7690 51838 7982
rect 51872 7690 51878 7982
rect 51832 7678 51878 7690
rect 52890 7982 52936 7994
rect 52890 7690 52896 7982
rect 52930 7690 52936 7982
rect 52890 7678 52936 7690
rect 47600 6888 47646 6900
rect 47600 6596 47606 6888
rect 47640 6596 47646 6888
rect 47600 6584 47646 6596
rect 48658 6888 48704 6900
rect 48658 6596 48664 6888
rect 48698 6596 48704 6888
rect 48658 6584 48704 6596
rect 49716 6888 49762 6900
rect 49716 6596 49722 6888
rect 49756 6596 49762 6888
rect 49716 6584 49762 6596
rect 50774 6888 50820 6900
rect 50774 6596 50780 6888
rect 50814 6596 50820 6888
rect 50774 6584 50820 6596
rect 51832 6888 51878 6900
rect 51832 6596 51838 6888
rect 51872 6596 51878 6888
rect 51832 6584 51878 6596
rect 52890 6888 52936 6900
rect 52890 6596 52896 6888
rect 52930 6596 52936 6888
rect 52890 6584 52936 6596
rect 41012 5772 41058 5784
rect 40480 5230 40514 5642
rect 41012 5480 41018 5772
rect 41052 5480 41058 5772
rect 41012 5468 41058 5480
rect 42070 5772 42116 5784
rect 42070 5480 42076 5772
rect 42110 5480 42116 5772
rect 42070 5468 42116 5480
rect 43128 5772 43174 5784
rect 43128 5480 43134 5772
rect 43168 5480 43174 5772
rect 43128 5468 43174 5480
rect 44186 5772 44232 5784
rect 44186 5480 44192 5772
rect 44226 5480 44232 5772
rect 44186 5468 44232 5480
rect 45244 5772 45290 5784
rect 45244 5480 45250 5772
rect 45284 5480 45290 5772
rect 45244 5468 45290 5480
rect 46302 5772 46348 5784
rect 46302 5480 46308 5772
rect 46342 5480 46348 5772
rect 46302 5468 46348 5480
rect 46836 5344 46974 6448
rect 40364 4906 40514 5230
rect 46952 5252 46974 5344
rect 47068 5684 47170 6448
rect 53442 6462 53776 11174
rect 59642 11168 59698 12542
rect 59934 11168 60012 12542
rect 62112 12778 62158 12790
rect 62112 12486 62118 12778
rect 62152 12486 62158 12778
rect 62112 12474 62158 12486
rect 63170 12778 63216 12790
rect 63170 12486 63176 12778
rect 63210 12486 63216 12778
rect 63170 12474 63216 12486
rect 64228 12778 64274 12790
rect 64228 12486 64234 12778
rect 64268 12486 64274 12778
rect 64228 12474 64274 12486
rect 65286 12778 65332 12790
rect 65286 12486 65292 12778
rect 65326 12486 65332 12778
rect 65286 12474 65332 12486
rect 66344 12778 66390 12790
rect 66344 12486 66350 12778
rect 66384 12486 66390 12778
rect 66344 12474 66390 12486
rect 67402 12778 67448 12790
rect 67402 12486 67408 12778
rect 67442 12486 67448 12778
rect 67402 12474 67448 12486
rect 59642 11002 60012 11168
rect 54096 10622 54142 10634
rect 54096 10330 54102 10622
rect 54136 10330 54142 10622
rect 54096 10318 54142 10330
rect 55154 10622 55200 10634
rect 55154 10330 55160 10622
rect 55194 10330 55200 10622
rect 55154 10318 55200 10330
rect 56212 10622 56258 10634
rect 56212 10330 56218 10622
rect 56252 10330 56258 10622
rect 56212 10318 56258 10330
rect 57270 10622 57316 10634
rect 57270 10330 57276 10622
rect 57310 10330 57316 10622
rect 57270 10318 57316 10330
rect 58328 10622 58374 10634
rect 58328 10330 58334 10622
rect 58368 10330 58374 10622
rect 58328 10318 58374 10330
rect 59386 10622 59432 10634
rect 59386 10330 59392 10622
rect 59426 10330 59432 10622
rect 59386 10318 59432 10330
rect 54096 9528 54142 9540
rect 54096 9236 54102 9528
rect 54136 9236 54142 9528
rect 54096 9224 54142 9236
rect 55154 9528 55200 9540
rect 55154 9236 55160 9528
rect 55194 9236 55200 9528
rect 55154 9224 55200 9236
rect 56212 9528 56258 9540
rect 56212 9236 56218 9528
rect 56252 9236 56258 9528
rect 56212 9224 56258 9236
rect 57270 9528 57316 9540
rect 57270 9236 57276 9528
rect 57310 9236 57316 9528
rect 57270 9224 57316 9236
rect 58328 9528 58374 9540
rect 58328 9236 58334 9528
rect 58368 9236 58374 9528
rect 58328 9224 58374 9236
rect 59386 9528 59432 9540
rect 59386 9236 59392 9528
rect 59426 9236 59432 9528
rect 59386 9224 59432 9236
rect 54114 7996 54160 8008
rect 54114 7704 54120 7996
rect 54154 7704 54160 7996
rect 54114 7692 54160 7704
rect 55172 7996 55218 8008
rect 55172 7704 55178 7996
rect 55212 7704 55218 7996
rect 55172 7692 55218 7704
rect 56230 7996 56276 8008
rect 56230 7704 56236 7996
rect 56270 7704 56276 7996
rect 56230 7692 56276 7704
rect 57288 7996 57334 8008
rect 57288 7704 57294 7996
rect 57328 7704 57334 7996
rect 57288 7692 57334 7704
rect 58346 7996 58392 8008
rect 58346 7704 58352 7996
rect 58386 7704 58392 7996
rect 58346 7692 58392 7704
rect 59404 7996 59450 8008
rect 59404 7704 59410 7996
rect 59444 7704 59450 7996
rect 59404 7692 59450 7704
rect 54114 6902 54160 6914
rect 54114 6610 54120 6902
rect 54154 6610 54160 6902
rect 54114 6598 54160 6610
rect 55172 6902 55218 6914
rect 55172 6610 55178 6902
rect 55212 6610 55218 6902
rect 55172 6598 55218 6610
rect 56230 6902 56276 6914
rect 56230 6610 56236 6902
rect 56270 6610 56276 6902
rect 56230 6598 56276 6610
rect 57288 6902 57334 6914
rect 57288 6610 57294 6902
rect 57328 6610 57334 6902
rect 57288 6598 57334 6610
rect 58346 6902 58392 6914
rect 58346 6610 58352 6902
rect 58386 6610 58392 6902
rect 58346 6598 58392 6610
rect 59404 6902 59450 6914
rect 59404 6610 59410 6902
rect 59444 6610 59450 6902
rect 59680 6812 60012 11002
rect 61464 12338 61614 12464
rect 61464 11142 61486 12338
rect 61580 11142 61614 12338
rect 67596 12336 68186 17012
rect 74374 16972 74642 18168
rect 74736 16972 74964 18168
rect 80820 18180 81372 22808
rect 87672 22802 87870 23606
rect 87964 23606 87998 23998
rect 94310 23996 94460 24122
rect 87964 22802 88224 23606
rect 88496 23344 88542 23356
rect 88496 23052 88502 23344
rect 88536 23052 88542 23344
rect 88496 23040 88542 23052
rect 89554 23344 89600 23356
rect 89554 23052 89560 23344
rect 89594 23052 89600 23344
rect 89554 23040 89600 23052
rect 90612 23344 90658 23356
rect 90612 23052 90618 23344
rect 90652 23052 90658 23344
rect 90612 23040 90658 23052
rect 91670 23344 91716 23356
rect 91670 23052 91676 23344
rect 91710 23052 91716 23344
rect 91670 23040 91716 23052
rect 92728 23344 92774 23356
rect 92728 23052 92734 23344
rect 92768 23052 92774 23344
rect 92728 23040 92774 23052
rect 93786 23344 93832 23356
rect 94310 23348 94332 23996
rect 93786 23052 93792 23344
rect 93826 23052 93832 23344
rect 93786 23040 93832 23052
rect 81724 22256 81770 22268
rect 81724 21964 81730 22256
rect 81764 21964 81770 22256
rect 81724 21952 81770 21964
rect 82782 22256 82828 22268
rect 82782 21964 82788 22256
rect 82822 21964 82828 22256
rect 82782 21952 82828 21964
rect 83840 22256 83886 22268
rect 83840 21964 83846 22256
rect 83880 21964 83886 22256
rect 83840 21952 83886 21964
rect 84898 22256 84944 22268
rect 84898 21964 84904 22256
rect 84938 21964 84944 22256
rect 84898 21952 84944 21964
rect 85956 22256 86002 22268
rect 85956 21964 85962 22256
rect 85996 21964 86002 22256
rect 85956 21952 86002 21964
rect 87014 22256 87060 22268
rect 87014 21964 87020 22256
rect 87054 21964 87060 22256
rect 87014 21952 87060 21964
rect 81724 21162 81770 21174
rect 81724 21038 81730 21162
rect 81718 20870 81730 21038
rect 81764 21038 81770 21162
rect 82782 21162 82828 21174
rect 81764 20870 81818 21038
rect 81718 19714 81818 20870
rect 82782 20870 82788 21162
rect 82822 20870 82828 21162
rect 82782 20858 82828 20870
rect 83840 21162 83886 21174
rect 83840 20870 83846 21162
rect 83880 20870 83886 21162
rect 83840 20858 83886 20870
rect 84898 21162 84944 21174
rect 84898 20870 84904 21162
rect 84938 20870 84944 21162
rect 84898 20858 84944 20870
rect 85956 21162 86002 21174
rect 85956 20870 85962 21162
rect 85996 20870 86002 21162
rect 87014 21162 87060 21174
rect 87014 21104 87020 21162
rect 85956 20858 86002 20870
rect 86978 20870 87020 21104
rect 87054 21104 87060 21162
rect 87054 20870 87110 21104
rect 81718 19586 81738 19714
rect 81732 19422 81738 19586
rect 81772 19586 81818 19714
rect 82790 19714 82836 19726
rect 81772 19422 81778 19586
rect 81732 19410 81778 19422
rect 82790 19422 82796 19714
rect 82830 19422 82836 19714
rect 82790 19410 82836 19422
rect 83848 19714 83894 19726
rect 83848 19422 83854 19714
rect 83888 19422 83894 19714
rect 83848 19410 83894 19422
rect 84906 19714 84952 19726
rect 84906 19422 84912 19714
rect 84946 19422 84952 19714
rect 84906 19410 84952 19422
rect 85964 19714 86010 19726
rect 85964 19422 85970 19714
rect 86004 19422 86010 19714
rect 86978 19714 87110 20870
rect 86978 19608 87028 19714
rect 85964 19410 86010 19422
rect 87022 19422 87028 19608
rect 87062 19608 87110 19714
rect 87062 19422 87068 19608
rect 87022 19410 87068 19422
rect 81732 18620 81778 18632
rect 81732 18328 81738 18620
rect 81772 18328 81778 18620
rect 81732 18316 81778 18328
rect 82790 18620 82836 18632
rect 82790 18328 82796 18620
rect 82830 18328 82836 18620
rect 82790 18316 82836 18328
rect 83848 18620 83894 18632
rect 83848 18328 83854 18620
rect 83888 18328 83894 18620
rect 83848 18316 83894 18328
rect 84906 18620 84952 18632
rect 84906 18328 84912 18620
rect 84946 18328 84952 18620
rect 84906 18316 84952 18328
rect 85964 18620 86010 18632
rect 85964 18328 85970 18620
rect 86004 18328 86010 18620
rect 85964 18316 86010 18328
rect 87022 18620 87068 18632
rect 87022 18328 87028 18620
rect 87062 18328 87068 18620
rect 87022 18316 87068 18328
rect 75268 17514 75314 17526
rect 75268 17222 75274 17514
rect 75308 17222 75314 17514
rect 75268 17210 75314 17222
rect 76326 17514 76372 17526
rect 76326 17222 76332 17514
rect 76366 17222 76372 17514
rect 76326 17210 76372 17222
rect 77384 17514 77430 17526
rect 77384 17222 77390 17514
rect 77424 17222 77430 17514
rect 77384 17210 77430 17222
rect 78442 17514 78488 17526
rect 78442 17222 78448 17514
rect 78482 17222 78488 17514
rect 78442 17210 78488 17222
rect 79500 17514 79546 17526
rect 79500 17222 79506 17514
rect 79540 17222 79546 17514
rect 79500 17210 79546 17222
rect 80558 17514 80604 17526
rect 80558 17222 80564 17514
rect 80598 17222 80604 17514
rect 80558 17210 80604 17222
rect 68576 16460 68622 16472
rect 68576 16168 68582 16460
rect 68616 16168 68622 16460
rect 68576 16156 68622 16168
rect 69634 16460 69680 16472
rect 69634 16168 69640 16460
rect 69674 16168 69680 16460
rect 69634 16156 69680 16168
rect 70692 16460 70738 16472
rect 70692 16168 70698 16460
rect 70732 16168 70738 16460
rect 70692 16156 70738 16168
rect 71750 16460 71796 16472
rect 71750 16168 71756 16460
rect 71790 16168 71796 16460
rect 71750 16156 71796 16168
rect 72808 16460 72854 16472
rect 72808 16168 72814 16460
rect 72848 16168 72854 16460
rect 72808 16156 72854 16168
rect 73866 16460 73912 16472
rect 73866 16168 73872 16460
rect 73906 16168 73912 16460
rect 73866 16156 73912 16168
rect 68576 15366 68622 15378
rect 68576 15180 68582 15366
rect 68518 15074 68582 15180
rect 68616 15074 68622 15366
rect 68518 15062 68622 15074
rect 69634 15366 69680 15378
rect 69634 15074 69640 15366
rect 69674 15074 69680 15366
rect 69634 15062 69680 15074
rect 70692 15366 70738 15378
rect 70692 15074 70698 15366
rect 70732 15074 70738 15366
rect 70692 15062 70738 15074
rect 71750 15366 71796 15378
rect 71750 15074 71756 15366
rect 71790 15074 71796 15366
rect 71750 15062 71796 15074
rect 72808 15366 72854 15378
rect 72808 15074 72814 15366
rect 72848 15074 72854 15366
rect 73866 15366 73912 15378
rect 73866 15180 73872 15366
rect 72808 15062 72854 15074
rect 73800 15074 73872 15180
rect 73906 15180 73912 15366
rect 73906 15074 73932 15180
rect 68518 13882 68618 15062
rect 68518 13870 68626 13882
rect 68518 13728 68586 13870
rect 68580 13578 68586 13728
rect 68620 13578 68626 13870
rect 68580 13566 68626 13578
rect 69638 13870 69684 13882
rect 69638 13578 69644 13870
rect 69678 13578 69684 13870
rect 69638 13566 69684 13578
rect 70696 13870 70742 13882
rect 70696 13578 70702 13870
rect 70736 13578 70742 13870
rect 70696 13566 70742 13578
rect 71754 13870 71800 13882
rect 71754 13578 71760 13870
rect 71794 13578 71800 13870
rect 71754 13566 71800 13578
rect 72812 13870 72858 13882
rect 72812 13578 72818 13870
rect 72852 13578 72858 13870
rect 73800 13870 73932 15074
rect 73800 13684 73876 13870
rect 72812 13566 72858 13578
rect 73870 13578 73876 13684
rect 73910 13684 73932 13870
rect 73910 13578 73916 13684
rect 73870 13566 73916 13578
rect 68580 12776 68626 12788
rect 68580 12484 68586 12776
rect 68620 12484 68626 12776
rect 68580 12472 68626 12484
rect 69638 12776 69684 12788
rect 69638 12484 69644 12776
rect 69678 12484 69684 12776
rect 69638 12472 69684 12484
rect 70696 12776 70742 12788
rect 70696 12484 70702 12776
rect 70736 12484 70742 12776
rect 70696 12472 70742 12484
rect 71754 12776 71800 12788
rect 71754 12484 71760 12776
rect 71794 12484 71800 12776
rect 71754 12472 71800 12484
rect 72812 12776 72858 12788
rect 72812 12484 72818 12776
rect 72852 12484 72858 12776
rect 72812 12472 72858 12484
rect 73870 12776 73916 12788
rect 73870 12484 73876 12776
rect 73910 12484 73916 12776
rect 73870 12472 73916 12484
rect 62112 11684 62158 11696
rect 62112 11392 62118 11684
rect 62152 11392 62158 11684
rect 62112 11380 62158 11392
rect 63170 11684 63216 11696
rect 63170 11392 63176 11684
rect 63210 11392 63216 11684
rect 63170 11380 63216 11392
rect 64228 11684 64274 11696
rect 64228 11392 64234 11684
rect 64268 11392 64274 11684
rect 64228 11380 64274 11392
rect 65286 11684 65332 11696
rect 65286 11392 65292 11684
rect 65326 11392 65332 11684
rect 65286 11380 65332 11392
rect 66344 11684 66390 11696
rect 66344 11392 66350 11684
rect 66384 11392 66390 11684
rect 66344 11380 66390 11392
rect 67402 11684 67448 11696
rect 67402 11392 67408 11684
rect 67442 11392 67448 11684
rect 67402 11380 67448 11392
rect 61464 10818 61614 11142
rect 67596 11140 67954 12336
rect 68048 11140 68186 12336
rect 74374 12310 74964 16972
rect 80820 16984 81106 18180
rect 81200 16984 81372 18180
rect 87672 18160 88224 22802
rect 94120 22800 94332 23348
rect 94426 23348 94460 23996
rect 94426 22800 94672 23348
rect 94958 23342 95004 23354
rect 94958 23050 94964 23342
rect 94998 23050 95004 23342
rect 94958 23038 95004 23050
rect 96016 23342 96062 23354
rect 96016 23050 96022 23342
rect 96056 23050 96062 23342
rect 96016 23038 96062 23050
rect 97074 23342 97120 23354
rect 97074 23050 97080 23342
rect 97114 23050 97120 23342
rect 97074 23038 97120 23050
rect 98132 23342 98178 23354
rect 98132 23050 98138 23342
rect 98172 23050 98178 23342
rect 98132 23038 98178 23050
rect 99190 23342 99236 23354
rect 99190 23050 99196 23342
rect 99230 23050 99236 23342
rect 99190 23038 99236 23050
rect 100248 23342 100294 23354
rect 100248 23050 100254 23342
rect 100288 23050 100294 23342
rect 100248 23038 100294 23050
rect 88496 22250 88542 22262
rect 88496 21958 88502 22250
rect 88536 21958 88542 22250
rect 88496 21946 88542 21958
rect 89554 22250 89600 22262
rect 89554 21958 89560 22250
rect 89594 21958 89600 22250
rect 89554 21946 89600 21958
rect 90612 22250 90658 22262
rect 90612 21958 90618 22250
rect 90652 21958 90658 22250
rect 90612 21946 90658 21958
rect 91670 22250 91716 22262
rect 91670 21958 91676 22250
rect 91710 21958 91716 22250
rect 91670 21946 91716 21958
rect 92728 22250 92774 22262
rect 92728 21958 92734 22250
rect 92768 21958 92774 22250
rect 92728 21946 92774 21958
rect 93786 22250 93832 22262
rect 93786 21958 93792 22250
rect 93826 21958 93832 22250
rect 93786 21946 93832 21958
rect 88496 21156 88542 21168
rect 88496 20976 88502 21156
rect 88470 20864 88502 20976
rect 88536 20976 88542 21156
rect 89554 21156 89600 21168
rect 88536 20864 88570 20976
rect 88470 19694 88570 20864
rect 89554 20864 89560 21156
rect 89594 20864 89600 21156
rect 89554 20852 89600 20864
rect 90612 21156 90658 21168
rect 90612 20864 90618 21156
rect 90652 20864 90658 21156
rect 90612 20852 90658 20864
rect 91670 21156 91716 21168
rect 91670 20864 91676 21156
rect 91710 20864 91716 21156
rect 91670 20852 91716 20864
rect 92728 21156 92774 21168
rect 92728 20864 92734 21156
rect 92768 20864 92774 21156
rect 93786 21156 93832 21168
rect 93786 21008 93792 21156
rect 92728 20852 92774 20864
rect 93764 20864 93792 21008
rect 93826 21008 93832 21156
rect 93826 20864 93864 21008
rect 88470 19524 88508 19694
rect 88502 19402 88508 19524
rect 88542 19524 88570 19694
rect 89560 19694 89606 19706
rect 88542 19402 88548 19524
rect 88502 19390 88548 19402
rect 89560 19402 89566 19694
rect 89600 19402 89606 19694
rect 89560 19390 89606 19402
rect 90618 19694 90664 19706
rect 90618 19402 90624 19694
rect 90658 19402 90664 19694
rect 90618 19390 90664 19402
rect 91676 19694 91722 19706
rect 91676 19402 91682 19694
rect 91716 19402 91722 19694
rect 91676 19390 91722 19402
rect 92734 19694 92780 19706
rect 92734 19402 92740 19694
rect 92774 19402 92780 19694
rect 93764 19694 93864 20864
rect 93764 19556 93798 19694
rect 92734 19390 92780 19402
rect 93792 19402 93798 19556
rect 93832 19556 93864 19694
rect 93832 19402 93838 19556
rect 93792 19390 93838 19402
rect 88502 18600 88548 18612
rect 88502 18308 88508 18600
rect 88542 18308 88548 18600
rect 88502 18296 88548 18308
rect 89560 18600 89606 18612
rect 89560 18308 89566 18600
rect 89600 18308 89606 18600
rect 89560 18296 89606 18308
rect 90618 18600 90664 18612
rect 90618 18308 90624 18600
rect 90658 18308 90664 18600
rect 90618 18296 90664 18308
rect 91676 18600 91722 18612
rect 91676 18308 91682 18600
rect 91716 18308 91722 18600
rect 91676 18296 91722 18308
rect 92734 18600 92780 18612
rect 92734 18308 92740 18600
rect 92774 18308 92780 18600
rect 92734 18296 92780 18308
rect 93792 18600 93838 18612
rect 93792 18308 93798 18600
rect 93832 18308 93838 18600
rect 93792 18296 93838 18308
rect 81732 17526 81778 17538
rect 81732 17234 81738 17526
rect 81772 17234 81778 17526
rect 81732 17222 81778 17234
rect 82790 17526 82836 17538
rect 82790 17234 82796 17526
rect 82830 17234 82836 17526
rect 82790 17222 82836 17234
rect 83848 17526 83894 17538
rect 83848 17234 83854 17526
rect 83888 17234 83894 17526
rect 83848 17222 83894 17234
rect 84906 17526 84952 17538
rect 84906 17234 84912 17526
rect 84946 17234 84952 17526
rect 84906 17222 84952 17234
rect 85964 17526 86010 17538
rect 85964 17234 85970 17526
rect 86004 17234 86010 17526
rect 85964 17222 86010 17234
rect 87022 17526 87068 17538
rect 87022 17234 87028 17526
rect 87062 17234 87068 17526
rect 87022 17222 87068 17234
rect 75268 16420 75314 16432
rect 75268 16128 75274 16420
rect 75308 16128 75314 16420
rect 75268 16116 75314 16128
rect 76326 16420 76372 16432
rect 76326 16128 76332 16420
rect 76366 16128 76372 16420
rect 76326 16116 76372 16128
rect 77384 16420 77430 16432
rect 77384 16128 77390 16420
rect 77424 16128 77430 16420
rect 77384 16116 77430 16128
rect 78442 16420 78488 16432
rect 78442 16128 78448 16420
rect 78482 16128 78488 16420
rect 78442 16116 78488 16128
rect 79500 16420 79546 16432
rect 79500 16128 79506 16420
rect 79540 16128 79546 16420
rect 79500 16116 79546 16128
rect 80558 16420 80604 16432
rect 80558 16128 80564 16420
rect 80598 16128 80604 16420
rect 80558 16116 80604 16128
rect 75268 15326 75314 15338
rect 75268 15118 75274 15326
rect 75236 15034 75274 15118
rect 75308 15118 75314 15326
rect 76326 15326 76372 15338
rect 75308 15034 75336 15118
rect 75236 13844 75336 15034
rect 76326 15034 76332 15326
rect 76366 15034 76372 15326
rect 76326 15022 76372 15034
rect 77384 15326 77430 15338
rect 77384 15034 77390 15326
rect 77424 15034 77430 15326
rect 77384 15022 77430 15034
rect 78442 15326 78488 15338
rect 78442 15034 78448 15326
rect 78482 15034 78488 15326
rect 78442 15022 78488 15034
rect 79500 15326 79546 15338
rect 79500 15034 79506 15326
rect 79540 15034 79546 15326
rect 80558 15326 80604 15338
rect 80558 15184 80564 15326
rect 79500 15022 79546 15034
rect 80530 15034 80564 15184
rect 80598 15184 80604 15326
rect 80598 15034 80630 15184
rect 75236 13666 75274 13844
rect 75268 13552 75274 13666
rect 75308 13666 75336 13844
rect 76326 13844 76372 13856
rect 75308 13552 75314 13666
rect 75268 13540 75314 13552
rect 76326 13552 76332 13844
rect 76366 13552 76372 13844
rect 76326 13540 76372 13552
rect 77384 13844 77430 13856
rect 77384 13552 77390 13844
rect 77424 13552 77430 13844
rect 77384 13540 77430 13552
rect 78442 13844 78488 13856
rect 78442 13552 78448 13844
rect 78482 13552 78488 13844
rect 78442 13540 78488 13552
rect 79500 13844 79546 13856
rect 79500 13552 79506 13844
rect 79540 13552 79546 13844
rect 80530 13844 80630 15034
rect 80530 13732 80564 13844
rect 79500 13540 79546 13552
rect 80558 13552 80564 13732
rect 80598 13732 80630 13844
rect 80598 13552 80604 13732
rect 80558 13540 80604 13552
rect 75268 12750 75314 12762
rect 75268 12458 75274 12750
rect 75308 12458 75314 12750
rect 75268 12446 75314 12458
rect 76326 12750 76372 12762
rect 76326 12458 76332 12750
rect 76366 12458 76372 12750
rect 76326 12446 76372 12458
rect 77384 12750 77430 12762
rect 77384 12458 77390 12750
rect 77424 12458 77430 12750
rect 77384 12446 77430 12458
rect 78442 12750 78488 12762
rect 78442 12458 78448 12750
rect 78482 12458 78488 12750
rect 78442 12446 78488 12458
rect 79500 12750 79546 12762
rect 79500 12458 79506 12750
rect 79540 12458 79546 12750
rect 79500 12446 79546 12458
rect 80558 12750 80604 12762
rect 80558 12458 80564 12750
rect 80598 12458 80604 12750
rect 80558 12446 80604 12458
rect 68580 11682 68626 11694
rect 68580 11390 68586 11682
rect 68620 11390 68626 11682
rect 68580 11378 68626 11390
rect 69638 11682 69684 11694
rect 69638 11390 69644 11682
rect 69678 11390 69684 11682
rect 69638 11378 69684 11390
rect 70696 11682 70742 11694
rect 70696 11390 70702 11682
rect 70736 11390 70742 11682
rect 70696 11378 70742 11390
rect 71754 11682 71800 11694
rect 71754 11390 71760 11682
rect 71794 11390 71800 11682
rect 71754 11378 71800 11390
rect 72812 11682 72858 11694
rect 72812 11390 72818 11682
rect 72852 11390 72858 11682
rect 72812 11378 72858 11390
rect 73870 11682 73916 11694
rect 73870 11390 73876 11682
rect 73910 11390 73916 11682
rect 73870 11378 73916 11390
rect 62112 10590 62158 10602
rect 62112 10298 62118 10590
rect 62152 10298 62158 10590
rect 62112 10286 62158 10298
rect 63170 10590 63216 10602
rect 63170 10298 63176 10590
rect 63210 10298 63216 10590
rect 63170 10286 63216 10298
rect 64228 10590 64274 10602
rect 64228 10298 64234 10590
rect 64268 10298 64274 10590
rect 64228 10286 64274 10298
rect 65286 10590 65332 10602
rect 65286 10298 65292 10590
rect 65326 10298 65332 10590
rect 65286 10286 65332 10298
rect 66344 10590 66390 10602
rect 66344 10298 66350 10590
rect 66384 10298 66390 10590
rect 66344 10286 66390 10298
rect 67402 10590 67448 10602
rect 67402 10298 67408 10590
rect 67442 10298 67448 10590
rect 67402 10286 67448 10298
rect 62112 9496 62158 9508
rect 62112 9292 62118 9496
rect 62092 9204 62118 9292
rect 62152 9292 62158 9496
rect 63170 9496 63216 9508
rect 62152 9204 62192 9292
rect 62092 8014 62192 9204
rect 63170 9204 63176 9496
rect 63210 9204 63216 9496
rect 63170 9192 63216 9204
rect 64228 9496 64274 9508
rect 64228 9204 64234 9496
rect 64268 9204 64274 9496
rect 64228 9192 64274 9204
rect 65286 9496 65332 9508
rect 65286 9204 65292 9496
rect 65326 9204 65332 9496
rect 65286 9192 65332 9204
rect 66344 9496 66390 9508
rect 66344 9204 66350 9496
rect 66384 9204 66390 9496
rect 67402 9496 67448 9508
rect 67402 9326 67408 9496
rect 66344 9192 66390 9204
rect 67362 9204 67408 9326
rect 67442 9326 67448 9496
rect 67442 9204 67462 9326
rect 62092 7840 62118 8014
rect 62112 7722 62118 7840
rect 62152 7840 62192 8014
rect 63170 8014 63216 8026
rect 62152 7722 62158 7840
rect 62112 7710 62158 7722
rect 63170 7722 63176 8014
rect 63210 7722 63216 8014
rect 63170 7710 63216 7722
rect 64228 8014 64274 8026
rect 64228 7722 64234 8014
rect 64268 7722 64274 8014
rect 64228 7710 64274 7722
rect 65286 8014 65332 8026
rect 65286 7722 65292 8014
rect 65326 7722 65332 8014
rect 65286 7710 65332 7722
rect 66344 8014 66390 8026
rect 66344 7722 66350 8014
rect 66384 7722 66390 8014
rect 67362 8014 67462 9204
rect 67362 7874 67408 8014
rect 66344 7710 66390 7722
rect 67402 7722 67408 7874
rect 67442 7874 67462 8014
rect 67442 7722 67448 7874
rect 67402 7710 67448 7722
rect 59404 6598 59450 6610
rect 59600 6714 60012 6812
rect 47600 5794 47646 5806
rect 47600 5684 47606 5794
rect 47068 5502 47606 5684
rect 47640 5684 47646 5794
rect 48658 5794 48704 5806
rect 47640 5502 47736 5684
rect 47068 5478 47736 5502
rect 48658 5502 48664 5794
rect 48698 5502 48704 5794
rect 48658 5490 48704 5502
rect 49716 5794 49762 5806
rect 49716 5502 49722 5794
rect 49756 5502 49762 5794
rect 49716 5490 49762 5502
rect 50774 5794 50820 5806
rect 50774 5502 50780 5794
rect 50814 5502 50820 5794
rect 50774 5490 50820 5502
rect 51832 5794 51878 5806
rect 51832 5502 51838 5794
rect 51872 5502 51878 5794
rect 51832 5490 51878 5502
rect 52890 5794 52936 5806
rect 52890 5502 52896 5794
rect 52930 5502 52936 5794
rect 53442 5720 53488 6462
rect 53392 5514 53488 5720
rect 52890 5490 52936 5502
rect 53442 5494 53488 5514
rect 47068 5344 47170 5478
rect 47068 5252 47102 5344
rect 46952 4928 47102 5252
rect 53466 5266 53488 5494
rect 53582 5720 53776 6462
rect 54114 5808 54160 5820
rect 54114 5720 54120 5808
rect 53582 5516 54120 5720
rect 54154 5720 54160 5808
rect 55172 5808 55218 5820
rect 54154 5516 54196 5720
rect 53582 5514 54196 5516
rect 55172 5516 55178 5808
rect 55212 5516 55218 5808
rect 53582 5494 53776 5514
rect 54114 5504 54160 5514
rect 55172 5504 55218 5516
rect 56230 5808 56276 5820
rect 56230 5516 56236 5808
rect 56270 5516 56276 5808
rect 56230 5504 56276 5516
rect 57288 5808 57334 5820
rect 57288 5516 57294 5808
rect 57328 5516 57334 5808
rect 57288 5504 57334 5516
rect 58346 5808 58392 5820
rect 58346 5516 58352 5808
rect 58386 5516 58392 5808
rect 59404 5808 59450 5820
rect 59404 5702 59410 5808
rect 58346 5504 58392 5516
rect 59364 5516 59410 5702
rect 59444 5702 59450 5808
rect 59600 5702 59684 6714
rect 59444 5516 59684 5702
rect 53582 5266 53616 5494
rect 59364 5478 59684 5516
rect 53466 4942 53616 5266
rect 59600 5340 59684 5478
rect 59850 5340 60012 6714
rect 62112 6920 62158 6932
rect 62112 6628 62118 6920
rect 62152 6628 62158 6920
rect 62112 6616 62158 6628
rect 63170 6920 63216 6932
rect 63170 6628 63176 6920
rect 63210 6628 63216 6920
rect 63170 6616 63216 6628
rect 64228 6920 64274 6932
rect 64228 6628 64234 6920
rect 64268 6628 64274 6920
rect 64228 6616 64274 6628
rect 65286 6920 65332 6932
rect 65286 6628 65292 6920
rect 65326 6628 65332 6920
rect 65286 6616 65332 6628
rect 66344 6920 66390 6932
rect 66344 6628 66350 6920
rect 66384 6628 66390 6920
rect 66344 6616 66390 6628
rect 67402 6920 67448 6932
rect 67402 6628 67408 6920
rect 67442 6628 67448 6920
rect 67402 6616 67448 6628
rect 59600 5174 60012 5340
rect 54114 4714 54160 4726
rect 47600 4700 47646 4712
rect 34522 4678 34568 4690
rect 34522 4386 34528 4678
rect 34562 4386 34568 4678
rect 34522 4374 34568 4386
rect 35580 4678 35626 4690
rect 35580 4386 35586 4678
rect 35620 4386 35626 4678
rect 35580 4374 35626 4386
rect 36638 4678 36684 4690
rect 36638 4386 36644 4678
rect 36678 4386 36684 4678
rect 36638 4374 36684 4386
rect 37696 4678 37742 4690
rect 37696 4386 37702 4678
rect 37736 4386 37742 4678
rect 37696 4374 37742 4386
rect 38754 4678 38800 4690
rect 38754 4386 38760 4678
rect 38794 4386 38800 4678
rect 38754 4374 38800 4386
rect 39812 4678 39858 4690
rect 39812 4386 39818 4678
rect 39852 4386 39858 4678
rect 39812 4374 39858 4386
rect 41012 4678 41058 4690
rect 41012 4386 41018 4678
rect 41052 4386 41058 4678
rect 41012 4374 41058 4386
rect 42070 4678 42116 4690
rect 42070 4386 42076 4678
rect 42110 4386 42116 4678
rect 42070 4374 42116 4386
rect 43128 4678 43174 4690
rect 43128 4386 43134 4678
rect 43168 4386 43174 4678
rect 43128 4374 43174 4386
rect 44186 4678 44232 4690
rect 44186 4386 44192 4678
rect 44226 4386 44232 4678
rect 44186 4374 44232 4386
rect 45244 4678 45290 4690
rect 45244 4386 45250 4678
rect 45284 4386 45290 4678
rect 45244 4374 45290 4386
rect 46302 4678 46348 4690
rect 46302 4386 46308 4678
rect 46342 4386 46348 4678
rect 47600 4408 47606 4700
rect 47640 4408 47646 4700
rect 47600 4396 47646 4408
rect 48658 4700 48704 4712
rect 48658 4408 48664 4700
rect 48698 4408 48704 4700
rect 48658 4396 48704 4408
rect 49716 4700 49762 4712
rect 49716 4408 49722 4700
rect 49756 4408 49762 4700
rect 49716 4396 49762 4408
rect 50774 4700 50820 4712
rect 50774 4408 50780 4700
rect 50814 4408 50820 4700
rect 50774 4396 50820 4408
rect 51832 4700 51878 4712
rect 51832 4408 51838 4700
rect 51872 4408 51878 4700
rect 51832 4396 51878 4408
rect 52890 4700 52936 4712
rect 52890 4408 52896 4700
rect 52930 4408 52936 4700
rect 54114 4422 54120 4714
rect 54154 4422 54160 4714
rect 54114 4410 54160 4422
rect 55172 4714 55218 4726
rect 55172 4422 55178 4714
rect 55212 4422 55218 4714
rect 55172 4410 55218 4422
rect 56230 4714 56276 4726
rect 56230 4422 56236 4714
rect 56270 4422 56276 4714
rect 56230 4410 56276 4422
rect 57288 4714 57334 4726
rect 57288 4422 57294 4714
rect 57328 4422 57334 4714
rect 57288 4410 57334 4422
rect 58346 4714 58392 4726
rect 58346 4422 58352 4714
rect 58386 4422 58392 4714
rect 58346 4410 58392 4422
rect 59404 4714 59450 4726
rect 59404 4422 59410 4714
rect 59444 4422 59450 4714
rect 59404 4410 59450 4422
rect 52890 4396 52936 4408
rect 46302 4374 46348 4386
rect 54114 3620 54160 3632
rect 47600 3606 47646 3618
rect 34522 3584 34568 3596
rect 34522 3292 34528 3584
rect 34562 3292 34568 3584
rect 34522 3280 34568 3292
rect 35580 3584 35626 3596
rect 35580 3292 35586 3584
rect 35620 3292 35626 3584
rect 35580 3280 35626 3292
rect 36638 3584 36684 3596
rect 36638 3292 36644 3584
rect 36678 3292 36684 3584
rect 36638 3280 36684 3292
rect 37696 3584 37742 3596
rect 37696 3292 37702 3584
rect 37736 3292 37742 3584
rect 37696 3280 37742 3292
rect 38754 3584 38800 3596
rect 38754 3292 38760 3584
rect 38794 3292 38800 3584
rect 39812 3584 39858 3596
rect 39812 3390 39818 3584
rect 38754 3280 38800 3292
rect 39690 3292 39818 3390
rect 39852 3390 39858 3584
rect 41012 3584 41058 3596
rect 39852 3292 39982 3390
rect 39690 2594 39982 3292
rect 41012 3292 41018 3584
rect 41052 3292 41058 3584
rect 41012 3280 41058 3292
rect 42070 3584 42116 3596
rect 42070 3292 42076 3584
rect 42110 3292 42116 3584
rect 42070 3280 42116 3292
rect 43128 3584 43174 3596
rect 43128 3292 43134 3584
rect 43168 3292 43174 3584
rect 43128 3280 43174 3292
rect 44186 3584 44232 3596
rect 44186 3292 44192 3584
rect 44226 3292 44232 3584
rect 44186 3280 44232 3292
rect 45244 3584 45290 3596
rect 45244 3292 45250 3584
rect 45284 3292 45290 3584
rect 45244 3280 45290 3292
rect 46302 3584 46348 3596
rect 46302 3292 46308 3584
rect 46342 3292 46348 3584
rect 47600 3314 47606 3606
rect 47640 3314 47646 3606
rect 47600 3302 47646 3314
rect 48658 3606 48704 3618
rect 48658 3314 48664 3606
rect 48698 3314 48704 3606
rect 48658 3302 48704 3314
rect 49716 3606 49762 3618
rect 49716 3314 49722 3606
rect 49756 3314 49762 3606
rect 49716 3302 49762 3314
rect 50774 3606 50820 3618
rect 50774 3314 50780 3606
rect 50814 3314 50820 3606
rect 50774 3302 50820 3314
rect 51832 3606 51878 3618
rect 51832 3314 51838 3606
rect 51872 3314 51878 3606
rect 51832 3302 51878 3314
rect 52890 3606 52936 3618
rect 52890 3314 52896 3606
rect 52930 3314 52936 3606
rect 54114 3328 54120 3620
rect 54154 3328 54160 3620
rect 54114 3316 54160 3328
rect 55172 3620 55218 3632
rect 55172 3328 55178 3620
rect 55212 3328 55218 3620
rect 55172 3316 55218 3328
rect 56230 3620 56276 3632
rect 56230 3328 56236 3620
rect 56270 3328 56276 3620
rect 56230 3316 56276 3328
rect 57288 3620 57334 3632
rect 57288 3328 57294 3620
rect 57328 3328 57334 3620
rect 57288 3316 57334 3328
rect 58346 3620 58392 3632
rect 58346 3328 58352 3620
rect 58386 3328 58392 3620
rect 58346 3316 58392 3328
rect 59404 3620 59450 3632
rect 59404 3328 59410 3620
rect 59444 3328 59450 3620
rect 59680 3574 60012 5174
rect 61464 6480 61614 6606
rect 61464 5284 61486 6480
rect 61580 5284 61614 6480
rect 67596 6478 68186 11140
rect 74374 11114 74642 12310
rect 74736 11114 74964 12310
rect 80820 12308 81372 16984
rect 87672 16964 87876 18160
rect 87970 16964 88224 18160
rect 94120 18172 94672 22800
rect 94958 22248 95004 22260
rect 94958 21956 94964 22248
rect 94998 21956 95004 22248
rect 94958 21944 95004 21956
rect 96016 22248 96062 22260
rect 96016 21956 96022 22248
rect 96056 21956 96062 22248
rect 96016 21944 96062 21956
rect 97074 22248 97120 22260
rect 97074 21956 97080 22248
rect 97114 21956 97120 22248
rect 97074 21944 97120 21956
rect 98132 22248 98178 22260
rect 98132 21956 98138 22248
rect 98172 21956 98178 22248
rect 98132 21944 98178 21956
rect 99190 22248 99236 22260
rect 99190 21956 99196 22248
rect 99230 21956 99236 22248
rect 99190 21944 99236 21956
rect 100248 22248 100294 22260
rect 100248 21956 100254 22248
rect 100288 21956 100294 22248
rect 100248 21944 100294 21956
rect 100676 21760 100786 24224
rect 101276 22686 101320 25032
rect 101276 21760 101376 22686
rect 94958 21154 95004 21166
rect 94958 21030 94964 21154
rect 94952 20862 94964 21030
rect 94998 21030 95004 21154
rect 96016 21154 96062 21166
rect 94998 20862 95052 21030
rect 94952 19706 95052 20862
rect 96016 20862 96022 21154
rect 96056 20862 96062 21154
rect 96016 20850 96062 20862
rect 97074 21154 97120 21166
rect 97074 20862 97080 21154
rect 97114 20862 97120 21154
rect 97074 20850 97120 20862
rect 98132 21154 98178 21166
rect 98132 20862 98138 21154
rect 98172 20862 98178 21154
rect 98132 20850 98178 20862
rect 99190 21154 99236 21166
rect 99190 20862 99196 21154
rect 99230 20862 99236 21154
rect 100248 21154 100294 21166
rect 100248 21096 100254 21154
rect 99190 20850 99236 20862
rect 100212 20862 100254 21096
rect 100288 21096 100294 21154
rect 100288 20862 100344 21096
rect 100676 21046 101376 21760
rect 94952 19578 94972 19706
rect 94966 19414 94972 19578
rect 95006 19578 95052 19706
rect 96024 19706 96070 19718
rect 95006 19414 95012 19578
rect 94966 19402 95012 19414
rect 96024 19414 96030 19706
rect 96064 19414 96070 19706
rect 96024 19402 96070 19414
rect 97082 19706 97128 19718
rect 97082 19414 97088 19706
rect 97122 19414 97128 19706
rect 97082 19402 97128 19414
rect 98140 19706 98186 19718
rect 98140 19414 98146 19706
rect 98180 19414 98186 19706
rect 98140 19402 98186 19414
rect 99198 19706 99244 19718
rect 99198 19414 99204 19706
rect 99238 19414 99244 19706
rect 100212 19706 100344 20862
rect 100212 19600 100262 19706
rect 99198 19402 99244 19414
rect 100256 19414 100262 19600
rect 100296 19600 100344 19706
rect 100296 19414 100302 19600
rect 100256 19402 100302 19414
rect 100788 19266 101376 21046
rect 100630 18976 101376 19266
rect 94966 18612 95012 18624
rect 94966 18320 94972 18612
rect 95006 18320 95012 18612
rect 94966 18308 95012 18320
rect 96024 18612 96070 18624
rect 96024 18320 96030 18612
rect 96064 18320 96070 18612
rect 96024 18308 96070 18320
rect 97082 18612 97128 18624
rect 97082 18320 97088 18612
rect 97122 18320 97128 18612
rect 97082 18308 97128 18320
rect 98140 18612 98186 18624
rect 98140 18320 98146 18612
rect 98180 18320 98186 18612
rect 98140 18308 98186 18320
rect 99198 18612 99244 18624
rect 99198 18320 99204 18612
rect 99238 18320 99244 18612
rect 99198 18308 99244 18320
rect 100256 18612 100302 18624
rect 100256 18320 100262 18612
rect 100296 18320 100302 18612
rect 100256 18308 100302 18320
rect 88502 17506 88548 17518
rect 88502 17214 88508 17506
rect 88542 17214 88548 17506
rect 88502 17202 88548 17214
rect 89560 17506 89606 17518
rect 89560 17214 89566 17506
rect 89600 17214 89606 17506
rect 89560 17202 89606 17214
rect 90618 17506 90664 17518
rect 90618 17214 90624 17506
rect 90658 17214 90664 17506
rect 90618 17202 90664 17214
rect 91676 17506 91722 17518
rect 91676 17214 91682 17506
rect 91716 17214 91722 17506
rect 91676 17202 91722 17214
rect 92734 17506 92780 17518
rect 92734 17214 92740 17506
rect 92774 17214 92780 17506
rect 92734 17202 92780 17214
rect 93792 17506 93838 17518
rect 93792 17214 93798 17506
rect 93832 17214 93838 17506
rect 93792 17202 93838 17214
rect 81732 16432 81778 16444
rect 81732 16140 81738 16432
rect 81772 16140 81778 16432
rect 81732 16128 81778 16140
rect 82790 16432 82836 16444
rect 82790 16140 82796 16432
rect 82830 16140 82836 16432
rect 82790 16128 82836 16140
rect 83848 16432 83894 16444
rect 83848 16140 83854 16432
rect 83888 16140 83894 16432
rect 83848 16128 83894 16140
rect 84906 16432 84952 16444
rect 84906 16140 84912 16432
rect 84946 16140 84952 16432
rect 84906 16128 84952 16140
rect 85964 16432 86010 16444
rect 85964 16140 85970 16432
rect 86004 16140 86010 16432
rect 85964 16128 86010 16140
rect 87022 16432 87068 16444
rect 87022 16140 87028 16432
rect 87062 16140 87068 16432
rect 87022 16128 87068 16140
rect 81732 15338 81778 15350
rect 81732 15152 81738 15338
rect 81674 15046 81738 15152
rect 81772 15046 81778 15338
rect 81674 15034 81778 15046
rect 82790 15338 82836 15350
rect 82790 15046 82796 15338
rect 82830 15046 82836 15338
rect 82790 15034 82836 15046
rect 83848 15338 83894 15350
rect 83848 15046 83854 15338
rect 83888 15046 83894 15338
rect 83848 15034 83894 15046
rect 84906 15338 84952 15350
rect 84906 15046 84912 15338
rect 84946 15046 84952 15338
rect 84906 15034 84952 15046
rect 85964 15338 86010 15350
rect 85964 15046 85970 15338
rect 86004 15046 86010 15338
rect 87022 15338 87068 15350
rect 87022 15152 87028 15338
rect 85964 15034 86010 15046
rect 86956 15046 87028 15152
rect 87062 15152 87068 15338
rect 87062 15046 87088 15152
rect 81674 13854 81774 15034
rect 81674 13842 81782 13854
rect 81674 13700 81742 13842
rect 81736 13550 81742 13700
rect 81776 13550 81782 13842
rect 81736 13538 81782 13550
rect 82794 13842 82840 13854
rect 82794 13550 82800 13842
rect 82834 13550 82840 13842
rect 82794 13538 82840 13550
rect 83852 13842 83898 13854
rect 83852 13550 83858 13842
rect 83892 13550 83898 13842
rect 83852 13538 83898 13550
rect 84910 13842 84956 13854
rect 84910 13550 84916 13842
rect 84950 13550 84956 13842
rect 84910 13538 84956 13550
rect 85968 13842 86014 13854
rect 85968 13550 85974 13842
rect 86008 13550 86014 13842
rect 86956 13842 87088 15046
rect 86956 13656 87032 13842
rect 85968 13538 86014 13550
rect 87026 13550 87032 13656
rect 87066 13656 87088 13842
rect 87066 13550 87072 13656
rect 87026 13538 87072 13550
rect 81736 12748 81782 12760
rect 81736 12456 81742 12748
rect 81776 12456 81782 12748
rect 81736 12444 81782 12456
rect 82794 12748 82840 12760
rect 82794 12456 82800 12748
rect 82834 12456 82840 12748
rect 82794 12444 82840 12456
rect 83852 12748 83898 12760
rect 83852 12456 83858 12748
rect 83892 12456 83898 12748
rect 83852 12444 83898 12456
rect 84910 12748 84956 12760
rect 84910 12456 84916 12748
rect 84950 12456 84956 12748
rect 84910 12444 84956 12456
rect 85968 12748 86014 12760
rect 85968 12456 85974 12748
rect 86008 12456 86014 12748
rect 85968 12444 86014 12456
rect 87026 12748 87072 12760
rect 87026 12456 87032 12748
rect 87066 12456 87072 12748
rect 87026 12444 87072 12456
rect 75268 11656 75314 11668
rect 75268 11364 75274 11656
rect 75308 11364 75314 11656
rect 75268 11352 75314 11364
rect 76326 11656 76372 11668
rect 76326 11364 76332 11656
rect 76366 11364 76372 11656
rect 76326 11352 76372 11364
rect 77384 11656 77430 11668
rect 77384 11364 77390 11656
rect 77424 11364 77430 11656
rect 77384 11352 77430 11364
rect 78442 11656 78488 11668
rect 78442 11364 78448 11656
rect 78482 11364 78488 11656
rect 78442 11352 78488 11364
rect 79500 11656 79546 11668
rect 79500 11364 79506 11656
rect 79540 11364 79546 11656
rect 79500 11352 79546 11364
rect 80558 11656 80604 11668
rect 80558 11364 80564 11656
rect 80598 11364 80604 11656
rect 80558 11352 80604 11364
rect 68580 10588 68626 10600
rect 68580 10296 68586 10588
rect 68620 10296 68626 10588
rect 68580 10284 68626 10296
rect 69638 10588 69684 10600
rect 69638 10296 69644 10588
rect 69678 10296 69684 10588
rect 69638 10284 69684 10296
rect 70696 10588 70742 10600
rect 70696 10296 70702 10588
rect 70736 10296 70742 10588
rect 70696 10284 70742 10296
rect 71754 10588 71800 10600
rect 71754 10296 71760 10588
rect 71794 10296 71800 10588
rect 71754 10284 71800 10296
rect 72812 10588 72858 10600
rect 72812 10296 72818 10588
rect 72852 10296 72858 10588
rect 72812 10284 72858 10296
rect 73870 10588 73916 10600
rect 73870 10296 73876 10588
rect 73910 10296 73916 10588
rect 73870 10284 73916 10296
rect 68580 9494 68626 9506
rect 68580 9348 68586 9494
rect 68550 9202 68586 9348
rect 68620 9348 68626 9494
rect 69638 9494 69684 9506
rect 68620 9202 68650 9348
rect 68550 8012 68650 9202
rect 69638 9202 69644 9494
rect 69678 9202 69684 9494
rect 69638 9190 69684 9202
rect 70696 9494 70742 9506
rect 70696 9202 70702 9494
rect 70736 9202 70742 9494
rect 70696 9190 70742 9202
rect 71754 9494 71800 9506
rect 71754 9202 71760 9494
rect 71794 9202 71800 9494
rect 71754 9190 71800 9202
rect 72812 9494 72858 9506
rect 72812 9202 72818 9494
rect 72852 9202 72858 9494
rect 73870 9494 73916 9506
rect 73870 9424 73876 9494
rect 72812 9190 72858 9202
rect 73832 9202 73876 9424
rect 73910 9424 73916 9494
rect 73910 9202 73964 9424
rect 68550 7896 68590 8012
rect 68584 7720 68590 7896
rect 68624 7896 68650 8012
rect 69642 8012 69688 8024
rect 68624 7720 68630 7896
rect 68584 7708 68630 7720
rect 69642 7720 69648 8012
rect 69682 7720 69688 8012
rect 69642 7708 69688 7720
rect 70700 8012 70746 8024
rect 70700 7720 70706 8012
rect 70740 7720 70746 8012
rect 70700 7708 70746 7720
rect 71758 8012 71804 8024
rect 71758 7720 71764 8012
rect 71798 7720 71804 8012
rect 71758 7708 71804 7720
rect 72816 8012 72862 8024
rect 72816 7720 72822 8012
rect 72856 7720 72862 8012
rect 73832 8012 73964 9202
rect 73832 7928 73880 8012
rect 72816 7708 72862 7720
rect 73874 7720 73880 7928
rect 73914 7928 73964 8012
rect 73914 7720 73920 7928
rect 73874 7708 73920 7720
rect 68584 6918 68630 6930
rect 68584 6626 68590 6918
rect 68624 6626 68630 6918
rect 68584 6614 68630 6626
rect 69642 6918 69688 6930
rect 69642 6626 69648 6918
rect 69682 6626 69688 6918
rect 69642 6614 69688 6626
rect 70700 6918 70746 6930
rect 70700 6626 70706 6918
rect 70740 6626 70746 6918
rect 70700 6614 70746 6626
rect 71758 6918 71804 6930
rect 71758 6626 71764 6918
rect 71798 6626 71804 6918
rect 71758 6614 71804 6626
rect 72816 6918 72862 6930
rect 72816 6626 72822 6918
rect 72856 6626 72862 6918
rect 72816 6614 72862 6626
rect 73874 6918 73920 6930
rect 73874 6626 73880 6918
rect 73914 6626 73920 6918
rect 73874 6614 73920 6626
rect 62112 5826 62158 5838
rect 62112 5534 62118 5826
rect 62152 5534 62158 5826
rect 62112 5522 62158 5534
rect 63170 5826 63216 5838
rect 63170 5534 63176 5826
rect 63210 5534 63216 5826
rect 63170 5522 63216 5534
rect 64228 5826 64274 5838
rect 64228 5534 64234 5826
rect 64268 5534 64274 5826
rect 64228 5522 64274 5534
rect 65286 5826 65332 5838
rect 65286 5534 65292 5826
rect 65326 5534 65332 5826
rect 65286 5522 65332 5534
rect 66344 5826 66390 5838
rect 66344 5534 66350 5826
rect 66384 5534 66390 5826
rect 66344 5522 66390 5534
rect 67402 5826 67448 5838
rect 67402 5534 67408 5826
rect 67442 5534 67448 5826
rect 67596 5592 67958 6478
rect 67402 5522 67448 5534
rect 61464 4960 61614 5284
rect 67936 5282 67958 5592
rect 68052 5592 68186 6478
rect 74374 6452 74964 11114
rect 80820 11112 81110 12308
rect 81204 11112 81372 12308
rect 87672 12302 88224 16964
rect 94120 16976 94340 18172
rect 94434 16976 94672 18172
rect 94966 17518 95012 17530
rect 94966 17226 94972 17518
rect 95006 17226 95012 17518
rect 94966 17214 95012 17226
rect 96024 17518 96070 17530
rect 96024 17226 96030 17518
rect 96064 17226 96070 17518
rect 96024 17214 96070 17226
rect 97082 17518 97128 17530
rect 97082 17226 97088 17518
rect 97122 17226 97128 17518
rect 97082 17214 97128 17226
rect 98140 17518 98186 17530
rect 98140 17226 98146 17518
rect 98180 17226 98186 17518
rect 98140 17214 98186 17226
rect 99198 17518 99244 17530
rect 99198 17226 99204 17518
rect 99238 17226 99244 17518
rect 99198 17214 99244 17226
rect 100256 17518 100302 17530
rect 100256 17226 100262 17518
rect 100296 17226 100302 17518
rect 100256 17214 100302 17226
rect 88502 16412 88548 16424
rect 88502 16120 88508 16412
rect 88542 16120 88548 16412
rect 88502 16108 88548 16120
rect 89560 16412 89606 16424
rect 89560 16120 89566 16412
rect 89600 16120 89606 16412
rect 89560 16108 89606 16120
rect 90618 16412 90664 16424
rect 90618 16120 90624 16412
rect 90658 16120 90664 16412
rect 90618 16108 90664 16120
rect 91676 16412 91722 16424
rect 91676 16120 91682 16412
rect 91716 16120 91722 16412
rect 91676 16108 91722 16120
rect 92734 16412 92780 16424
rect 92734 16120 92740 16412
rect 92774 16120 92780 16412
rect 92734 16108 92780 16120
rect 93792 16412 93838 16424
rect 93792 16120 93798 16412
rect 93832 16120 93838 16412
rect 93792 16108 93838 16120
rect 88502 15318 88548 15330
rect 88502 15110 88508 15318
rect 88470 15026 88508 15110
rect 88542 15110 88548 15318
rect 89560 15318 89606 15330
rect 88542 15026 88570 15110
rect 88470 13836 88570 15026
rect 89560 15026 89566 15318
rect 89600 15026 89606 15318
rect 89560 15014 89606 15026
rect 90618 15318 90664 15330
rect 90618 15026 90624 15318
rect 90658 15026 90664 15318
rect 90618 15014 90664 15026
rect 91676 15318 91722 15330
rect 91676 15026 91682 15318
rect 91716 15026 91722 15318
rect 91676 15014 91722 15026
rect 92734 15318 92780 15330
rect 92734 15026 92740 15318
rect 92774 15026 92780 15318
rect 93792 15318 93838 15330
rect 93792 15176 93798 15318
rect 92734 15014 92780 15026
rect 93764 15026 93798 15176
rect 93832 15176 93838 15318
rect 93832 15026 93864 15176
rect 88470 13658 88508 13836
rect 88502 13544 88508 13658
rect 88542 13658 88570 13836
rect 89560 13836 89606 13848
rect 88542 13544 88548 13658
rect 88502 13532 88548 13544
rect 89560 13544 89566 13836
rect 89600 13544 89606 13836
rect 89560 13532 89606 13544
rect 90618 13836 90664 13848
rect 90618 13544 90624 13836
rect 90658 13544 90664 13836
rect 90618 13532 90664 13544
rect 91676 13836 91722 13848
rect 91676 13544 91682 13836
rect 91716 13544 91722 13836
rect 91676 13532 91722 13544
rect 92734 13836 92780 13848
rect 92734 13544 92740 13836
rect 92774 13544 92780 13836
rect 93764 13836 93864 15026
rect 93764 13724 93798 13836
rect 92734 13532 92780 13544
rect 93792 13544 93798 13724
rect 93832 13724 93864 13836
rect 93832 13544 93838 13724
rect 93792 13532 93838 13544
rect 88502 12742 88548 12754
rect 88502 12450 88508 12742
rect 88542 12450 88548 12742
rect 88502 12438 88548 12450
rect 89560 12742 89606 12754
rect 89560 12450 89566 12742
rect 89600 12450 89606 12742
rect 89560 12438 89606 12450
rect 90618 12742 90664 12754
rect 90618 12450 90624 12742
rect 90658 12450 90664 12742
rect 90618 12438 90664 12450
rect 91676 12742 91722 12754
rect 91676 12450 91682 12742
rect 91716 12450 91722 12742
rect 91676 12438 91722 12450
rect 92734 12742 92780 12754
rect 92734 12450 92740 12742
rect 92774 12450 92780 12742
rect 92734 12438 92780 12450
rect 93792 12742 93838 12754
rect 93792 12450 93798 12742
rect 93832 12450 93838 12742
rect 93792 12438 93838 12450
rect 81736 11654 81782 11666
rect 81736 11362 81742 11654
rect 81776 11362 81782 11654
rect 81736 11350 81782 11362
rect 82794 11654 82840 11666
rect 82794 11362 82800 11654
rect 82834 11362 82840 11654
rect 82794 11350 82840 11362
rect 83852 11654 83898 11666
rect 83852 11362 83858 11654
rect 83892 11362 83898 11654
rect 83852 11350 83898 11362
rect 84910 11654 84956 11666
rect 84910 11362 84916 11654
rect 84950 11362 84956 11654
rect 84910 11350 84956 11362
rect 85968 11654 86014 11666
rect 85968 11362 85974 11654
rect 86008 11362 86014 11654
rect 85968 11350 86014 11362
rect 87026 11654 87072 11666
rect 87026 11362 87032 11654
rect 87066 11362 87072 11654
rect 87026 11350 87072 11362
rect 75268 10562 75314 10574
rect 75268 10270 75274 10562
rect 75308 10270 75314 10562
rect 75268 10258 75314 10270
rect 76326 10562 76372 10574
rect 76326 10270 76332 10562
rect 76366 10270 76372 10562
rect 76326 10258 76372 10270
rect 77384 10562 77430 10574
rect 77384 10270 77390 10562
rect 77424 10270 77430 10562
rect 77384 10258 77430 10270
rect 78442 10562 78488 10574
rect 78442 10270 78448 10562
rect 78482 10270 78488 10562
rect 78442 10258 78488 10270
rect 79500 10562 79546 10574
rect 79500 10270 79506 10562
rect 79540 10270 79546 10562
rect 79500 10258 79546 10270
rect 80558 10562 80604 10574
rect 80558 10270 80564 10562
rect 80598 10270 80604 10562
rect 80558 10258 80604 10270
rect 75268 9468 75314 9480
rect 75268 9264 75274 9468
rect 75248 9176 75274 9264
rect 75308 9264 75314 9468
rect 76326 9468 76372 9480
rect 75308 9176 75348 9264
rect 75248 7986 75348 9176
rect 76326 9176 76332 9468
rect 76366 9176 76372 9468
rect 76326 9164 76372 9176
rect 77384 9468 77430 9480
rect 77384 9176 77390 9468
rect 77424 9176 77430 9468
rect 77384 9164 77430 9176
rect 78442 9468 78488 9480
rect 78442 9176 78448 9468
rect 78482 9176 78488 9468
rect 78442 9164 78488 9176
rect 79500 9468 79546 9480
rect 79500 9176 79506 9468
rect 79540 9176 79546 9468
rect 80558 9468 80604 9480
rect 80558 9298 80564 9468
rect 79500 9164 79546 9176
rect 80518 9176 80564 9298
rect 80598 9298 80604 9468
rect 80598 9176 80618 9298
rect 75248 7812 75274 7986
rect 75268 7694 75274 7812
rect 75308 7812 75348 7986
rect 76326 7986 76372 7998
rect 75308 7694 75314 7812
rect 75268 7682 75314 7694
rect 76326 7694 76332 7986
rect 76366 7694 76372 7986
rect 76326 7682 76372 7694
rect 77384 7986 77430 7998
rect 77384 7694 77390 7986
rect 77424 7694 77430 7986
rect 77384 7682 77430 7694
rect 78442 7986 78488 7998
rect 78442 7694 78448 7986
rect 78482 7694 78488 7986
rect 78442 7682 78488 7694
rect 79500 7986 79546 7998
rect 79500 7694 79506 7986
rect 79540 7694 79546 7986
rect 80518 7986 80618 9176
rect 80518 7846 80564 7986
rect 79500 7682 79546 7694
rect 80558 7694 80564 7846
rect 80598 7846 80618 7986
rect 80598 7694 80604 7846
rect 80558 7682 80604 7694
rect 75268 6892 75314 6904
rect 75268 6600 75274 6892
rect 75308 6600 75314 6892
rect 75268 6588 75314 6600
rect 76326 6892 76372 6904
rect 76326 6600 76332 6892
rect 76366 6600 76372 6892
rect 76326 6588 76372 6600
rect 77384 6892 77430 6904
rect 77384 6600 77390 6892
rect 77424 6600 77430 6892
rect 77384 6588 77430 6600
rect 78442 6892 78488 6904
rect 78442 6600 78448 6892
rect 78482 6600 78488 6892
rect 78442 6588 78488 6600
rect 79500 6892 79546 6904
rect 79500 6600 79506 6892
rect 79540 6600 79546 6892
rect 79500 6588 79546 6600
rect 80558 6892 80604 6904
rect 80558 6600 80564 6892
rect 80598 6600 80604 6892
rect 80558 6588 80604 6600
rect 68584 5824 68630 5836
rect 68052 5282 68086 5592
rect 68584 5532 68590 5824
rect 68624 5532 68630 5824
rect 68584 5520 68630 5532
rect 69642 5824 69688 5836
rect 69642 5532 69648 5824
rect 69682 5532 69688 5824
rect 69642 5520 69688 5532
rect 70700 5824 70746 5836
rect 70700 5532 70706 5824
rect 70740 5532 70746 5824
rect 70700 5520 70746 5532
rect 71758 5824 71804 5836
rect 71758 5532 71764 5824
rect 71798 5532 71804 5824
rect 71758 5520 71804 5532
rect 72816 5824 72862 5836
rect 72816 5532 72822 5824
rect 72856 5532 72862 5824
rect 72816 5520 72862 5532
rect 73874 5824 73920 5836
rect 73874 5532 73880 5824
rect 73914 5532 73920 5824
rect 73874 5520 73920 5532
rect 74374 5408 74642 6452
rect 67936 4958 68086 5282
rect 74620 5256 74642 5408
rect 74736 5408 74964 6452
rect 80820 6450 81372 11112
rect 87672 11106 87876 12302
rect 87970 11106 88224 12302
rect 94120 12300 94672 16976
rect 94966 16424 95012 16436
rect 94966 16132 94972 16424
rect 95006 16132 95012 16424
rect 94966 16120 95012 16132
rect 96024 16424 96070 16436
rect 96024 16132 96030 16424
rect 96064 16132 96070 16424
rect 96024 16120 96070 16132
rect 97082 16424 97128 16436
rect 97082 16132 97088 16424
rect 97122 16132 97128 16424
rect 97082 16120 97128 16132
rect 98140 16424 98186 16436
rect 98140 16132 98146 16424
rect 98180 16132 98186 16424
rect 98140 16120 98186 16132
rect 99198 16424 99244 16436
rect 99198 16132 99204 16424
rect 99238 16132 99244 16424
rect 99198 16120 99244 16132
rect 100256 16424 100302 16436
rect 100256 16132 100262 16424
rect 100296 16132 100302 16424
rect 100256 16120 100302 16132
rect 100630 15392 100742 18976
rect 101120 15392 101376 18976
rect 94966 15330 95012 15342
rect 94966 15144 94972 15330
rect 94908 15038 94972 15144
rect 95006 15038 95012 15330
rect 94908 15026 95012 15038
rect 96024 15330 96070 15342
rect 96024 15038 96030 15330
rect 96064 15038 96070 15330
rect 96024 15026 96070 15038
rect 97082 15330 97128 15342
rect 97082 15038 97088 15330
rect 97122 15038 97128 15330
rect 97082 15026 97128 15038
rect 98140 15330 98186 15342
rect 98140 15038 98146 15330
rect 98180 15038 98186 15330
rect 98140 15026 98186 15038
rect 99198 15330 99244 15342
rect 99198 15038 99204 15330
rect 99238 15038 99244 15330
rect 100256 15330 100302 15342
rect 100256 15144 100262 15330
rect 99198 15026 99244 15038
rect 100190 15038 100262 15144
rect 100296 15144 100302 15330
rect 100296 15038 100322 15144
rect 94908 13846 95008 15026
rect 94908 13834 95016 13846
rect 94908 13692 94976 13834
rect 94970 13542 94976 13692
rect 95010 13542 95016 13834
rect 94970 13530 95016 13542
rect 96028 13834 96074 13846
rect 96028 13542 96034 13834
rect 96068 13542 96074 13834
rect 96028 13530 96074 13542
rect 97086 13834 97132 13846
rect 97086 13542 97092 13834
rect 97126 13542 97132 13834
rect 97086 13530 97132 13542
rect 98144 13834 98190 13846
rect 98144 13542 98150 13834
rect 98184 13542 98190 13834
rect 98144 13530 98190 13542
rect 99202 13834 99248 13846
rect 99202 13542 99208 13834
rect 99242 13542 99248 13834
rect 100190 13834 100322 15038
rect 100630 14880 101376 15392
rect 100788 13902 101376 14880
rect 100190 13648 100266 13834
rect 99202 13530 99248 13542
rect 100260 13542 100266 13648
rect 100300 13648 100322 13834
rect 100300 13542 100306 13648
rect 100260 13530 100306 13542
rect 100630 13456 101376 13902
rect 94970 12740 95016 12752
rect 94970 12448 94976 12740
rect 95010 12448 95016 12740
rect 94970 12436 95016 12448
rect 96028 12740 96074 12752
rect 96028 12448 96034 12740
rect 96068 12448 96074 12740
rect 96028 12436 96074 12448
rect 97086 12740 97132 12752
rect 97086 12448 97092 12740
rect 97126 12448 97132 12740
rect 97086 12436 97132 12448
rect 98144 12740 98190 12752
rect 98144 12448 98150 12740
rect 98184 12448 98190 12740
rect 98144 12436 98190 12448
rect 99202 12740 99248 12752
rect 99202 12448 99208 12740
rect 99242 12448 99248 12740
rect 99202 12436 99248 12448
rect 100260 12740 100306 12752
rect 100260 12448 100266 12740
rect 100300 12448 100306 12740
rect 100260 12436 100306 12448
rect 88502 11648 88548 11660
rect 88502 11356 88508 11648
rect 88542 11356 88548 11648
rect 88502 11344 88548 11356
rect 89560 11648 89606 11660
rect 89560 11356 89566 11648
rect 89600 11356 89606 11648
rect 89560 11344 89606 11356
rect 90618 11648 90664 11660
rect 90618 11356 90624 11648
rect 90658 11356 90664 11648
rect 90618 11344 90664 11356
rect 91676 11648 91722 11660
rect 91676 11356 91682 11648
rect 91716 11356 91722 11648
rect 91676 11344 91722 11356
rect 92734 11648 92780 11660
rect 92734 11356 92740 11648
rect 92774 11356 92780 11648
rect 92734 11344 92780 11356
rect 93792 11648 93838 11660
rect 93792 11356 93798 11648
rect 93832 11356 93838 11648
rect 93792 11344 93838 11356
rect 81736 10560 81782 10572
rect 81736 10268 81742 10560
rect 81776 10268 81782 10560
rect 81736 10256 81782 10268
rect 82794 10560 82840 10572
rect 82794 10268 82800 10560
rect 82834 10268 82840 10560
rect 82794 10256 82840 10268
rect 83852 10560 83898 10572
rect 83852 10268 83858 10560
rect 83892 10268 83898 10560
rect 83852 10256 83898 10268
rect 84910 10560 84956 10572
rect 84910 10268 84916 10560
rect 84950 10268 84956 10560
rect 84910 10256 84956 10268
rect 85968 10560 86014 10572
rect 85968 10268 85974 10560
rect 86008 10268 86014 10560
rect 85968 10256 86014 10268
rect 87026 10560 87072 10572
rect 87026 10268 87032 10560
rect 87066 10268 87072 10560
rect 87026 10256 87072 10268
rect 81736 9466 81782 9478
rect 81736 9320 81742 9466
rect 81706 9174 81742 9320
rect 81776 9320 81782 9466
rect 82794 9466 82840 9478
rect 81776 9174 81806 9320
rect 81706 7984 81806 9174
rect 82794 9174 82800 9466
rect 82834 9174 82840 9466
rect 82794 9162 82840 9174
rect 83852 9466 83898 9478
rect 83852 9174 83858 9466
rect 83892 9174 83898 9466
rect 83852 9162 83898 9174
rect 84910 9466 84956 9478
rect 84910 9174 84916 9466
rect 84950 9174 84956 9466
rect 84910 9162 84956 9174
rect 85968 9466 86014 9478
rect 85968 9174 85974 9466
rect 86008 9174 86014 9466
rect 87026 9466 87072 9478
rect 87026 9396 87032 9466
rect 85968 9162 86014 9174
rect 86988 9174 87032 9396
rect 87066 9396 87072 9466
rect 87066 9174 87120 9396
rect 81706 7868 81746 7984
rect 81740 7692 81746 7868
rect 81780 7868 81806 7984
rect 82798 7984 82844 7996
rect 81780 7692 81786 7868
rect 81740 7680 81786 7692
rect 82798 7692 82804 7984
rect 82838 7692 82844 7984
rect 82798 7680 82844 7692
rect 83856 7984 83902 7996
rect 83856 7692 83862 7984
rect 83896 7692 83902 7984
rect 83856 7680 83902 7692
rect 84914 7984 84960 7996
rect 84914 7692 84920 7984
rect 84954 7692 84960 7984
rect 84914 7680 84960 7692
rect 85972 7984 86018 7996
rect 85972 7692 85978 7984
rect 86012 7692 86018 7984
rect 86988 7984 87120 9174
rect 86988 7900 87036 7984
rect 85972 7680 86018 7692
rect 87030 7692 87036 7900
rect 87070 7900 87120 7984
rect 87070 7692 87076 7900
rect 87030 7680 87076 7692
rect 81740 6890 81786 6902
rect 81740 6598 81746 6890
rect 81780 6598 81786 6890
rect 81740 6586 81786 6598
rect 82798 6890 82844 6902
rect 82798 6598 82804 6890
rect 82838 6598 82844 6890
rect 82798 6586 82844 6598
rect 83856 6890 83902 6902
rect 83856 6598 83862 6890
rect 83896 6598 83902 6890
rect 83856 6586 83902 6598
rect 84914 6890 84960 6902
rect 84914 6598 84920 6890
rect 84954 6598 84960 6890
rect 84914 6586 84960 6598
rect 85972 6890 86018 6902
rect 85972 6598 85978 6890
rect 86012 6598 86018 6890
rect 85972 6586 86018 6598
rect 87030 6890 87076 6902
rect 87030 6598 87036 6890
rect 87070 6598 87076 6890
rect 87030 6586 87076 6598
rect 75268 5798 75314 5810
rect 75268 5506 75274 5798
rect 75308 5506 75314 5798
rect 75268 5494 75314 5506
rect 76326 5798 76372 5810
rect 76326 5506 76332 5798
rect 76366 5506 76372 5798
rect 76326 5494 76372 5506
rect 77384 5798 77430 5810
rect 77384 5506 77390 5798
rect 77424 5506 77430 5798
rect 77384 5494 77430 5506
rect 78442 5798 78488 5810
rect 78442 5506 78448 5798
rect 78482 5506 78488 5798
rect 78442 5494 78488 5506
rect 79500 5798 79546 5810
rect 79500 5506 79506 5798
rect 79540 5506 79546 5798
rect 79500 5494 79546 5506
rect 80558 5798 80604 5810
rect 80558 5506 80564 5798
rect 80598 5506 80604 5798
rect 80558 5494 80604 5506
rect 74736 5256 74770 5408
rect 74620 4932 74770 5256
rect 80820 5254 81114 6450
rect 81208 5254 81372 6450
rect 87672 6444 88224 11106
rect 94120 11104 94344 12300
rect 94438 11104 94672 12300
rect 94970 11646 95016 11658
rect 94970 11354 94976 11646
rect 95010 11354 95016 11646
rect 94970 11342 95016 11354
rect 96028 11646 96074 11658
rect 96028 11354 96034 11646
rect 96068 11354 96074 11646
rect 96028 11342 96074 11354
rect 97086 11646 97132 11658
rect 97086 11354 97092 11646
rect 97126 11354 97132 11646
rect 97086 11342 97132 11354
rect 98144 11646 98190 11658
rect 98144 11354 98150 11646
rect 98184 11354 98190 11646
rect 98144 11342 98190 11354
rect 99202 11646 99248 11658
rect 99202 11354 99208 11646
rect 99242 11354 99248 11646
rect 99202 11342 99248 11354
rect 100260 11646 100306 11658
rect 100260 11354 100266 11646
rect 100300 11354 100306 11646
rect 100260 11342 100306 11354
rect 88502 10554 88548 10566
rect 88502 10262 88508 10554
rect 88542 10262 88548 10554
rect 88502 10250 88548 10262
rect 89560 10554 89606 10566
rect 89560 10262 89566 10554
rect 89600 10262 89606 10554
rect 89560 10250 89606 10262
rect 90618 10554 90664 10566
rect 90618 10262 90624 10554
rect 90658 10262 90664 10554
rect 90618 10250 90664 10262
rect 91676 10554 91722 10566
rect 91676 10262 91682 10554
rect 91716 10262 91722 10554
rect 91676 10250 91722 10262
rect 92734 10554 92780 10566
rect 92734 10262 92740 10554
rect 92774 10262 92780 10554
rect 92734 10250 92780 10262
rect 93792 10554 93838 10566
rect 93792 10262 93798 10554
rect 93832 10262 93838 10554
rect 93792 10250 93838 10262
rect 88502 9460 88548 9472
rect 88502 9256 88508 9460
rect 88482 9168 88508 9256
rect 88542 9256 88548 9460
rect 89560 9460 89606 9472
rect 88542 9168 88582 9256
rect 88482 7978 88582 9168
rect 89560 9168 89566 9460
rect 89600 9168 89606 9460
rect 89560 9156 89606 9168
rect 90618 9460 90664 9472
rect 90618 9168 90624 9460
rect 90658 9168 90664 9460
rect 90618 9156 90664 9168
rect 91676 9460 91722 9472
rect 91676 9168 91682 9460
rect 91716 9168 91722 9460
rect 91676 9156 91722 9168
rect 92734 9460 92780 9472
rect 92734 9168 92740 9460
rect 92774 9168 92780 9460
rect 93792 9460 93838 9472
rect 93792 9290 93798 9460
rect 92734 9156 92780 9168
rect 93752 9168 93798 9290
rect 93832 9290 93838 9460
rect 93832 9168 93852 9290
rect 88482 7804 88508 7978
rect 88502 7686 88508 7804
rect 88542 7804 88582 7978
rect 89560 7978 89606 7990
rect 88542 7686 88548 7804
rect 88502 7674 88548 7686
rect 89560 7686 89566 7978
rect 89600 7686 89606 7978
rect 89560 7674 89606 7686
rect 90618 7978 90664 7990
rect 90618 7686 90624 7978
rect 90658 7686 90664 7978
rect 90618 7674 90664 7686
rect 91676 7978 91722 7990
rect 91676 7686 91682 7978
rect 91716 7686 91722 7978
rect 91676 7674 91722 7686
rect 92734 7978 92780 7990
rect 92734 7686 92740 7978
rect 92774 7686 92780 7978
rect 93752 7978 93852 9168
rect 93752 7838 93798 7978
rect 92734 7674 92780 7686
rect 93792 7686 93798 7838
rect 93832 7838 93852 7978
rect 93832 7686 93838 7838
rect 93792 7674 93838 7686
rect 88502 6884 88548 6896
rect 88502 6592 88508 6884
rect 88542 6592 88548 6884
rect 88502 6580 88548 6592
rect 89560 6884 89606 6896
rect 89560 6592 89566 6884
rect 89600 6592 89606 6884
rect 89560 6580 89606 6592
rect 90618 6884 90664 6896
rect 90618 6592 90624 6884
rect 90658 6592 90664 6884
rect 90618 6580 90664 6592
rect 91676 6884 91722 6896
rect 91676 6592 91682 6884
rect 91716 6592 91722 6884
rect 91676 6580 91722 6592
rect 92734 6884 92780 6896
rect 92734 6592 92740 6884
rect 92774 6592 92780 6884
rect 92734 6580 92780 6592
rect 93792 6884 93838 6896
rect 93792 6592 93798 6884
rect 93832 6592 93838 6884
rect 93792 6580 93838 6592
rect 81740 5796 81786 5808
rect 81740 5504 81746 5796
rect 81780 5504 81786 5796
rect 81740 5492 81786 5504
rect 82798 5796 82844 5808
rect 82798 5504 82804 5796
rect 82838 5504 82844 5796
rect 82798 5492 82844 5504
rect 83856 5796 83902 5808
rect 83856 5504 83862 5796
rect 83896 5504 83902 5796
rect 83856 5492 83902 5504
rect 84914 5796 84960 5808
rect 84914 5504 84920 5796
rect 84954 5504 84960 5796
rect 84914 5492 84960 5504
rect 85972 5796 86018 5808
rect 85972 5504 85978 5796
rect 86012 5504 86018 5796
rect 85972 5492 86018 5504
rect 87030 5796 87076 5808
rect 87030 5504 87036 5796
rect 87070 5504 87076 5796
rect 87030 5492 87076 5504
rect 62112 4732 62158 4744
rect 62112 4440 62118 4732
rect 62152 4440 62158 4732
rect 62112 4428 62158 4440
rect 63170 4732 63216 4744
rect 63170 4440 63176 4732
rect 63210 4440 63216 4732
rect 63170 4428 63216 4440
rect 64228 4732 64274 4744
rect 64228 4440 64234 4732
rect 64268 4440 64274 4732
rect 64228 4428 64274 4440
rect 65286 4732 65332 4744
rect 65286 4440 65292 4732
rect 65326 4440 65332 4732
rect 65286 4428 65332 4440
rect 66344 4732 66390 4744
rect 66344 4440 66350 4732
rect 66384 4440 66390 4732
rect 66344 4428 66390 4440
rect 67402 4732 67448 4744
rect 67402 4440 67408 4732
rect 67442 4440 67448 4732
rect 67402 4428 67448 4440
rect 68584 4730 68630 4742
rect 68584 4438 68590 4730
rect 68624 4438 68630 4730
rect 68584 4426 68630 4438
rect 69642 4730 69688 4742
rect 69642 4438 69648 4730
rect 69682 4438 69688 4730
rect 69642 4426 69688 4438
rect 70700 4730 70746 4742
rect 70700 4438 70706 4730
rect 70740 4438 70746 4730
rect 70700 4426 70746 4438
rect 71758 4730 71804 4742
rect 71758 4438 71764 4730
rect 71798 4438 71804 4730
rect 71758 4426 71804 4438
rect 72816 4730 72862 4742
rect 72816 4438 72822 4730
rect 72856 4438 72862 4730
rect 72816 4426 72862 4438
rect 73874 4730 73920 4742
rect 73874 4438 73880 4730
rect 73914 4438 73920 4730
rect 73874 4426 73920 4438
rect 75268 4704 75314 4716
rect 75268 4412 75274 4704
rect 75308 4412 75314 4704
rect 75268 4400 75314 4412
rect 76326 4704 76372 4716
rect 76326 4412 76332 4704
rect 76366 4412 76372 4704
rect 76326 4400 76372 4412
rect 77384 4704 77430 4716
rect 77384 4412 77390 4704
rect 77424 4412 77430 4704
rect 77384 4400 77430 4412
rect 78442 4704 78488 4716
rect 78442 4412 78448 4704
rect 78482 4412 78488 4704
rect 78442 4400 78488 4412
rect 79500 4704 79546 4716
rect 79500 4412 79506 4704
rect 79540 4412 79546 4704
rect 79500 4400 79546 4412
rect 80558 4704 80604 4716
rect 80558 4412 80564 4704
rect 80598 4412 80604 4704
rect 80558 4400 80604 4412
rect 62112 3638 62158 3650
rect 62112 3346 62118 3638
rect 62152 3346 62158 3638
rect 62112 3334 62158 3346
rect 63170 3638 63216 3650
rect 63170 3346 63176 3638
rect 63210 3346 63216 3638
rect 63170 3334 63216 3346
rect 64228 3638 64274 3650
rect 64228 3346 64234 3638
rect 64268 3346 64274 3638
rect 64228 3334 64274 3346
rect 65286 3638 65332 3650
rect 65286 3346 65292 3638
rect 65326 3346 65332 3638
rect 65286 3334 65332 3346
rect 66344 3638 66390 3650
rect 66344 3346 66350 3638
rect 66384 3346 66390 3638
rect 66344 3334 66390 3346
rect 67402 3638 67448 3650
rect 67402 3346 67408 3638
rect 67442 3346 67448 3638
rect 67402 3334 67448 3346
rect 68584 3636 68630 3648
rect 68584 3344 68590 3636
rect 68624 3344 68630 3636
rect 68584 3332 68630 3344
rect 69642 3636 69688 3648
rect 69642 3344 69648 3636
rect 69682 3344 69688 3636
rect 69642 3332 69688 3344
rect 70700 3636 70746 3648
rect 70700 3344 70706 3636
rect 70740 3344 70746 3636
rect 70700 3332 70746 3344
rect 71758 3636 71804 3648
rect 71758 3344 71764 3636
rect 71798 3344 71804 3636
rect 71758 3332 71804 3344
rect 72816 3636 72862 3648
rect 72816 3344 72822 3636
rect 72856 3344 72862 3636
rect 72816 3332 72862 3344
rect 73874 3636 73920 3648
rect 73874 3344 73880 3636
rect 73914 3344 73920 3636
rect 75268 3610 75314 3622
rect 75268 3416 75274 3610
rect 73874 3332 73920 3344
rect 59404 3316 59450 3328
rect 75142 3318 75274 3416
rect 75308 3416 75314 3610
rect 76326 3610 76372 3622
rect 75308 3318 75380 3416
rect 52890 3302 52936 3314
rect 46302 3280 46348 3292
rect 75142 2594 75380 3318
rect 76326 3318 76332 3610
rect 76366 3318 76372 3610
rect 76326 3306 76372 3318
rect 77384 3610 77430 3622
rect 77384 3318 77390 3610
rect 77424 3318 77430 3610
rect 77384 3306 77430 3318
rect 78442 3610 78488 3622
rect 78442 3318 78448 3610
rect 78482 3318 78488 3610
rect 78442 3306 78488 3318
rect 79500 3610 79546 3622
rect 79500 3318 79506 3610
rect 79540 3318 79546 3610
rect 79500 3306 79546 3318
rect 80558 3610 80604 3622
rect 80558 3318 80564 3610
rect 80598 3318 80604 3610
rect 80558 3306 80604 3318
rect 39688 2392 75380 2594
rect 75142 2284 75380 2392
rect 67068 840 69266 846
rect 59508 -184 60606 -178
rect 39824 -496 41570 -490
rect 39824 -1246 39836 -496
rect 41558 -1246 41570 -496
rect 59508 -682 59520 -184
rect 60594 -682 60606 -184
rect 67068 -192 67080 840
rect 69254 -192 69266 840
rect 67068 -198 69266 -192
rect 73662 804 75860 810
rect 59508 -688 60606 -682
rect 39824 -1252 41570 -1246
rect 40284 -3192 40658 -1252
rect 59810 -3192 60142 -688
rect 67632 -3192 68480 -198
rect 73662 -228 73674 804
rect 75848 -228 75860 804
rect 73662 -234 75860 -228
rect 74154 -3192 75258 -234
rect 80820 -3192 81372 5254
rect 87672 5248 87876 6444
rect 87970 5248 88224 6444
rect 94120 6442 94672 11104
rect 94970 10552 95016 10564
rect 94970 10260 94976 10552
rect 95010 10260 95016 10552
rect 94970 10248 95016 10260
rect 96028 10552 96074 10564
rect 96028 10260 96034 10552
rect 96068 10260 96074 10552
rect 96028 10248 96074 10260
rect 97086 10552 97132 10564
rect 97086 10260 97092 10552
rect 97126 10260 97132 10552
rect 97086 10248 97132 10260
rect 98144 10552 98190 10564
rect 98144 10260 98150 10552
rect 98184 10260 98190 10552
rect 98144 10248 98190 10260
rect 99202 10552 99248 10564
rect 99202 10260 99208 10552
rect 99242 10260 99248 10552
rect 99202 10248 99248 10260
rect 100260 10552 100306 10564
rect 100260 10260 100266 10552
rect 100300 10260 100306 10552
rect 100260 10248 100306 10260
rect 100630 9760 100876 13456
rect 101098 9760 101376 13456
rect 94970 9458 95016 9470
rect 94970 9312 94976 9458
rect 94940 9166 94976 9312
rect 95010 9312 95016 9458
rect 96028 9458 96074 9470
rect 95010 9166 95040 9312
rect 94940 7976 95040 9166
rect 96028 9166 96034 9458
rect 96068 9166 96074 9458
rect 96028 9154 96074 9166
rect 97086 9458 97132 9470
rect 97086 9166 97092 9458
rect 97126 9166 97132 9458
rect 97086 9154 97132 9166
rect 98144 9458 98190 9470
rect 98144 9166 98150 9458
rect 98184 9166 98190 9458
rect 98144 9154 98190 9166
rect 99202 9458 99248 9470
rect 99202 9166 99208 9458
rect 99242 9166 99248 9458
rect 100260 9458 100306 9470
rect 100260 9388 100266 9458
rect 99202 9154 99248 9166
rect 100222 9166 100266 9388
rect 100300 9388 100306 9458
rect 100300 9166 100354 9388
rect 100630 9294 101376 9760
rect 94940 7860 94980 7976
rect 94974 7684 94980 7860
rect 95014 7860 95040 7976
rect 96032 7976 96078 7988
rect 95014 7684 95020 7860
rect 94974 7672 95020 7684
rect 96032 7684 96038 7976
rect 96072 7684 96078 7976
rect 96032 7672 96078 7684
rect 97090 7976 97136 7988
rect 97090 7684 97096 7976
rect 97130 7684 97136 7976
rect 97090 7672 97136 7684
rect 98148 7976 98194 7988
rect 98148 7684 98154 7976
rect 98188 7684 98194 7976
rect 98148 7672 98194 7684
rect 99206 7976 99252 7988
rect 99206 7684 99212 7976
rect 99246 7684 99252 7976
rect 100222 7976 100354 9166
rect 100222 7892 100270 7976
rect 99206 7672 99252 7684
rect 100264 7684 100270 7892
rect 100304 7892 100354 7976
rect 100304 7684 100310 7892
rect 100788 7712 101376 9294
rect 100264 7672 100310 7684
rect 100608 7268 101376 7712
rect 94974 6882 95020 6894
rect 94974 6590 94980 6882
rect 95014 6590 95020 6882
rect 94974 6578 95020 6590
rect 96032 6882 96078 6894
rect 96032 6590 96038 6882
rect 96072 6590 96078 6882
rect 96032 6578 96078 6590
rect 97090 6882 97136 6894
rect 97090 6590 97096 6882
rect 97130 6590 97136 6882
rect 97090 6578 97136 6590
rect 98148 6882 98194 6894
rect 98148 6590 98154 6882
rect 98188 6590 98194 6882
rect 98148 6578 98194 6590
rect 99206 6882 99252 6894
rect 99206 6590 99212 6882
rect 99246 6590 99252 6882
rect 99206 6578 99252 6590
rect 100264 6882 100310 6894
rect 100264 6590 100270 6882
rect 100304 6590 100310 6882
rect 100264 6578 100310 6590
rect 88502 5790 88548 5802
rect 88502 5498 88508 5790
rect 88542 5498 88548 5790
rect 88502 5486 88548 5498
rect 89560 5790 89606 5802
rect 89560 5498 89566 5790
rect 89600 5498 89606 5790
rect 89560 5486 89606 5498
rect 90618 5790 90664 5802
rect 90618 5498 90624 5790
rect 90658 5498 90664 5790
rect 90618 5486 90664 5498
rect 91676 5790 91722 5802
rect 91676 5498 91682 5790
rect 91716 5498 91722 5790
rect 91676 5486 91722 5498
rect 92734 5790 92780 5802
rect 92734 5498 92740 5790
rect 92774 5498 92780 5790
rect 92734 5486 92780 5498
rect 93792 5790 93838 5802
rect 93792 5498 93798 5790
rect 93832 5498 93838 5790
rect 93792 5486 93838 5498
rect 81740 4702 81786 4714
rect 81740 4410 81746 4702
rect 81780 4410 81786 4702
rect 81740 4398 81786 4410
rect 82798 4702 82844 4714
rect 82798 4410 82804 4702
rect 82838 4410 82844 4702
rect 82798 4398 82844 4410
rect 83856 4702 83902 4714
rect 83856 4410 83862 4702
rect 83896 4410 83902 4702
rect 83856 4398 83902 4410
rect 84914 4702 84960 4714
rect 84914 4410 84920 4702
rect 84954 4410 84960 4702
rect 84914 4398 84960 4410
rect 85972 4702 86018 4714
rect 85972 4410 85978 4702
rect 86012 4410 86018 4702
rect 85972 4398 86018 4410
rect 87030 4702 87076 4714
rect 87030 4410 87036 4702
rect 87070 4410 87076 4702
rect 87030 4398 87076 4410
rect 81740 3608 81786 3620
rect 81740 3316 81746 3608
rect 81780 3316 81786 3608
rect 81740 3304 81786 3316
rect 82798 3608 82844 3620
rect 82798 3316 82804 3608
rect 82838 3316 82844 3608
rect 82798 3304 82844 3316
rect 83856 3608 83902 3620
rect 83856 3316 83862 3608
rect 83896 3316 83902 3608
rect 83856 3304 83902 3316
rect 84914 3608 84960 3620
rect 84914 3316 84920 3608
rect 84954 3316 84960 3608
rect 84914 3304 84960 3316
rect 85972 3608 86018 3620
rect 85972 3316 85978 3608
rect 86012 3316 86018 3608
rect 87030 3608 87076 3620
rect 87030 3590 87036 3608
rect 87006 3340 87036 3590
rect 85972 3304 86018 3316
rect 87030 3316 87036 3340
rect 87070 3590 87076 3608
rect 87672 3590 88224 5248
rect 94120 5246 94348 6442
rect 94442 5246 94672 6442
rect 94974 5788 95020 5800
rect 94974 5496 94980 5788
rect 95014 5496 95020 5788
rect 94974 5484 95020 5496
rect 96032 5788 96078 5800
rect 96032 5496 96038 5788
rect 96072 5496 96078 5788
rect 96032 5484 96078 5496
rect 97090 5788 97136 5800
rect 97090 5496 97096 5788
rect 97130 5496 97136 5788
rect 97090 5484 97136 5496
rect 98148 5788 98194 5800
rect 98148 5496 98154 5788
rect 98188 5496 98194 5788
rect 98148 5484 98194 5496
rect 99206 5788 99252 5800
rect 99206 5496 99212 5788
rect 99246 5496 99252 5788
rect 99206 5484 99252 5496
rect 100264 5788 100310 5800
rect 100264 5496 100270 5788
rect 100304 5496 100310 5788
rect 100264 5484 100310 5496
rect 88502 4696 88548 4708
rect 88502 4404 88508 4696
rect 88542 4404 88548 4696
rect 88502 4392 88548 4404
rect 89560 4696 89606 4708
rect 89560 4404 89566 4696
rect 89600 4404 89606 4696
rect 89560 4392 89606 4404
rect 90618 4696 90664 4708
rect 90618 4404 90624 4696
rect 90658 4404 90664 4696
rect 90618 4392 90664 4404
rect 91676 4696 91722 4708
rect 91676 4404 91682 4696
rect 91716 4404 91722 4696
rect 91676 4392 91722 4404
rect 92734 4696 92780 4708
rect 92734 4404 92740 4696
rect 92774 4404 92780 4696
rect 92734 4392 92780 4404
rect 93792 4696 93838 4708
rect 93792 4404 93798 4696
rect 93832 4404 93838 4696
rect 93792 4392 93838 4404
rect 87070 3340 88224 3590
rect 87070 3316 87076 3340
rect 87030 3304 87076 3316
rect 87672 -3192 88224 3340
rect 88502 3602 88548 3614
rect 88502 3310 88508 3602
rect 88542 3310 88548 3602
rect 88502 3298 88548 3310
rect 89560 3602 89606 3614
rect 89560 3310 89566 3602
rect 89600 3310 89606 3602
rect 89560 3298 89606 3310
rect 90618 3602 90664 3614
rect 90618 3310 90624 3602
rect 90658 3310 90664 3602
rect 90618 3298 90664 3310
rect 91676 3602 91722 3614
rect 91676 3310 91682 3602
rect 91716 3310 91722 3602
rect 91676 3298 91722 3310
rect 92734 3602 92780 3614
rect 92734 3310 92740 3602
rect 92774 3310 92780 3602
rect 92734 3298 92780 3310
rect 93792 3602 93838 3614
rect 93792 3310 93798 3602
rect 93832 3310 93838 3602
rect 93792 3298 93838 3310
rect 94120 -3192 94672 5246
rect 94974 4694 95020 4706
rect 94974 4402 94980 4694
rect 95014 4402 95020 4694
rect 94974 4390 95020 4402
rect 96032 4694 96078 4706
rect 96032 4402 96038 4694
rect 96072 4402 96078 4694
rect 96032 4390 96078 4402
rect 97090 4694 97136 4706
rect 97090 4402 97096 4694
rect 97130 4402 97136 4694
rect 97090 4390 97136 4402
rect 98148 4694 98194 4706
rect 98148 4402 98154 4694
rect 98188 4402 98194 4694
rect 98148 4390 98194 4402
rect 99206 4694 99252 4706
rect 99206 4402 99212 4694
rect 99246 4402 99252 4694
rect 99206 4390 99252 4402
rect 100264 4694 100310 4706
rect 100264 4402 100270 4694
rect 100304 4402 100310 4694
rect 100264 4390 100310 4402
rect 94974 3600 95020 3612
rect 94974 3308 94980 3600
rect 95014 3308 95020 3600
rect 94974 3296 95020 3308
rect 96032 3600 96078 3612
rect 96032 3308 96038 3600
rect 96072 3308 96078 3600
rect 96032 3296 96078 3308
rect 97090 3600 97136 3612
rect 97090 3308 97096 3600
rect 97130 3308 97136 3600
rect 97090 3296 97136 3308
rect 98148 3600 98194 3612
rect 98148 3308 98154 3600
rect 98188 3308 98194 3600
rect 98148 3296 98194 3308
rect 99206 3600 99252 3612
rect 99206 3308 99212 3600
rect 99246 3308 99252 3600
rect 99206 3296 99252 3308
rect 100264 3600 100310 3612
rect 100264 3308 100270 3600
rect 100304 3308 100310 3600
rect 100264 3296 100310 3308
rect 100608 3594 100898 7268
rect 101098 3594 101376 7268
rect 100608 3172 101376 3594
rect 100788 -3192 101376 3172
rect 101856 -3192 111286 -3176
rect -588 -9218 111286 -3192
rect 101856 -9328 111286 -9218
<< via1 >>
rect 38848 65126 39974 65882
rect 59236 56850 59510 57262
rect 30980 55430 31268 55738
rect 82976 53912 83164 54070
rect 82558 53468 82674 53658
rect 83008 53424 83100 53498
rect 88276 51730 88474 51918
rect 38424 47838 39756 48764
rect 66824 45974 67244 46688
rect 68198 47424 68884 47812
rect 75724 47308 76368 47790
rect 73060 46020 73674 46882
rect 79170 43104 79870 43578
rect 88552 42666 89804 43684
<< metal2 >>
rect 38848 67730 39922 67740
rect 38848 66930 39922 66940
rect 39152 65892 39538 66930
rect 38848 65882 39974 65892
rect 38848 65116 39974 65126
rect 60520 57272 60932 57282
rect 59236 57262 59510 57272
rect 59510 56956 60520 57174
rect 59236 56840 59510 56850
rect 60520 56770 60932 56780
rect 31454 55766 31654 55776
rect 30980 55738 31268 55748
rect 31268 55524 31454 55630
rect 30980 55420 31268 55430
rect 31454 55398 31654 55408
rect 82976 54070 83164 54080
rect 82976 53902 83164 53912
rect 82558 53658 82674 53668
rect 82674 53468 82680 53654
rect 83018 53508 83086 53902
rect 82558 53458 82680 53468
rect 82568 51232 82680 53458
rect 83008 53498 83100 53508
rect 83008 53414 83100 53424
rect 89286 51966 89526 51976
rect 88276 51918 88474 51928
rect 88474 51860 89118 51864
rect 88474 51794 89286 51860
rect 89034 51790 89286 51794
rect 88276 51720 88474 51730
rect 89526 51790 89544 51860
rect 89286 51720 89526 51730
rect 82500 51222 82792 51232
rect 82500 50964 82792 50974
rect 38454 50414 39552 50424
rect 38454 49652 39552 49662
rect 68170 50012 68902 50022
rect 38540 48774 39118 49652
rect 68170 49466 68902 49476
rect 38424 48764 39756 48774
rect 38424 47828 39756 47838
rect 68312 47822 68620 49466
rect 68198 47812 68884 47822
rect 68198 47414 68884 47424
rect 75724 47790 76368 47800
rect 75724 47298 76368 47308
rect 73060 46882 73674 46892
rect 66824 46688 67244 46698
rect 67244 46212 73060 46578
rect 73060 46010 73674 46020
rect 66824 45964 67244 45974
rect 75884 45904 76188 47298
rect 77922 45994 78764 46004
rect 75856 45858 76958 45904
rect 75828 45650 77922 45858
rect 75856 45560 77922 45650
rect 75856 45180 76182 45560
rect 76398 45544 77922 45560
rect 77922 45280 78764 45290
rect 88708 45818 89786 45828
rect 88708 45240 89786 45250
rect 75856 45076 76228 45180
rect 75856 45054 76188 45076
rect 75866 43464 76188 45054
rect 88982 43694 89414 45240
rect 88552 43684 89804 43694
rect 79170 43578 79870 43588
rect 75866 43200 79170 43464
rect 75866 43190 76188 43200
rect 79170 43100 79870 43104
rect 79170 43094 79608 43100
rect 79798 43094 79870 43100
rect 88552 42656 89804 42666
<< via2 >>
rect 38848 66940 39922 67730
rect 60520 56780 60932 57272
rect 31454 55408 31654 55766
rect 89286 51730 89526 51966
rect 82500 50974 82792 51222
rect 38454 49662 39552 50414
rect 68170 49476 68902 50012
rect 77922 45290 78764 45994
rect 88708 45250 89786 45818
<< metal3 >>
rect 33014 64584 38214 68598
rect 39024 68250 39034 69308
rect 39622 68250 39632 69308
rect 39184 67735 39488 68250
rect 38838 67730 39932 67735
rect 38838 66940 38848 67730
rect 39922 66940 39932 67730
rect 38838 66935 39932 66940
rect 33014 64410 38884 64584
rect 33014 64384 33042 64410
rect 33004 64346 33042 64384
rect 38186 64346 38884 64410
rect 33004 64248 38884 64346
rect 33014 64180 38884 64248
rect 33014 60264 38214 64180
rect 38508 60264 38884 64180
rect 33014 60118 38884 60264
rect 33014 60092 33042 60118
rect 33004 60054 33042 60092
rect 38186 60054 38884 60118
rect 33004 59956 38884 60054
rect 33014 59860 38884 59956
rect 33014 55970 38214 59860
rect 38508 55970 38884 59860
rect 62432 59874 67632 63980
rect 62432 59792 68654 59874
rect 62432 59728 62460 59792
rect 67604 59728 68654 59792
rect 62432 59568 68654 59728
rect 60510 57272 60942 57277
rect 60510 56780 60520 57272
rect 60932 57148 60942 57272
rect 61028 57148 61038 57236
rect 60932 56928 61038 57148
rect 60932 56780 60942 56928
rect 61028 56780 61038 56928
rect 61372 56780 61382 57236
rect 60510 56775 60942 56780
rect 33014 55826 38884 55970
rect 33014 55800 33042 55826
rect 31444 55766 31664 55771
rect 31444 55408 31454 55766
rect 31654 55644 31664 55766
rect 31760 55644 31770 55766
rect 31654 55508 31770 55644
rect 31654 55408 31664 55508
rect 31444 55403 31664 55408
rect 31760 55386 31770 55508
rect 32028 55386 32038 55766
rect 33002 55762 33042 55800
rect 38186 55762 38884 55826
rect 33002 55664 38884 55762
rect 33014 55566 38884 55664
rect 33014 51696 38214 55566
rect 38508 51802 38884 55566
rect 62432 55574 67632 59568
rect 68138 55574 68654 59568
rect 62432 55500 68654 55574
rect 62432 55476 62460 55500
rect 62430 55436 62460 55476
rect 67604 55436 68654 55500
rect 62430 55334 68654 55436
rect 62432 55270 68654 55334
rect 62432 55268 68550 55270
rect 38508 51696 38946 51802
rect 33014 51534 38946 51696
rect 33014 51508 33042 51534
rect 33012 51470 33042 51508
rect 38186 51470 38946 51534
rect 33012 51372 38946 51470
rect 33014 51292 38946 51372
rect 33014 47242 38214 51292
rect 38508 51274 38946 51292
rect 38598 50419 38946 51274
rect 62432 51208 67632 55268
rect 62432 51144 62460 51208
rect 67604 51144 67632 51208
rect 62432 51124 67632 51144
rect 68320 53232 68550 55268
rect 38444 50414 39562 50419
rect 38444 49662 38454 50414
rect 39552 49662 39562 50414
rect 68320 50017 68576 53232
rect 89276 51966 89536 51971
rect 82490 51222 82802 51227
rect 82490 50974 82500 51222
rect 82792 50974 82802 51222
rect 82490 50969 82802 50974
rect 82562 50666 82690 50969
rect 82428 50454 82438 50666
rect 82798 50454 82808 50666
rect 38444 49657 39562 49662
rect 68160 50012 68912 50017
rect 68160 49476 68170 50012
rect 68902 49476 68912 50012
rect 68160 49471 68912 49476
rect 83036 47658 88236 51752
rect 89276 51730 89286 51966
rect 89526 51730 89536 51966
rect 89276 51725 89536 51730
rect 89340 51408 89478 51725
rect 89350 47658 89462 51408
rect 83032 47638 88248 47658
rect 88904 47638 89472 47658
rect 83032 47564 89472 47638
rect 83032 47500 83064 47564
rect 88208 47500 89472 47564
rect 83032 47384 89472 47500
rect 83032 47346 88248 47384
rect 33014 47178 33042 47242
rect 38186 47178 38214 47242
rect 33014 47158 38214 47178
rect 77912 45994 78774 45999
rect 77912 45290 77922 45994
rect 78764 45818 78774 45994
rect 81260 45818 81270 46190
rect 78764 45408 81270 45818
rect 78764 45290 78774 45408
rect 77912 45285 78774 45290
rect 81260 45270 81270 45408
rect 81936 45270 81946 46190
rect 83036 43272 88236 47346
rect 88904 45823 89472 47384
rect 88698 45818 89796 45823
rect 88698 45250 88708 45818
rect 89786 45250 89796 45818
rect 88698 45245 89796 45250
rect 83036 43208 83064 43272
rect 88208 43208 88236 43272
rect 83036 43188 88236 43208
<< via3 >>
rect 39034 68250 39622 69308
rect 33042 64346 38186 64410
rect 33042 60054 38186 60118
rect 62460 59728 67604 59792
rect 61038 56780 61372 57236
rect 31770 55386 32028 55766
rect 33042 55762 38186 55826
rect 62460 55436 67604 55500
rect 33042 51470 38186 51534
rect 62460 51144 67604 51208
rect 82438 50454 82798 50666
rect 83064 47500 88208 47564
rect 33042 47178 38186 47242
rect 81270 45270 81936 46190
rect 83064 43208 88208 43272
<< mimcap >>
rect 33114 67086 38114 68498
rect 33114 65910 33154 67086
rect 38074 65910 38114 67086
rect 33114 64498 38114 65910
rect 33114 62794 38114 64206
rect 33114 61618 33154 62794
rect 38074 61618 38114 62794
rect 33114 60206 38114 61618
rect 62532 62468 67532 63880
rect 62532 61292 62572 62468
rect 67492 61292 67532 62468
rect 33114 58502 38114 59914
rect 62532 59880 67532 61292
rect 33114 57326 33154 58502
rect 38074 57326 38114 58502
rect 33114 55914 38114 57326
rect 62532 58176 67532 59588
rect 62532 57000 62572 58176
rect 67492 57000 67532 58176
rect 33114 54210 38114 55622
rect 62532 55588 67532 57000
rect 33114 53034 33154 54210
rect 38074 53034 38114 54210
rect 33114 51622 38114 53034
rect 62532 53884 67532 55296
rect 62532 52708 62572 53884
rect 67492 52708 67532 53884
rect 33114 49918 38114 51330
rect 62532 51296 67532 52708
rect 33114 48742 33154 49918
rect 38074 48742 38114 49918
rect 33114 47330 38114 48742
rect 83136 50240 88136 51652
rect 83136 49064 83176 50240
rect 88096 49064 88136 50240
rect 83136 47652 88136 49064
rect 83136 45948 88136 47360
rect 83136 44772 83176 45948
rect 88096 44772 88136 45948
rect 83136 43360 88136 44772
<< mimcapcontact >>
rect 33154 65910 38074 67086
rect 33154 61618 38074 62794
rect 62572 61292 67492 62468
rect 33154 57326 38074 58502
rect 62572 57000 67492 58176
rect 33154 53034 38074 54210
rect 62572 52708 67492 53884
rect 33154 48742 38074 49918
rect 83176 49064 88096 50240
rect 83176 44772 88096 45948
<< metal4 >>
rect 39033 69308 39623 69309
rect 39033 69224 39034 69308
rect 32146 68754 39034 69224
rect 32162 66698 32516 68754
rect 39033 68250 39034 68754
rect 39622 68250 39623 69308
rect 39033 68249 39623 68250
rect 33153 67086 38075 67087
rect 33153 66698 33154 67086
rect 32120 66696 33154 66698
rect 32098 66258 33154 66696
rect 32098 62508 32540 66258
rect 33153 65910 33154 66258
rect 38074 65910 38075 67086
rect 33153 65909 38075 65910
rect 33026 64410 38202 64426
rect 33026 64346 33042 64410
rect 38186 64346 38202 64410
rect 33026 64330 38202 64346
rect 33153 62794 38075 62795
rect 32094 62496 32598 62508
rect 33153 62496 33154 62794
rect 32094 62056 33154 62496
rect 32094 58138 32598 62056
rect 33153 61618 33154 62056
rect 38074 61618 38075 62794
rect 62571 62468 67493 62469
rect 33153 61617 38075 61618
rect 61604 62272 61972 62296
rect 62571 62272 62572 62468
rect 61604 61734 62572 62272
rect 33026 60118 38202 60134
rect 33026 60054 33042 60118
rect 38186 60054 38202 60118
rect 33026 60038 38202 60054
rect 33153 58502 38075 58503
rect 33153 58138 33154 58502
rect 32094 57698 33154 58138
rect 31769 55766 32029 55767
rect 31769 55386 31770 55766
rect 32028 55624 32029 55766
rect 32094 55624 32598 57698
rect 33153 57326 33154 57698
rect 38074 57326 38075 58502
rect 33153 57325 38075 57326
rect 61604 57832 61972 61734
rect 62571 61292 62572 61734
rect 67492 61292 67493 62468
rect 62571 61291 67493 61292
rect 62444 59792 67620 59808
rect 62444 59728 62460 59792
rect 67604 59728 67620 59792
rect 62444 59712 67620 59728
rect 62571 58176 67493 58177
rect 62571 57832 62572 58176
rect 61604 57294 62572 57832
rect 61037 57236 61373 57237
rect 61037 56780 61038 57236
rect 61372 57130 61373 57236
rect 61604 57130 61972 57294
rect 61372 56928 61972 57130
rect 62571 57000 62572 57294
rect 67492 57000 67493 58176
rect 62571 56999 67493 57000
rect 61372 56780 61373 56928
rect 61037 56779 61373 56780
rect 33026 55826 38202 55842
rect 33026 55762 33042 55826
rect 38186 55762 38202 55826
rect 33026 55746 38202 55762
rect 32028 55494 32598 55624
rect 32028 55386 32029 55494
rect 31769 55385 32029 55386
rect 32094 53846 32598 55494
rect 33153 54210 38075 54211
rect 33153 53846 33154 54210
rect 32094 53406 33154 53846
rect 32094 49554 32598 53406
rect 33153 53034 33154 53406
rect 38074 53034 38075 54210
rect 33153 53033 38075 53034
rect 61604 53566 61972 56928
rect 62444 55500 67620 55516
rect 62444 55436 62460 55500
rect 67604 55436 67620 55500
rect 62444 55420 67620 55436
rect 62571 53884 67493 53885
rect 62571 53566 62572 53884
rect 61604 53028 62572 53566
rect 61604 53026 61972 53028
rect 62571 52708 62572 53028
rect 67492 52708 67493 53884
rect 62571 52707 67493 52708
rect 33026 51534 38202 51550
rect 33026 51470 33042 51534
rect 38186 51470 38202 51534
rect 33026 51454 38202 51470
rect 62444 51208 67620 51224
rect 62444 51144 62460 51208
rect 67604 51144 67620 51208
rect 62444 51128 67620 51144
rect 82437 50666 82799 50667
rect 82437 50454 82438 50666
rect 82798 50454 82799 50666
rect 82437 50453 82799 50454
rect 82546 50030 82702 50453
rect 83175 50240 88097 50241
rect 82462 50010 82908 50030
rect 83175 50010 83176 50240
rect 33153 49918 38075 49919
rect 33153 49554 33154 49918
rect 32094 49114 33154 49554
rect 32094 49050 32598 49114
rect 33153 48742 33154 49114
rect 38074 48742 38075 49918
rect 33153 48741 38075 48742
rect 82462 49486 83176 50010
rect 82462 48376 82908 49486
rect 83175 49064 83176 49486
rect 88096 49064 88097 50240
rect 83175 49063 88097 49064
rect 82446 47596 82908 48376
rect 33026 47242 38202 47258
rect 33026 47178 33042 47242
rect 38186 47178 38202 47242
rect 33026 47162 38202 47178
rect 81269 46190 81937 46191
rect 81269 45270 81270 46190
rect 81936 46092 81937 46190
rect 82462 46092 82908 47596
rect 83048 47564 88224 47580
rect 83048 47500 83064 47564
rect 88208 47500 88224 47564
rect 83048 47484 88224 47500
rect 81936 45686 82908 46092
rect 83175 45948 88097 45949
rect 83175 45686 83176 45948
rect 81936 45642 83176 45686
rect 81936 45270 81937 45642
rect 81269 45269 81937 45270
rect 82462 45144 83176 45642
rect 83175 44772 83176 45144
rect 88096 44772 88097 45948
rect 83175 44771 88097 44772
rect 83048 43272 88224 43288
rect 83048 43208 83064 43272
rect 88208 43208 88224 43272
rect 83048 43192 88224 43208
<< labels >>
flabel poly 30710 44036 30710 44036 0 FreeSans 4800 0 0 0 vin1
flabel metal1 21456 45972 21456 45972 0 FreeSans 1600 0 0 0 vout
flabel locali 21634 55558 21634 55558 0 FreeSans 1600 0 0 0 vout1
flabel locali 61674 46392 61674 46392 0 FreeSans 1600 0 0 0 vout2
flabel metal1 4286 77500 4286 77500 0 FreeSans 1600 0 0 0 vdda
rlabel metal3 88528 47472 88528 47472 5 bot
flabel locali 76018 49066 76018 49066 0 FreeSans 1600 0 0 0 vout3
flabel metal1 86350 53606 86350 53606 0 FreeSans 800 0 0 0 dfout
flabel metal1 83702 53468 83702 53468 0 FreeSans 800 0 0 0 reset
flabel metal1 83258 53670 83258 53670 0 FreeSans 800 0 0 0 clkin
flabel metal1 1910 -6426 1910 -6426 0 FreeSans 1600 0 0 0 vssa
flabel metal1 46520 2470 46520 2470 0 FreeSans 1600 0 0 0 vcap
flabel poly 80634 26412 80658 26412 0 FreeSans 1600 0 0 0 vin2
flabel locali 67518 3174 67518 3174 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_0/nmos5555_0/d
flabel locali 62016 8226 62016 8226 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_0/nmos5555_0/s
flabel poly 66228 8416 66228 8416 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_0/nmos5555_0/g
flabel locali 67518 9032 67518 9032 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_0/nmos5555_1/d
flabel locali 62016 14084 62016 14084 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_0/nmos5555_1/s
flabel poly 66228 14274 66228 14274 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_0/nmos5555_1/g
flabel locali 67518 14890 67518 14890 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_0/nmos5555_2/d
flabel locali 62016 19942 62016 19942 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_0/nmos5555_2/s
flabel poly 66228 20132 66228 20132 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_0/nmos5555_2/g
flabel locali 67512 20728 67512 20728 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_0/nmos5555_3/d
flabel locali 62010 25780 62010 25780 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_0/nmos5555_3/s
flabel poly 66222 25970 66222 25970 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_0/nmos5555_3/g
flabel locali 73990 3172 73990 3172 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_0/nmos5555_4/d
flabel locali 68488 8224 68488 8224 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_0/nmos5555_4/s
flabel poly 72700 8414 72700 8414 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_0/nmos5555_4/g
flabel locali 73986 9030 73986 9030 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_0/nmos5555_5/d
flabel locali 68484 14082 68484 14082 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_0/nmos5555_5/s
flabel poly 72696 14272 72696 14272 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_0/nmos5555_5/g
flabel locali 73982 14902 73982 14902 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_0/nmos5555_6/d
flabel locali 68480 19954 68480 19954 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_0/nmos5555_6/s
flabel poly 72692 20144 72692 20144 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_0/nmos5555_6/g
flabel locali 73974 20726 73974 20726 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_0/nmos5555_7/d
flabel locali 68472 25778 68472 25778 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_0/nmos5555_7/s
flabel poly 72684 25968 72684 25968 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_0/nmos5555_7/g
flabel locali 80674 3146 80674 3146 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_1/nmos5555_0/d
flabel locali 75172 8198 75172 8198 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_1/nmos5555_0/s
flabel poly 79384 8388 79384 8388 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_1/nmos5555_0/g
flabel locali 80674 9004 80674 9004 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_1/nmos5555_1/d
flabel locali 75172 14056 75172 14056 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_1/nmos5555_1/s
flabel poly 79384 14246 79384 14246 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_1/nmos5555_1/g
flabel locali 80674 14862 80674 14862 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_1/nmos5555_2/d
flabel locali 75172 19914 75172 19914 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_1/nmos5555_2/s
flabel poly 79384 20104 79384 20104 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_1/nmos5555_2/g
flabel locali 80668 20700 80668 20700 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_1/nmos5555_3/d
flabel locali 75166 25752 75166 25752 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_1/nmos5555_3/s
flabel poly 79378 25942 79378 25942 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_1/nmos5555_3/g
flabel locali 87146 3144 87146 3144 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_1/nmos5555_4/d
flabel locali 81644 8196 81644 8196 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_1/nmos5555_4/s
flabel poly 85856 8386 85856 8386 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_1/nmos5555_4/g
flabel locali 87142 9002 87142 9002 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_1/nmos5555_5/d
flabel locali 81640 14054 81640 14054 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_1/nmos5555_5/s
flabel poly 85852 14244 85852 14244 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_1/nmos5555_5/g
flabel locali 87138 14874 87138 14874 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_1/nmos5555_6/d
flabel locali 81636 19926 81636 19926 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_1/nmos5555_6/s
flabel poly 85848 20116 85848 20116 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_1/nmos5555_6/g
flabel locali 87130 20698 87130 20698 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_1/nmos5555_7/d
flabel locali 81628 25750 81628 25750 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_1/nmos5555_7/s
flabel poly 85840 25940 85840 25940 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_1/nmos5555_7/g
flabel locali 93908 3138 93908 3138 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_2/nmos5555_0/d
flabel locali 88406 8190 88406 8190 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_2/nmos5555_0/s
flabel poly 92618 8380 92618 8380 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_2/nmos5555_0/g
flabel locali 93908 8996 93908 8996 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_2/nmos5555_1/d
flabel locali 88406 14048 88406 14048 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_2/nmos5555_1/s
flabel poly 92618 14238 92618 14238 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_2/nmos5555_1/g
flabel locali 93908 14854 93908 14854 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_2/nmos5555_2/d
flabel locali 88406 19906 88406 19906 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_2/nmos5555_2/s
flabel poly 92618 20096 92618 20096 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_2/nmos5555_2/g
flabel locali 93902 20692 93902 20692 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_2/nmos5555_3/d
flabel locali 88400 25744 88400 25744 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_2/nmos5555_3/s
flabel poly 92612 25934 92612 25934 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_2/nmos5555_3/g
flabel locali 100380 3136 100380 3136 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_2/nmos5555_4/d
flabel locali 94878 8188 94878 8188 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_2/nmos5555_4/s
flabel poly 99090 8378 99090 8378 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_2/nmos5555_4/g
flabel locali 100376 8994 100376 8994 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_2/nmos5555_5/d
flabel locali 94874 14046 94874 14046 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_2/nmos5555_5/s
flabel poly 99086 14236 99086 14236 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_2/nmos5555_5/g
flabel locali 100372 14866 100372 14866 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_2/nmos5555_6/d
flabel locali 94870 19918 94870 19918 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_2/nmos5555_6/s
flabel poly 99082 20108 99082 20108 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_2/nmos5555_6/g
flabel locali 100364 20690 100364 20690 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_2/nmos5555_7/d
flabel locali 94862 25742 94862 25742 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_2/nmos5555_7/s
flabel poly 99074 25932 99074 25932 0 FreeSans 1600 0 0 0 nmos551020guard_0/nmos551020_2/nmos5555_7/g
flabel locali 83760 39310 83760 39310 0 FreeSans 1600 0 0 0 nmos3346guard_0/nmos3346_2/d
flabel poly 85250 39378 85250 39378 0 FreeSans 1600 0 0 0 nmos3346guard_0/nmos3346_2/g
flabel locali 84868 35144 84868 35144 0 FreeSans 1600 0 0 0 nmos3346guard_0/nmos3346_2/s
flabel metal1 83366 38924 83366 38924 0 FreeSans 1600 0 0 0 nmos3346guard_0/nmos3346_2/sub
flabel locali 77124 39316 77124 39316 0 FreeSans 1600 0 0 0 nmos3346guard_0/nmos3346_0/d
flabel poly 78614 39384 78614 39384 0 FreeSans 1600 0 0 0 nmos3346guard_0/nmos3346_0/g
flabel locali 78232 35150 78232 35150 0 FreeSans 1600 0 0 0 nmos3346guard_0/nmos3346_0/s
flabel metal1 76730 38930 76730 38930 0 FreeSans 1600 0 0 0 nmos3346guard_0/nmos3346_0/sub
flabel locali 80450 39310 80450 39310 0 FreeSans 1600 0 0 0 nmos3346guard_0/nmos3346_1/d
flabel poly 81940 39378 81940 39378 0 FreeSans 1600 0 0 0 nmos3346guard_0/nmos3346_1/g
flabel locali 81558 35144 81558 35144 0 FreeSans 1600 0 0 0 nmos3346guard_0/nmos3346_1/s
flabel metal1 80056 38924 80056 38924 0 FreeSans 1600 0 0 0 nmos3346guard_0/nmos3346_1/sub
flabel locali 74046 73256 74046 73256 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_0/pmos3345_5/s
flabel locali 73378 70036 73378 70036 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_0/pmos3345_5/d
flabel poly 72378 73386 72378 73386 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_0/pmos3345_5/g
flabel locali 74042 69480 74042 69480 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_0/pmos3345_4/s
flabel locali 73374 66260 73374 66260 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_0/pmos3345_4/d
flabel poly 72374 69610 72374 69610 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_0/pmos3345_4/g
flabel locali 74042 65710 74042 65710 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_0/pmos3345_3/s
flabel locali 73374 62490 73374 62490 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_0/pmos3345_3/d
flabel poly 72374 65840 72374 65840 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_0/pmos3345_3/g
flabel locali 74042 61946 74042 61946 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_0/pmos3345_2/s
flabel locali 73374 58726 73374 58726 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_0/pmos3345_2/d
flabel poly 72374 62076 72374 62076 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_0/pmos3345_2/g
flabel locali 74042 58170 74042 58170 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_0/pmos3345_1/s
flabel locali 73374 54950 73374 54950 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_0/pmos3345_1/d
flabel poly 72374 58300 72374 58300 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_0/pmos3345_1/g
flabel locali 74046 54398 74046 54398 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_0/pmos3345_0/s
flabel locali 73378 51178 73378 51178 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_0/pmos3345_0/d
flabel poly 72378 54528 72378 54528 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_0/pmos3345_0/g
flabel locali 77910 73236 77910 73236 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_1/pmos3345_5/s
flabel locali 77242 70016 77242 70016 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_1/pmos3345_5/d
flabel poly 76242 73366 76242 73366 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_1/pmos3345_5/g
flabel locali 77906 69460 77906 69460 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_1/pmos3345_4/s
flabel locali 77238 66240 77238 66240 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_1/pmos3345_4/d
flabel poly 76238 69590 76238 69590 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_1/pmos3345_4/g
flabel locali 77906 65690 77906 65690 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_1/pmos3345_3/s
flabel locali 77238 62470 77238 62470 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_1/pmos3345_3/d
flabel poly 76238 65820 76238 65820 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_1/pmos3345_3/g
flabel locali 77906 61926 77906 61926 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_1/pmos3345_2/s
flabel locali 77238 58706 77238 58706 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_1/pmos3345_2/d
flabel poly 76238 62056 76238 62056 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_1/pmos3345_2/g
flabel locali 77906 58150 77906 58150 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_1/pmos3345_1/s
flabel locali 77238 54930 77238 54930 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_1/pmos3345_1/d
flabel poly 76238 58280 76238 58280 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_1/pmos3345_1/g
flabel locali 77910 54378 77910 54378 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_1/pmos3345_0/s
flabel locali 77242 51158 77242 51158 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_1/pmos3345_0/d
flabel poly 76242 54508 76242 54508 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_1/pmos3345_0/g
flabel locali 81760 73250 81760 73250 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_2/pmos3345_5/s
flabel locali 81092 70030 81092 70030 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_2/pmos3345_5/d
flabel poly 80092 73380 80092 73380 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_2/pmos3345_5/g
flabel locali 81756 69474 81756 69474 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_2/pmos3345_4/s
flabel locali 81088 66254 81088 66254 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_2/pmos3345_4/d
flabel poly 80088 69604 80088 69604 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_2/pmos3345_4/g
flabel locali 81756 65704 81756 65704 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_2/pmos3345_3/s
flabel locali 81088 62484 81088 62484 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_2/pmos3345_3/d
flabel poly 80088 65834 80088 65834 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_2/pmos3345_3/g
flabel locali 81756 61940 81756 61940 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_2/pmos3345_2/s
flabel locali 81088 58720 81088 58720 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_2/pmos3345_2/d
flabel poly 80088 62070 80088 62070 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_2/pmos3345_2/g
flabel locali 81756 58164 81756 58164 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_2/pmos3345_1/s
flabel locali 81088 54944 81088 54944 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_2/pmos3345_1/d
flabel poly 80088 58294 80088 58294 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_2/pmos3345_1/g
flabel locali 81760 54392 81760 54392 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_2/pmos3345_0/s
flabel locali 81092 51172 81092 51172 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_2/pmos3345_0/d
flabel poly 80092 54522 80092 54522 0 FreeSans 1600 0 0 0 pmos33431guard_0/pmos33431_2/pmos3345_0/g
flabel locali 20714 59322 20714 59322 0 FreeSans 1600 0 0 0 pmos33823guard_0/d
flabel locali 18562 59764 18562 59764 0 FreeSans 1600 0 0 0 pmos33823guard_0/sub
flabel poly 20690 55516 20690 55516 0 FreeSans 1600 0 0 0 pmos33823guard_0/g
flabel metal1 18770 53884 18770 53884 0 FreeSans 1600 0 0 0 pmos33823guard_0/s
flabel locali 30178 55640 30178 55640 0 FreeSans 1600 0 0 0 nmos33210guard_0/d
flabel locali 23346 54920 23346 54920 0 FreeSans 1600 0 0 0 nmos33210guard_0/s
flabel poly 30404 54952 30404 54952 0 FreeSans 1600 0 0 0 nmos33210guard_0/g
flabel locali 29658 54032 29658 54032 0 FreeSans 1600 0 0 0 nmos33210guard_0/sub
rlabel metal4 32340 58294 32340 58294 3 cap5p_0/top
rlabel metal3 38766 56832 38766 56832 3 cap5p_0/bot
flabel locali 57760 64534 57760 64534 0 FreeSans 1600 0 0 0 pmos331020guard_0/d
flabel locali 57802 57040 57802 57040 0 FreeSans 1600 0 0 0 pmos331020guard_0/s
flabel locali 53526 65020 53526 65020 0 FreeSans 1600 0 0 0 pmos331020guard_0/sub
flabel poly 57946 61004 57946 61004 0 FreeSans 1600 0 0 0 pmos331020guard_0/g
rlabel metal3 68498 57998 68498 57998 3 cap3p_0/bot
rlabel metal4 61752 57942 61752 57942 3 cap3p_0/top
flabel poly 67860 43534 67860 43534 0 FreeSans 1600 0 0 0 nmos3355guard_0/g
flabel locali 66306 43396 66306 43396 0 FreeSans 1600 0 0 0 nmos3355guard_0/d
flabel locali 69622 43428 69622 43428 0 FreeSans 1600 0 0 0 nmos3355guard_0/s
flabel locali 65984 42764 65984 42764 0 FreeSans 1600 0 0 0 nmos3355guard_0/sub
rlabel comment 83272 53268 83272 53268 4 sky130_fd_sc_hvl__dfrtp_1_0/dfrtp_1
flabel metal1 83272 53319 86344 53393 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__dfrtp_1_0/VGND
flabel metal1 83272 53268 86344 53291 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__dfrtp_1_0/VNB
flabel metal1 83272 53957 86344 54031 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__dfrtp_1_0/VPWR
flabel metal1 83272 54059 86344 54082 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__dfrtp_1_0/VPB
flabel locali 83975 53436 84009 53470 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__dfrtp_1_0/D
flabel locali 83975 53510 84009 53544 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__dfrtp_1_0/D
flabel locali 83975 53584 84009 53618 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__dfrtp_1_0/D
flabel locali 83399 53510 83433 53544 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__dfrtp_1_0/CLK
flabel locali 83399 53584 83433 53618 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__dfrtp_1_0/CLK
flabel locali 83399 53658 83433 53692 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__dfrtp_1_0/CLK
flabel locali 83879 53732 83913 53766 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__dfrtp_1_0/RESET_B
flabel locali 86279 53436 86313 53470 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__dfrtp_1_0/Q
flabel locali 86279 53510 86313 53544 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__dfrtp_1_0/Q
flabel locali 86279 53584 86313 53618 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__dfrtp_1_0/Q
flabel locali 86279 53658 86313 53692 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__dfrtp_1_0/Q
flabel locali 86279 53732 86313 53766 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__dfrtp_1_0/Q
flabel locali 86279 53806 86313 53840 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__dfrtp_1_0/Q
flabel locali 86279 53880 86313 53914 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__dfrtp_1_0/Q
flabel poly 30500 43816 30500 43816 0 FreeSans 3200 0 0 0 nmos551535_0/g
flabel locali 39832 43608 39832 43608 0 FreeSans 3200 0 0 0 nmos551535_0/S
flabel locali 21058 43282 21058 43282 0 FreeSans 3200 0 0 0 nmos551535_0/D
flabel locali 59492 38270 59492 38270 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_3/nmos5555_6/d
flabel locali 53990 43322 53990 43322 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_3/nmos5555_6/s
flabel poly 58202 43512 58202 43512 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_3/nmos5555_6/g
flabel locali 59492 32454 59492 32454 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_3/nmos5555_5/d
flabel locali 53990 37506 53990 37506 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_3/nmos5555_5/s
flabel poly 58202 37696 58202 37696 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_3/nmos5555_5/g
flabel locali 59492 26620 59492 26620 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_3/nmos5555_4/d
flabel locali 53990 31672 53990 31672 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_3/nmos5555_4/s
flabel poly 58202 31862 58202 31862 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_3/nmos5555_4/g
flabel locali 59492 20784 59492 20784 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_3/nmos5555_3/d
flabel locali 53990 25836 53990 25836 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_3/nmos5555_3/s
flabel poly 58202 26026 58202 26026 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_3/nmos5555_3/g
flabel locali 59492 14920 59492 14920 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_3/nmos5555_2/d
flabel locali 53990 19972 53990 19972 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_3/nmos5555_2/s
flabel poly 58202 20162 58202 20162 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_3/nmos5555_2/g
flabel locali 59502 9064 59502 9064 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_3/nmos5555_1/d
flabel locali 54000 14116 54000 14116 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_3/nmos5555_1/s
flabel poly 58212 14306 58212 14306 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_3/nmos5555_1/g
flabel locali 59520 3156 59520 3156 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_3/nmos5555_0/d
flabel locali 54018 8208 54018 8208 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_3/nmos5555_0/s
flabel poly 58230 8398 58230 8398 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_3/nmos5555_0/g
flabel locali 52978 38256 52978 38256 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_2/nmos5555_6/d
flabel locali 47476 43308 47476 43308 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_2/nmos5555_6/s
flabel poly 51688 43498 51688 43498 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_2/nmos5555_6/g
flabel locali 52978 32440 52978 32440 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_2/nmos5555_5/d
flabel locali 47476 37492 47476 37492 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_2/nmos5555_5/s
flabel poly 51688 37682 51688 37682 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_2/nmos5555_5/g
flabel locali 52978 26606 52978 26606 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_2/nmos5555_4/d
flabel locali 47476 31658 47476 31658 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_2/nmos5555_4/s
flabel poly 51688 31848 51688 31848 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_2/nmos5555_4/g
flabel locali 52978 20770 52978 20770 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_2/nmos5555_3/d
flabel locali 47476 25822 47476 25822 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_2/nmos5555_3/s
flabel poly 51688 26012 51688 26012 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_2/nmos5555_3/g
flabel locali 52978 14906 52978 14906 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_2/nmos5555_2/d
flabel locali 47476 19958 47476 19958 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_2/nmos5555_2/s
flabel poly 51688 20148 51688 20148 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_2/nmos5555_2/g
flabel locali 52988 9050 52988 9050 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_2/nmos5555_1/d
flabel locali 47486 14102 47486 14102 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_2/nmos5555_1/s
flabel poly 51698 14292 51698 14292 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_2/nmos5555_1/g
flabel locali 53006 3142 53006 3142 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_2/nmos5555_0/d
flabel locali 47504 8194 47504 8194 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_2/nmos5555_0/s
flabel poly 51716 8384 51716 8384 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_2/nmos5555_0/g
flabel locali 46390 38234 46390 38234 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_1/nmos5555_6/d
flabel locali 40888 43286 40888 43286 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_1/nmos5555_6/s
flabel poly 45100 43476 45100 43476 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_1/nmos5555_6/g
flabel locali 46390 32418 46390 32418 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_1/nmos5555_5/d
flabel locali 40888 37470 40888 37470 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_1/nmos5555_5/s
flabel poly 45100 37660 45100 37660 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_1/nmos5555_5/g
flabel locali 46390 26584 46390 26584 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_1/nmos5555_4/d
flabel locali 40888 31636 40888 31636 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_1/nmos5555_4/s
flabel poly 45100 31826 45100 31826 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_1/nmos5555_4/g
flabel locali 46390 20748 46390 20748 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_1/nmos5555_3/d
flabel locali 40888 25800 40888 25800 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_1/nmos5555_3/s
flabel poly 45100 25990 45100 25990 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_1/nmos5555_3/g
flabel locali 46390 14884 46390 14884 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_1/nmos5555_2/d
flabel locali 40888 19936 40888 19936 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_1/nmos5555_2/s
flabel poly 45100 20126 45100 20126 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_1/nmos5555_2/g
flabel locali 46400 9028 46400 9028 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_1/nmos5555_1/d
flabel locali 40898 14080 40898 14080 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_1/nmos5555_1/s
flabel poly 45110 14270 45110 14270 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_1/nmos5555_1/g
flabel locali 46418 3120 46418 3120 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_1/nmos5555_0/d
flabel locali 40916 8172 40916 8172 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_1/nmos5555_0/s
flabel poly 45128 8362 45128 8362 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_1/nmos5555_0/g
flabel locali 39900 38234 39900 38234 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_0/nmos5555_6/d
flabel locali 34398 43286 34398 43286 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_0/nmos5555_6/s
flabel poly 38610 43476 38610 43476 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_0/nmos5555_6/g
flabel locali 39900 32418 39900 32418 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_0/nmos5555_5/d
flabel locali 34398 37470 34398 37470 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_0/nmos5555_5/s
flabel poly 38610 37660 38610 37660 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_0/nmos5555_5/g
flabel locali 39900 26584 39900 26584 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_0/nmos5555_4/d
flabel locali 34398 31636 34398 31636 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_0/nmos5555_4/s
flabel poly 38610 31826 38610 31826 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_0/nmos5555_4/g
flabel locali 39900 20748 39900 20748 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_0/nmos5555_3/d
flabel locali 34398 25800 34398 25800 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_0/nmos5555_3/s
flabel poly 38610 25990 38610 25990 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_0/nmos5555_3/g
flabel locali 39900 14884 39900 14884 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_0/nmos5555_2/d
flabel locali 34398 19936 34398 19936 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_0/nmos5555_2/s
flabel poly 38610 20126 38610 20126 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_0/nmos5555_2/g
flabel locali 39910 9028 39910 9028 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_0/nmos5555_1/d
flabel locali 34408 14080 34408 14080 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_0/nmos5555_1/s
flabel poly 38620 14270 38620 14270 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_0/nmos5555_1/g
flabel locali 39928 3120 39928 3120 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_0/nmos5555_0/d
flabel locali 34426 8172 34426 8172 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_0/nmos5555_0/s
flabel poly 38638 8362 38638 8362 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_0/nmos5555_0/g
flabel locali 33390 38228 33390 38228 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_8/nmos5555_6/d
flabel locali 27888 43280 27888 43280 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_8/nmos5555_6/s
flabel poly 32100 43470 32100 43470 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_8/nmos5555_6/g
flabel locali 33390 32412 33390 32412 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_8/nmos5555_5/d
flabel locali 27888 37464 27888 37464 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_8/nmos5555_5/s
flabel poly 32100 37654 32100 37654 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_8/nmos5555_5/g
flabel locali 33390 26578 33390 26578 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_8/nmos5555_4/d
flabel locali 27888 31630 27888 31630 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_8/nmos5555_4/s
flabel poly 32100 31820 32100 31820 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_8/nmos5555_4/g
flabel locali 33390 20742 33390 20742 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_8/nmos5555_3/d
flabel locali 27888 25794 27888 25794 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_8/nmos5555_3/s
flabel poly 32100 25984 32100 25984 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_8/nmos5555_3/g
flabel locali 33390 14878 33390 14878 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_8/nmos5555_2/d
flabel locali 27888 19930 27888 19930 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_8/nmos5555_2/s
flabel poly 32100 20120 32100 20120 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_8/nmos5555_2/g
flabel locali 33400 9022 33400 9022 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_8/nmos5555_1/d
flabel locali 27898 14074 27898 14074 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_8/nmos5555_1/s
flabel poly 32110 14264 32110 14264 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_8/nmos5555_1/g
flabel locali 33418 3114 33418 3114 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_8/nmos5555_0/d
flabel locali 27916 8166 27916 8166 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_8/nmos5555_0/s
flabel poly 32128 8356 32128 8356 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_8/nmos5555_0/g
flabel locali 26868 38212 26868 38212 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_7/nmos5555_6/d
flabel locali 21366 43264 21366 43264 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_7/nmos5555_6/s
flabel poly 25578 43454 25578 43454 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_7/nmos5555_6/g
flabel locali 26868 32396 26868 32396 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_7/nmos5555_5/d
flabel locali 21366 37448 21366 37448 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_7/nmos5555_5/s
flabel poly 25578 37638 25578 37638 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_7/nmos5555_5/g
flabel locali 26868 26562 26868 26562 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_7/nmos5555_4/d
flabel locali 21366 31614 21366 31614 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_7/nmos5555_4/s
flabel poly 25578 31804 25578 31804 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_7/nmos5555_4/g
flabel locali 26868 20726 26868 20726 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_7/nmos5555_3/d
flabel locali 21366 25778 21366 25778 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_7/nmos5555_3/s
flabel poly 25578 25968 25578 25968 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_7/nmos5555_3/g
flabel locali 26868 14862 26868 14862 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_7/nmos5555_2/d
flabel locali 21366 19914 21366 19914 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_7/nmos5555_2/s
flabel poly 25578 20104 25578 20104 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_7/nmos5555_2/g
flabel locali 26878 9006 26878 9006 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_7/nmos5555_1/d
flabel locali 21376 14058 21376 14058 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_7/nmos5555_1/s
flabel poly 25588 14248 25588 14248 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_7/nmos5555_1/g
flabel locali 26896 3098 26896 3098 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_7/nmos5555_0/d
flabel locali 21394 8150 21394 8150 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_7/nmos5555_0/s
flabel poly 25606 8340 25606 8340 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_7/nmos5555_0/g
flabel locali 20378 38228 20378 38228 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_6/nmos5555_6/d
flabel locali 14876 43280 14876 43280 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_6/nmos5555_6/s
flabel poly 19088 43470 19088 43470 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_6/nmos5555_6/g
flabel locali 20378 32412 20378 32412 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_6/nmos5555_5/d
flabel locali 14876 37464 14876 37464 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_6/nmos5555_5/s
flabel poly 19088 37654 19088 37654 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_6/nmos5555_5/g
flabel locali 20378 26578 20378 26578 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_6/nmos5555_4/d
flabel locali 14876 31630 14876 31630 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_6/nmos5555_4/s
flabel poly 19088 31820 19088 31820 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_6/nmos5555_4/g
flabel locali 20378 20742 20378 20742 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_6/nmos5555_3/d
flabel locali 14876 25794 14876 25794 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_6/nmos5555_3/s
flabel poly 19088 25984 19088 25984 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_6/nmos5555_3/g
flabel locali 20378 14878 20378 14878 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_6/nmos5555_2/d
flabel locali 14876 19930 14876 19930 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_6/nmos5555_2/s
flabel poly 19088 20120 19088 20120 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_6/nmos5555_2/g
flabel locali 20388 9022 20388 9022 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_6/nmos5555_1/d
flabel locali 14886 14074 14886 14074 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_6/nmos5555_1/s
flabel poly 19098 14264 19098 14264 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_6/nmos5555_1/g
flabel locali 20406 3114 20406 3114 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_6/nmos5555_0/d
flabel locali 14904 8166 14904 8166 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_6/nmos5555_0/s
flabel poly 19116 8356 19116 8356 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_6/nmos5555_0/g
flabel locali 13872 38220 13872 38220 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_5/nmos5555_6/d
flabel locali 8370 43272 8370 43272 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_5/nmos5555_6/s
flabel poly 12582 43462 12582 43462 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_5/nmos5555_6/g
flabel locali 13872 32404 13872 32404 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_5/nmos5555_5/d
flabel locali 8370 37456 8370 37456 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_5/nmos5555_5/s
flabel poly 12582 37646 12582 37646 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_5/nmos5555_5/g
flabel locali 13872 26570 13872 26570 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_5/nmos5555_4/d
flabel locali 8370 31622 8370 31622 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_5/nmos5555_4/s
flabel poly 12582 31812 12582 31812 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_5/nmos5555_4/g
flabel locali 13872 20734 13872 20734 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_5/nmos5555_3/d
flabel locali 8370 25786 8370 25786 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_5/nmos5555_3/s
flabel poly 12582 25976 12582 25976 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_5/nmos5555_3/g
flabel locali 13872 14870 13872 14870 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_5/nmos5555_2/d
flabel locali 8370 19922 8370 19922 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_5/nmos5555_2/s
flabel poly 12582 20112 12582 20112 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_5/nmos5555_2/g
flabel locali 13882 9014 13882 9014 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_5/nmos5555_1/d
flabel locali 8380 14066 8380 14066 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_5/nmos5555_1/s
flabel poly 12592 14256 12592 14256 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_5/nmos5555_1/g
flabel locali 13900 3106 13900 3106 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_5/nmos5555_0/d
flabel locali 8398 8158 8398 8158 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_5/nmos5555_0/s
flabel poly 12610 8348 12610 8348 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_5/nmos5555_0/g
flabel locali 7358 38212 7358 38212 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_4/nmos5555_6/d
flabel locali 1856 43264 1856 43264 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_4/nmos5555_6/s
flabel poly 6068 43454 6068 43454 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_4/nmos5555_6/g
flabel locali 7358 32396 7358 32396 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_4/nmos5555_5/d
flabel locali 1856 37448 1856 37448 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_4/nmos5555_5/s
flabel poly 6068 37638 6068 37638 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_4/nmos5555_5/g
flabel locali 7358 26562 7358 26562 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_4/nmos5555_4/d
flabel locali 1856 31614 1856 31614 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_4/nmos5555_4/s
flabel poly 6068 31804 6068 31804 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_4/nmos5555_4/g
flabel locali 7358 20726 7358 20726 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_4/nmos5555_3/d
flabel locali 1856 25778 1856 25778 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_4/nmos5555_3/s
flabel poly 6068 25968 6068 25968 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_4/nmos5555_3/g
flabel locali 7358 14862 7358 14862 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_4/nmos5555_2/d
flabel locali 1856 19914 1856 19914 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_4/nmos5555_2/s
flabel poly 6068 20104 6068 20104 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_4/nmos5555_2/g
flabel locali 7368 9006 7368 9006 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_4/nmos5555_1/d
flabel locali 1866 14058 1866 14058 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_4/nmos5555_1/s
flabel poly 6078 14248 6078 14248 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_4/nmos5555_1/g
flabel locali 7386 3098 7386 3098 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_4/nmos5555_0/d
flabel locali 1884 8150 1884 8150 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_4/nmos5555_0/s
flabel poly 6096 8340 6096 8340 0 FreeSans 1600 0 0 0 nmos551535_0/nmos55535_4/nmos5555_0/g
<< end >>
