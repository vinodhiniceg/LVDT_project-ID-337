magic
tech sky130A
timestamp 1634553547
<< pwell >>
rect 162 12816 703 12830
rect 19731 12816 20496 12830
rect 162 12448 20496 12816
rect 162 12268 703 12448
rect 19731 12200 20496 12448
rect 187 -30 20450 338
<< mvpsubdiff >>
rect 162 12816 703 12830
rect 162 12483 20425 12816
rect 162 12448 20459 12483
rect 162 12268 703 12448
rect 194 338 701 12268
rect 19952 11642 20459 12448
rect 19952 9716 20093 11642
rect 20349 9716 20459 11642
rect 19952 8603 20459 9716
rect 19952 6544 20082 8603
rect 20327 6544 20459 8603
rect 19952 5898 20459 6544
rect 19952 3806 20104 5898
rect 20349 3806 20459 5898
rect 19952 2782 20459 3806
rect 19952 723 20126 2782
rect 20316 723 20459 2782
rect 19952 338 20459 723
rect 187 253 20459 338
rect 187 -30 20450 253
<< mvpsubdiffcont >>
rect 20093 9716 20349 11642
rect 20082 6544 20327 8603
rect 20104 3806 20349 5898
rect 20126 723 20316 2782
<< polycont >>
rect 3526 12142 3875 12208
rect 16730 12126 16946 12192
<< locali >>
rect 3506 12208 3889 12222
rect 3506 12142 3526 12208
rect 3875 12142 3889 12208
rect 3506 12128 3889 12142
rect 16707 12192 16972 12206
rect 3663 11899 3772 12128
rect 16707 12126 16730 12192
rect 16946 12126 16972 12192
rect 16707 12115 16972 12126
rect 6659 11962 6696 11965
rect 6125 11911 6696 11962
rect 6659 11774 6696 11911
rect 16804 11887 16918 12115
rect 19302 11961 19900 11967
rect 19302 11887 19911 11961
rect 19832 11733 19911 11887
rect 20071 11642 20393 11831
rect 20071 9716 20093 11642
rect 20349 11564 20393 11642
rect 20371 9928 20393 11564
rect 20349 9716 20393 9928
rect 20071 9571 20393 9716
rect 20048 8603 20371 8681
rect 20048 6544 20082 8603
rect 20327 6544 20371 8603
rect 20048 6488 20371 6544
rect 20048 5898 20382 5999
rect 20048 3806 20104 5898
rect 20349 3806 20382 5898
rect 20048 3695 20382 3806
rect 20037 2782 20382 2904
rect 20037 723 20126 2782
rect 20316 723 20382 2782
rect 20037 634 20382 723
<< viali >>
rect 3583 12156 3823 12205
rect 16764 12143 16929 12183
rect 20126 9928 20349 11564
rect 20349 9928 20371 11564
rect 20104 6744 20293 8536
rect 20171 3928 20282 5776
rect 20182 845 20282 2682
<< metal1 >>
rect 3506 12205 3889 12222
rect 3506 12156 3583 12205
rect 3823 12156 3889 12205
rect 3506 12128 3889 12156
rect 16707 12183 16972 12206
rect 16707 12143 16764 12183
rect 16929 12143 16972 12183
rect 16707 12115 16972 12143
rect 20071 11564 20393 11831
rect 20071 11223 20126 11564
rect 19849 11160 20126 11223
rect 488 10625 806 10688
rect 20071 9928 20126 11160
rect 20371 9928 20393 11564
rect 20071 9571 20393 9928
rect 20048 8536 20371 8681
rect 20048 6744 20104 8536
rect 20293 6744 20371 8536
rect 20048 6488 20371 6744
rect 20048 5776 20382 5999
rect 20048 3928 20171 5776
rect 20282 3928 20382 5776
rect 20048 3695 20382 3928
rect 20037 2682 20382 2904
rect 20037 845 20182 2682
rect 20282 845 20382 2682
rect 20037 634 20382 845
use nmos551020  nmos551020_2
timestamp 1634552665
transform 1 0 13605 0 1 444
box -410 -462 6891 12086
use nmos551020  nmos551020_1
timestamp 1634552665
transform 1 0 6988 0 1 448
box -410 -462 6891 12086
use nmos551020  nmos551020_0
timestamp 1634552665
transform 1 0 410 0 1 462
box -410 -462 6891 12086
<< end >>
