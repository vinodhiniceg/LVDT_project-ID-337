magic
tech sky130A
magscale 1 2
timestamp 1634127529
<< mvnmos >>
rect -958 2823 -358 3423
rect -300 2823 300 3423
rect 358 2823 958 3423
rect -958 2129 -358 2729
rect -300 2129 300 2729
rect 358 2129 958 2729
rect -958 1435 -358 2035
rect -300 1435 300 2035
rect 358 1435 958 2035
rect -958 741 -358 1341
rect -300 741 300 1341
rect 358 741 958 1341
rect -958 47 -358 647
rect -300 47 300 647
rect 358 47 958 647
rect -958 -647 -358 -47
rect -300 -647 300 -47
rect 358 -647 958 -47
rect -958 -1341 -358 -741
rect -300 -1341 300 -741
rect 358 -1341 958 -741
rect -958 -2035 -358 -1435
rect -300 -2035 300 -1435
rect 358 -2035 958 -1435
rect -958 -2729 -358 -2129
rect -300 -2729 300 -2129
rect 358 -2729 958 -2129
rect -958 -3423 -358 -2823
rect -300 -3423 300 -2823
rect 358 -3423 958 -2823
<< mvndiff >>
rect -1016 3209 -958 3423
rect -1016 3037 -1004 3209
rect -970 3037 -958 3209
rect -1016 2823 -958 3037
rect -358 3209 -300 3423
rect -358 3037 -346 3209
rect -312 3037 -300 3209
rect -358 2823 -300 3037
rect 300 3209 358 3423
rect 300 3037 312 3209
rect 346 3037 358 3209
rect 300 2823 358 3037
rect 958 3209 1016 3423
rect 958 3037 970 3209
rect 1004 3037 1016 3209
rect 958 2823 1016 3037
rect -1016 2515 -958 2729
rect -1016 2343 -1004 2515
rect -970 2343 -958 2515
rect -1016 2129 -958 2343
rect -358 2515 -300 2729
rect -358 2343 -346 2515
rect -312 2343 -300 2515
rect -358 2129 -300 2343
rect 300 2515 358 2729
rect 300 2343 312 2515
rect 346 2343 358 2515
rect 300 2129 358 2343
rect 958 2515 1016 2729
rect 958 2343 970 2515
rect 1004 2343 1016 2515
rect 958 2129 1016 2343
rect -1016 1821 -958 2035
rect -1016 1649 -1004 1821
rect -970 1649 -958 1821
rect -1016 1435 -958 1649
rect -358 1821 -300 2035
rect -358 1649 -346 1821
rect -312 1649 -300 1821
rect -358 1435 -300 1649
rect 300 1821 358 2035
rect 300 1649 312 1821
rect 346 1649 358 1821
rect 300 1435 358 1649
rect 958 1821 1016 2035
rect 958 1649 970 1821
rect 1004 1649 1016 1821
rect 958 1435 1016 1649
rect -1016 1127 -958 1341
rect -1016 955 -1004 1127
rect -970 955 -958 1127
rect -1016 741 -958 955
rect -358 1127 -300 1341
rect -358 955 -346 1127
rect -312 955 -300 1127
rect -358 741 -300 955
rect 300 1127 358 1341
rect 300 955 312 1127
rect 346 955 358 1127
rect 300 741 358 955
rect 958 1127 1016 1341
rect 958 955 970 1127
rect 1004 955 1016 1127
rect 958 741 1016 955
rect -1016 433 -958 647
rect -1016 261 -1004 433
rect -970 261 -958 433
rect -1016 47 -958 261
rect -358 433 -300 647
rect -358 261 -346 433
rect -312 261 -300 433
rect -358 47 -300 261
rect 300 433 358 647
rect 300 261 312 433
rect 346 261 358 433
rect 300 47 358 261
rect 958 433 1016 647
rect 958 261 970 433
rect 1004 261 1016 433
rect 958 47 1016 261
rect -1016 -261 -958 -47
rect -1016 -433 -1004 -261
rect -970 -433 -958 -261
rect -1016 -647 -958 -433
rect -358 -261 -300 -47
rect -358 -433 -346 -261
rect -312 -433 -300 -261
rect -358 -647 -300 -433
rect 300 -261 358 -47
rect 300 -433 312 -261
rect 346 -433 358 -261
rect 300 -647 358 -433
rect 958 -261 1016 -47
rect 958 -433 970 -261
rect 1004 -433 1016 -261
rect 958 -647 1016 -433
rect -1016 -955 -958 -741
rect -1016 -1127 -1004 -955
rect -970 -1127 -958 -955
rect -1016 -1341 -958 -1127
rect -358 -955 -300 -741
rect -358 -1127 -346 -955
rect -312 -1127 -300 -955
rect -358 -1341 -300 -1127
rect 300 -955 358 -741
rect 300 -1127 312 -955
rect 346 -1127 358 -955
rect 300 -1341 358 -1127
rect 958 -955 1016 -741
rect 958 -1127 970 -955
rect 1004 -1127 1016 -955
rect 958 -1341 1016 -1127
rect -1016 -1649 -958 -1435
rect -1016 -1821 -1004 -1649
rect -970 -1821 -958 -1649
rect -1016 -2035 -958 -1821
rect -358 -1649 -300 -1435
rect -358 -1821 -346 -1649
rect -312 -1821 -300 -1649
rect -358 -2035 -300 -1821
rect 300 -1649 358 -1435
rect 300 -1821 312 -1649
rect 346 -1821 358 -1649
rect 300 -2035 358 -1821
rect 958 -1649 1016 -1435
rect 958 -1821 970 -1649
rect 1004 -1821 1016 -1649
rect 958 -2035 1016 -1821
rect -1016 -2343 -958 -2129
rect -1016 -2515 -1004 -2343
rect -970 -2515 -958 -2343
rect -1016 -2729 -958 -2515
rect -358 -2343 -300 -2129
rect -358 -2515 -346 -2343
rect -312 -2515 -300 -2343
rect -358 -2729 -300 -2515
rect 300 -2343 358 -2129
rect 300 -2515 312 -2343
rect 346 -2515 358 -2343
rect 300 -2729 358 -2515
rect 958 -2343 1016 -2129
rect 958 -2515 970 -2343
rect 1004 -2515 1016 -2343
rect 958 -2729 1016 -2515
rect -1016 -3037 -958 -2823
rect -1016 -3209 -1004 -3037
rect -970 -3209 -958 -3037
rect -1016 -3423 -958 -3209
rect -358 -3037 -300 -2823
rect -358 -3209 -346 -3037
rect -312 -3209 -300 -3037
rect -358 -3423 -300 -3209
rect 300 -3037 358 -2823
rect 300 -3209 312 -3037
rect 346 -3209 358 -3037
rect 300 -3423 358 -3209
rect 958 -3037 1016 -2823
rect 958 -3209 970 -3037
rect 1004 -3209 1016 -3037
rect 958 -3423 1016 -3209
<< mvndiffc >>
rect -1004 3037 -970 3209
rect -346 3037 -312 3209
rect 312 3037 346 3209
rect 970 3037 1004 3209
rect -1004 2343 -970 2515
rect -346 2343 -312 2515
rect 312 2343 346 2515
rect 970 2343 1004 2515
rect -1004 1649 -970 1821
rect -346 1649 -312 1821
rect 312 1649 346 1821
rect 970 1649 1004 1821
rect -1004 955 -970 1127
rect -346 955 -312 1127
rect 312 955 346 1127
rect 970 955 1004 1127
rect -1004 261 -970 433
rect -346 261 -312 433
rect 312 261 346 433
rect 970 261 1004 433
rect -1004 -433 -970 -261
rect -346 -433 -312 -261
rect 312 -433 346 -261
rect 970 -433 1004 -261
rect -1004 -1127 -970 -955
rect -346 -1127 -312 -955
rect 312 -1127 346 -955
rect 970 -1127 1004 -955
rect -1004 -1821 -970 -1649
rect -346 -1821 -312 -1649
rect 312 -1821 346 -1649
rect 970 -1821 1004 -1649
rect -1004 -2515 -970 -2343
rect -346 -2515 -312 -2343
rect 312 -2515 346 -2343
rect 970 -2515 1004 -2343
rect -1004 -3209 -970 -3037
rect -346 -3209 -312 -3037
rect 312 -3209 346 -3037
rect 970 -3209 1004 -3037
<< poly >>
rect -958 3423 -358 3449
rect -300 3423 300 3449
rect 358 3423 958 3449
rect -958 2797 -358 2823
rect -300 2797 300 2823
rect 358 2797 958 2823
rect -958 2729 -358 2755
rect -300 2729 300 2755
rect 358 2729 958 2755
rect -958 2103 -358 2129
rect -300 2103 300 2129
rect 358 2103 958 2129
rect -958 2035 -358 2061
rect -300 2035 300 2061
rect 358 2035 958 2061
rect -958 1409 -358 1435
rect -300 1409 300 1435
rect 358 1409 958 1435
rect -958 1341 -358 1367
rect -300 1341 300 1367
rect 358 1341 958 1367
rect -958 715 -358 741
rect -300 715 300 741
rect 358 715 958 741
rect -958 647 -358 673
rect -300 647 300 673
rect 358 647 958 673
rect -958 21 -358 47
rect -300 21 300 47
rect 358 21 958 47
rect -958 -47 -358 -21
rect -300 -47 300 -21
rect 358 -47 958 -21
rect -958 -673 -358 -647
rect -300 -673 300 -647
rect 358 -673 958 -647
rect -958 -741 -358 -715
rect -300 -741 300 -715
rect 358 -741 958 -715
rect -958 -1367 -358 -1341
rect -300 -1367 300 -1341
rect 358 -1367 958 -1341
rect -958 -1435 -358 -1409
rect -300 -1435 300 -1409
rect 358 -1435 958 -1409
rect -958 -2061 -358 -2035
rect -300 -2061 300 -2035
rect 358 -2061 958 -2035
rect -958 -2129 -358 -2103
rect -300 -2129 300 -2103
rect 358 -2129 958 -2103
rect -958 -2755 -358 -2729
rect -300 -2755 300 -2729
rect 358 -2755 958 -2729
rect -958 -2823 -358 -2797
rect -300 -2823 300 -2797
rect 358 -2823 958 -2797
rect -958 -3449 -358 -3423
rect -300 -3449 300 -3423
rect 358 -3449 958 -3423
<< locali >>
rect -1004 3209 -970 3225
rect -1004 3021 -970 3037
rect -346 3209 -312 3225
rect -346 3021 -312 3037
rect 312 3209 346 3225
rect 312 3021 346 3037
rect 970 3209 1004 3225
rect 970 3021 1004 3037
rect -1004 2515 -970 2531
rect -1004 2327 -970 2343
rect -346 2515 -312 2531
rect -346 2327 -312 2343
rect 312 2515 346 2531
rect 312 2327 346 2343
rect 970 2515 1004 2531
rect 970 2327 1004 2343
rect -1004 1821 -970 1837
rect -1004 1633 -970 1649
rect -346 1821 -312 1837
rect -346 1633 -312 1649
rect 312 1821 346 1837
rect 312 1633 346 1649
rect 970 1821 1004 1837
rect 970 1633 1004 1649
rect -1004 1127 -970 1143
rect -1004 939 -970 955
rect -346 1127 -312 1143
rect -346 939 -312 955
rect 312 1127 346 1143
rect 312 939 346 955
rect 970 1127 1004 1143
rect 970 939 1004 955
rect -1004 433 -970 449
rect -1004 245 -970 261
rect -346 433 -312 449
rect -346 245 -312 261
rect 312 433 346 449
rect 312 245 346 261
rect 970 433 1004 449
rect 970 245 1004 261
rect -1004 -261 -970 -245
rect -1004 -449 -970 -433
rect -346 -261 -312 -245
rect -346 -449 -312 -433
rect 312 -261 346 -245
rect 312 -449 346 -433
rect 970 -261 1004 -245
rect 970 -449 1004 -433
rect -1004 -955 -970 -939
rect -1004 -1143 -970 -1127
rect -346 -955 -312 -939
rect -346 -1143 -312 -1127
rect 312 -955 346 -939
rect 312 -1143 346 -1127
rect 970 -955 1004 -939
rect 970 -1143 1004 -1127
rect -1004 -1649 -970 -1633
rect -1004 -1837 -970 -1821
rect -346 -1649 -312 -1633
rect -346 -1837 -312 -1821
rect 312 -1649 346 -1633
rect 312 -1837 346 -1821
rect 970 -1649 1004 -1633
rect 970 -1837 1004 -1821
rect -1004 -2343 -970 -2327
rect -1004 -2531 -970 -2515
rect -346 -2343 -312 -2327
rect -346 -2531 -312 -2515
rect 312 -2343 346 -2327
rect 312 -2531 346 -2515
rect 970 -2343 1004 -2327
rect 970 -2531 1004 -2515
rect -1004 -3037 -970 -3021
rect -1004 -3225 -970 -3209
rect -346 -3037 -312 -3021
rect -346 -3225 -312 -3209
rect 312 -3037 346 -3021
rect 312 -3225 346 -3209
rect 970 -3037 1004 -3021
rect 970 -3225 1004 -3209
<< viali >>
rect -1004 3037 -970 3209
rect -346 3037 -312 3209
rect 312 3037 346 3209
rect 970 3037 1004 3209
rect -1004 2343 -970 2515
rect -346 2343 -312 2515
rect 312 2343 346 2515
rect 970 2343 1004 2515
rect -1004 1649 -970 1821
rect -346 1649 -312 1821
rect 312 1649 346 1821
rect 970 1649 1004 1821
rect -1004 955 -970 1127
rect -346 955 -312 1127
rect 312 955 346 1127
rect 970 955 1004 1127
rect -1004 261 -970 433
rect -346 261 -312 433
rect 312 261 346 433
rect 970 261 1004 433
rect -1004 -433 -970 -261
rect -346 -433 -312 -261
rect 312 -433 346 -261
rect 970 -433 1004 -261
rect -1004 -1127 -970 -955
rect -346 -1127 -312 -955
rect 312 -1127 346 -955
rect 970 -1127 1004 -955
rect -1004 -1821 -970 -1649
rect -346 -1821 -312 -1649
rect 312 -1821 346 -1649
rect 970 -1821 1004 -1649
rect -1004 -2515 -970 -2343
rect -346 -2515 -312 -2343
rect 312 -2515 346 -2343
rect 970 -2515 1004 -2343
rect -1004 -3209 -970 -3037
rect -346 -3209 -312 -3037
rect 312 -3209 346 -3037
rect 970 -3209 1004 -3037
<< metal1 >>
rect -1010 3209 -964 3221
rect -1010 3037 -1004 3209
rect -970 3037 -964 3209
rect -1010 3025 -964 3037
rect -352 3209 -306 3221
rect -352 3037 -346 3209
rect -312 3037 -306 3209
rect -352 3025 -306 3037
rect 306 3209 352 3221
rect 306 3037 312 3209
rect 346 3037 352 3209
rect 306 3025 352 3037
rect 964 3209 1010 3221
rect 964 3037 970 3209
rect 1004 3037 1010 3209
rect 964 3025 1010 3037
rect -1010 2515 -964 2527
rect -1010 2343 -1004 2515
rect -970 2343 -964 2515
rect -1010 2331 -964 2343
rect -352 2515 -306 2527
rect -352 2343 -346 2515
rect -312 2343 -306 2515
rect -352 2331 -306 2343
rect 306 2515 352 2527
rect 306 2343 312 2515
rect 346 2343 352 2515
rect 306 2331 352 2343
rect 964 2515 1010 2527
rect 964 2343 970 2515
rect 1004 2343 1010 2515
rect 964 2331 1010 2343
rect -1010 1821 -964 1833
rect -1010 1649 -1004 1821
rect -970 1649 -964 1821
rect -1010 1637 -964 1649
rect -352 1821 -306 1833
rect -352 1649 -346 1821
rect -312 1649 -306 1821
rect -352 1637 -306 1649
rect 306 1821 352 1833
rect 306 1649 312 1821
rect 346 1649 352 1821
rect 306 1637 352 1649
rect 964 1821 1010 1833
rect 964 1649 970 1821
rect 1004 1649 1010 1821
rect 964 1637 1010 1649
rect -1010 1127 -964 1139
rect -1010 955 -1004 1127
rect -970 955 -964 1127
rect -1010 943 -964 955
rect -352 1127 -306 1139
rect -352 955 -346 1127
rect -312 955 -306 1127
rect -352 943 -306 955
rect 306 1127 352 1139
rect 306 955 312 1127
rect 346 955 352 1127
rect 306 943 352 955
rect 964 1127 1010 1139
rect 964 955 970 1127
rect 1004 955 1010 1127
rect 964 943 1010 955
rect -1010 433 -964 445
rect -1010 261 -1004 433
rect -970 261 -964 433
rect -1010 249 -964 261
rect -352 433 -306 445
rect -352 261 -346 433
rect -312 261 -306 433
rect -352 249 -306 261
rect 306 433 352 445
rect 306 261 312 433
rect 346 261 352 433
rect 306 249 352 261
rect 964 433 1010 445
rect 964 261 970 433
rect 1004 261 1010 433
rect 964 249 1010 261
rect -1010 -261 -964 -249
rect -1010 -433 -1004 -261
rect -970 -433 -964 -261
rect -1010 -445 -964 -433
rect -352 -261 -306 -249
rect -352 -433 -346 -261
rect -312 -433 -306 -261
rect -352 -445 -306 -433
rect 306 -261 352 -249
rect 306 -433 312 -261
rect 346 -433 352 -261
rect 306 -445 352 -433
rect 964 -261 1010 -249
rect 964 -433 970 -261
rect 1004 -433 1010 -261
rect 964 -445 1010 -433
rect -1010 -955 -964 -943
rect -1010 -1127 -1004 -955
rect -970 -1127 -964 -955
rect -1010 -1139 -964 -1127
rect -352 -955 -306 -943
rect -352 -1127 -346 -955
rect -312 -1127 -306 -955
rect -352 -1139 -306 -1127
rect 306 -955 352 -943
rect 306 -1127 312 -955
rect 346 -1127 352 -955
rect 306 -1139 352 -1127
rect 964 -955 1010 -943
rect 964 -1127 970 -955
rect 1004 -1127 1010 -955
rect 964 -1139 1010 -1127
rect -1010 -1649 -964 -1637
rect -1010 -1821 -1004 -1649
rect -970 -1821 -964 -1649
rect -1010 -1833 -964 -1821
rect -352 -1649 -306 -1637
rect -352 -1821 -346 -1649
rect -312 -1821 -306 -1649
rect -352 -1833 -306 -1821
rect 306 -1649 352 -1637
rect 306 -1821 312 -1649
rect 346 -1821 352 -1649
rect 306 -1833 352 -1821
rect 964 -1649 1010 -1637
rect 964 -1821 970 -1649
rect 1004 -1821 1010 -1649
rect 964 -1833 1010 -1821
rect -1010 -2343 -964 -2331
rect -1010 -2515 -1004 -2343
rect -970 -2515 -964 -2343
rect -1010 -2527 -964 -2515
rect -352 -2343 -306 -2331
rect -352 -2515 -346 -2343
rect -312 -2515 -306 -2343
rect -352 -2527 -306 -2515
rect 306 -2343 352 -2331
rect 306 -2515 312 -2343
rect 346 -2515 352 -2343
rect 306 -2527 352 -2515
rect 964 -2343 1010 -2331
rect 964 -2515 970 -2343
rect 1004 -2515 1010 -2343
rect 964 -2527 1010 -2515
rect -1010 -3037 -964 -3025
rect -1010 -3209 -1004 -3037
rect -970 -3209 -964 -3037
rect -1010 -3221 -964 -3209
rect -352 -3037 -306 -3025
rect -352 -3209 -346 -3037
rect -312 -3209 -306 -3037
rect -352 -3221 -306 -3209
rect 306 -3037 352 -3025
rect 306 -3209 312 -3037
rect 346 -3209 352 -3037
rect 306 -3221 352 -3209
rect 964 -3037 1010 -3025
rect 964 -3209 970 -3037
rect 1004 -3209 1010 -3037
rect 964 -3221 1010 -3209
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string parameters w 3 l 3 m 10 nf 3 diffcov 30 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 30 viadrn 30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
