magic
tech sky130A
timestamp 1634050450
<< pwell >>
rect -19 15982 21179 16419
rect -191 -211 21200 15982
rect -191 -550 21211 -211
rect -11 -700 21211 -550
rect 169 -717 21211 -700
<< mvpsubdiff >>
rect -19 16389 21179 16419
rect -78 15994 21179 16389
rect -78 15941 21187 15994
rect -78 15620 430 15941
rect -78 15402 482 15620
rect -5 188 482 15402
rect 20580 14831 21187 15941
rect 20580 10876 20722 14831
rect 21064 10876 21187 14831
rect 20580 9035 21187 10876
rect 20580 5340 20670 9035
rect 21012 5340 21187 9035
rect 20580 3975 21187 5340
rect 20580 695 20774 3975
rect 21042 695 21187 3975
rect -11 -211 503 188
rect 20580 -211 21187 695
rect -11 -700 21211 -211
rect 169 -717 21211 -700
<< mvpsubdiffcont >>
rect 20722 10876 21064 14831
rect 20670 5340 21012 9035
rect 20774 695 21042 3975
<< poly >>
rect 10848 15511 11250 15648
<< polycont >>
rect 3888 15504 4002 15531
rect 18115 15501 18239 15534
<< locali >>
rect 3872 15531 4011 15541
rect 3872 15504 3888 15531
rect 4002 15504 4011 15531
rect 3872 15493 4011 15504
rect 18091 15534 18266 15540
rect 18091 15501 18115 15534
rect 18239 15501 18266 15534
rect 3912 15183 3961 15493
rect 18091 15488 18266 15501
rect 5433 15093 6629 15221
rect 7323 15051 7553 15289
rect 13578 14989 13808 15203
rect 18136 15153 18204 15488
rect 19290 15095 20548 15234
rect 20672 14831 21123 14897
rect 20672 10876 20722 14831
rect 21064 10876 21123 14831
rect 20672 10652 21123 10876
rect 20626 9035 21116 9139
rect 20626 5340 20670 9035
rect 21012 5340 21116 9035
rect 20626 5140 21116 5340
rect 20708 3975 21123 4101
rect 20708 695 20774 3975
rect 21042 695 21123 3975
rect 20708 569 21123 695
<< viali >>
rect 3911 15511 3970 15529
rect 18140 15507 18210 15533
rect 20767 11091 21012 14667
rect 20715 5437 20938 8924
rect 20811 932 20997 3901
<< metal1 >>
rect 3872 15529 4011 15541
rect 3872 15511 3911 15529
rect 3970 15511 4011 15529
rect 3872 15493 4011 15511
rect 18091 15533 18266 15540
rect 18091 15507 18140 15533
rect 18210 15507 18266 15533
rect 18091 15488 18266 15507
rect 20672 14667 21123 14897
rect 20672 11091 20767 14667
rect 21012 11091 21123 14667
rect 20672 10652 21123 11091
rect 20626 8924 21116 9139
rect 20626 5437 20715 8924
rect 20938 5437 21116 8924
rect 20626 5140 21116 5437
rect 20708 3901 21123 4101
rect 20708 932 20811 3901
rect 20997 932 21123 3901
rect 20708 569 21123 932
use nmos1010514  nmos1010514_2
timestamp 1634049493
transform 1 0 14014 0 1 4294
box -89 -4296 6980 11300
use nmos1010514  nmos1010514_1
timestamp 1634049493
transform 1 0 7060 0 1 4287
box -89 -4296 6980 11300
use nmos1010514  nmos1010514_0
timestamp 1634049493
transform 1 0 89 0 1 4296
box -89 -4296 6980 11300
<< labels >>
flabel locali 7382 15160 7382 15160 0 FreeSans 800 0 0 0 d
flabel locali 13691 15086 13691 15086 0 FreeSans 800 0 0 0 s
flabel poly 11024 15589 11024 15589 0 FreeSans 800 0 0 0 g
<< end >>
