magic
tech sky130A
timestamp 1634123280
<< nwell >>
rect 8751 10312 8881 10359
rect 125 80 9621 266
<< mvnsubdiff >>
rect 122 10407 9620 10518
rect 125 10270 315 10407
rect 133 266 311 10270
rect 9438 10206 9620 10407
rect 9438 9697 9489 10206
rect 9567 9697 9620 10206
rect 9438 9153 9620 9697
rect 9438 8493 9474 9153
rect 9547 8493 9620 9153
rect 9438 7783 9620 8493
rect 9438 7078 9485 7783
rect 9565 7078 9620 7783
rect 9438 5258 9620 7078
rect 9438 4528 9476 5258
rect 9556 4528 9620 5258
rect 9438 2161 9620 4528
rect 9438 1265 9493 2161
rect 9558 1265 9620 2161
rect 9438 266 9620 1265
rect 125 80 9621 266
<< mvnsubdiffcont >>
rect 9489 9697 9567 10206
rect 9474 8493 9547 9153
rect 9485 7078 9565 7783
rect 9476 4528 9556 5258
rect 9493 1265 9558 2161
<< poly >>
rect 1082 10368 1196 10382
rect 1082 10348 1114 10368
rect 582 10326 1114 10348
rect 1151 10348 1196 10368
rect 1151 10326 2941 10348
rect 8751 10344 8881 10359
rect 582 10305 2941 10326
rect 3638 10289 5997 10332
rect 8751 10325 8807 10344
rect 6830 10308 8807 10325
rect 8833 10325 8881 10344
rect 8833 10308 9271 10325
rect 6830 10291 9271 10308
<< polycont >>
rect 1114 10326 1151 10368
rect 8807 10308 8833 10344
<< locali >>
rect 1106 10368 1162 10374
rect 1106 10326 1114 10368
rect 1151 10326 1162 10368
rect 1106 10315 1162 10326
rect 209 10169 405 10230
rect 695 10167 720 10292
rect 1118 10222 1143 10315
rect 3486 10184 3560 10389
rect 8799 10344 8845 10352
rect 8799 10308 8807 10344
rect 8833 10308 8845 10344
rect 8799 10296 8845 10308
rect 8809 10230 8829 10296
rect 8985 10137 9019 10248
rect 9472 10206 9583 10231
rect 9472 10174 9489 10206
rect 9295 10109 9489 10174
rect 9472 9697 9489 10109
rect 9567 9697 9583 10206
rect 9472 9672 9583 9697
rect 3277 9089 3407 9309
rect 9461 9153 9575 9176
rect 9461 8493 9474 9153
rect 9547 8493 9575 9153
rect 9461 8450 9575 8493
rect 9470 7783 9584 7817
rect 9470 7078 9485 7783
rect 9565 7078 9584 7783
rect 9470 7051 9584 7078
rect 9463 5258 9577 5286
rect 9463 4528 9476 5258
rect 9556 4528 9577 5258
rect 9463 4488 9577 4528
rect 9478 2161 9573 2177
rect 9478 1265 9493 2161
rect 9558 1265 9573 2161
rect 9478 1199 9573 1265
<< viali >>
rect 1122 10335 1141 10360
rect 8814 10314 8831 10340
rect 9496 9760 9550 10182
rect 9481 8528 9532 9133
rect 9498 7165 9556 7705
rect 9481 4578 9545 5226
rect 9511 1334 9549 2118
<< metal1 >>
rect 1106 10360 1162 10374
rect 1106 10335 1122 10360
rect 1141 10335 1162 10360
rect 1106 10315 1162 10335
rect 8799 10340 8845 10352
rect 8799 10314 8814 10340
rect 8831 10314 8845 10340
rect 8799 10296 8845 10314
rect 9472 10182 9583 10231
rect 9472 9760 9496 10182
rect 9550 9760 9583 10182
rect 9472 9672 9583 9760
rect 5790 9327 6315 9402
rect 9461 9133 9575 9176
rect 9461 8528 9481 9133
rect 9532 8528 9575 9133
rect 9461 8450 9575 8528
rect 9470 7705 9584 7817
rect 9470 7165 9498 7705
rect 9556 7165 9584 7705
rect 9470 7051 9584 7165
rect 9463 5226 9577 5286
rect 9463 4578 9481 5226
rect 9545 4578 9577 5226
rect 9463 4488 9577 4578
rect 9478 2118 9573 2177
rect 9478 1334 9511 2118
rect 9549 1334 9573 2118
rect 9478 1199 9573 1334
use pmos33823  pmos33823_0 ~/layout test
timestamp 1634123280
transform 1 0 137 0 1 172
box -137 -172 3296 10404
use pmos33823  pmos33823_1
timestamp 1634123280
transform 1 0 3271 0 1 158
box -137 -172 3296 10404
use pmos33823  pmos33823_2
timestamp 1634123280
transform 1 0 6454 0 1 158
box -137 -172 3296 10404
<< labels >>
flabel locali 3517 10326 3517 10326 0 FreeSans 800 0 0 0 d
flabel locali 3296 9250 3296 9250 0 FreeSans 800 0 0 0 sub
flabel poly 5420 10314 5420 10314 0 FreeSans 800 0 0 0 g
flabel metal1 6236 9354 6236 9354 0 FreeSans 800 0 0 0 s
<< end >>
