magic
tech sky130A
timestamp 1634552665
<< pwell >>
rect -410 -462 6891 12086
<< poly >>
rect 4000 11772 4102 11774
rect 4000 11770 4111 11772
rect 2086 11663 4111 11770
rect 2090 11566 2347 11663
rect 4000 11559 4111 11663
rect 676 8640 826 8853
rect 1107 8643 1257 8856
rect 1661 8641 1811 8854
rect 2138 8638 2288 8851
rect 2622 8639 2772 8852
rect 3884 8654 4018 8850
rect 4310 8654 4444 8850
rect 4920 8657 5054 8853
rect 5394 8656 5528 8852
rect 5858 8658 5992 8854
rect 682 5715 836 5935
rect 1041 5714 1195 5934
rect 1720 5712 1874 5932
rect 2086 5717 2240 5937
rect 2638 5714 2792 5934
rect 3892 5724 4037 5942
rect 4308 5717 4461 5940
rect 4829 5718 4982 5941
rect 5382 5715 5535 5938
rect 5920 5716 6073 5939
rect 656 2787 810 3007
rect 1075 2788 1229 3008
rect 1610 2787 1764 3007
rect 2134 2783 2288 3003
rect 2745 2783 2899 3003
rect 3890 2781 4043 3004
rect 4373 2778 4526 3001
rect 4805 2781 4958 3004
rect 5386 2782 5539 3005
rect 5908 2780 6061 3003
<< locali >>
rect 2476 11441 3785 11518
rect 3032 152 4193 207
<< metal1 >>
rect 363 8366 413 9092
rect 3010 8382 3060 9108
rect 3604 8393 3654 9119
rect 6234 8404 6300 9152
rect 363 5433 413 6159
rect 3010 5466 3060 6192
rect 3582 5450 3632 6176
rect 6223 5428 6289 6176
rect 369 2506 419 3232
rect 3004 2523 3054 3249
rect 3598 2534 3648 3260
rect 6239 2550 6305 3298
use nmos5555  nmos5555_7
timestamp 1634301196
transform 1 0 3604 0 1 8845
box -376 -69 2845 2828
use nmos5555  nmos5555_6
timestamp 1634301196
transform 1 0 3608 0 1 5933
box -376 -69 2845 2828
use nmos5555  nmos5555_5
timestamp 1634301196
transform 1 0 3610 0 1 2997
box -376 -69 2845 2828
use nmos5555  nmos5555_4
timestamp 1634301196
transform 1 0 3612 0 1 68
box -376 -69 2845 2828
use nmos5555  nmos5555_3
timestamp 1634301196
transform 1 0 373 0 1 8846
box -376 -69 2845 2828
use nmos5555  nmos5555_2
timestamp 1634301196
transform 1 0 376 0 1 5927
box -376 -69 2845 2828
use nmos5555  nmos5555_1
timestamp 1634301196
transform 1 0 376 0 1 2998
box -376 -69 2845 2828
use nmos5555  nmos5555_0
timestamp 1634301196
transform 1 0 376 0 1 69
box -376 -69 2845 2828
<< end >>
