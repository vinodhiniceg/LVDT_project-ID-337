magic
tech sky130A
magscale 1 2
timestamp 1634046683
<< mvnmos >>
rect -2029 2141 -29 4141
rect 29 2141 2029 4141
rect -2029 47 -29 2047
rect 29 47 2029 2047
rect -2029 -2047 -29 -47
rect 29 -2047 2029 -47
rect -2029 -4141 -29 -2141
rect 29 -4141 2029 -2141
<< mvndiff >>
rect -2087 3437 -2029 4141
rect -2087 2845 -2075 3437
rect -2041 2845 -2029 3437
rect -2087 2141 -2029 2845
rect -29 3437 29 4141
rect -29 2845 -17 3437
rect 17 2845 29 3437
rect -29 2141 29 2845
rect 2029 3437 2087 4141
rect 2029 2845 2041 3437
rect 2075 2845 2087 3437
rect 2029 2141 2087 2845
rect -2087 1343 -2029 2047
rect -2087 751 -2075 1343
rect -2041 751 -2029 1343
rect -2087 47 -2029 751
rect -29 1343 29 2047
rect -29 751 -17 1343
rect 17 751 29 1343
rect -29 47 29 751
rect 2029 1343 2087 2047
rect 2029 751 2041 1343
rect 2075 751 2087 1343
rect 2029 47 2087 751
rect -2087 -751 -2029 -47
rect -2087 -1343 -2075 -751
rect -2041 -1343 -2029 -751
rect -2087 -2047 -2029 -1343
rect -29 -751 29 -47
rect -29 -1343 -17 -751
rect 17 -1343 29 -751
rect -29 -2047 29 -1343
rect 2029 -751 2087 -47
rect 2029 -1343 2041 -751
rect 2075 -1343 2087 -751
rect 2029 -2047 2087 -1343
rect -2087 -2845 -2029 -2141
rect -2087 -3437 -2075 -2845
rect -2041 -3437 -2029 -2845
rect -2087 -4141 -2029 -3437
rect -29 -2845 29 -2141
rect -29 -3437 -17 -2845
rect 17 -3437 29 -2845
rect -29 -4141 29 -3437
rect 2029 -2845 2087 -2141
rect 2029 -3437 2041 -2845
rect 2075 -3437 2087 -2845
rect 2029 -4141 2087 -3437
<< mvndiffc >>
rect -2075 2845 -2041 3437
rect -17 2845 17 3437
rect 2041 2845 2075 3437
rect -2075 751 -2041 1343
rect -17 751 17 1343
rect 2041 751 2075 1343
rect -2075 -1343 -2041 -751
rect -17 -1343 17 -751
rect 2041 -1343 2075 -751
rect -2075 -3437 -2041 -2845
rect -17 -3437 17 -2845
rect 2041 -3437 2075 -2845
<< poly >>
rect -2029 4141 -29 4167
rect 29 4141 2029 4167
rect -2029 2115 -29 2141
rect 29 2115 2029 2141
rect -2029 2047 -29 2073
rect 29 2047 2029 2073
rect -2029 21 -29 47
rect 29 21 2029 47
rect -2029 -47 -29 -21
rect 29 -47 2029 -21
rect -2029 -2073 -29 -2047
rect 29 -2073 2029 -2047
rect -2029 -2141 -29 -2115
rect 29 -2141 2029 -2115
rect -2029 -4167 -29 -4141
rect 29 -4167 2029 -4141
<< locali >>
rect -2075 3437 -2041 3453
rect -2075 2829 -2041 2845
rect -17 3437 17 3453
rect -17 2829 17 2845
rect 2041 3437 2075 3453
rect 2041 2829 2075 2845
rect -2075 1343 -2041 1359
rect -2075 735 -2041 751
rect -17 1343 17 1359
rect -17 735 17 751
rect 2041 1343 2075 1359
rect 2041 735 2075 751
rect -2075 -751 -2041 -735
rect -2075 -1359 -2041 -1343
rect -17 -751 17 -735
rect -17 -1359 17 -1343
rect 2041 -751 2075 -735
rect 2041 -1359 2075 -1343
rect -2075 -2845 -2041 -2829
rect -2075 -3453 -2041 -3437
rect -17 -2845 17 -2829
rect -17 -3453 17 -3437
rect 2041 -2845 2075 -2829
rect 2041 -3453 2075 -3437
<< viali >>
rect -2075 2845 -2041 3437
rect -17 2845 17 3437
rect 2041 2845 2075 3437
rect -2075 751 -2041 1343
rect -17 751 17 1343
rect 2041 751 2075 1343
rect -2075 -1343 -2041 -751
rect -17 -1343 17 -751
rect 2041 -1343 2075 -751
rect -2075 -3437 -2041 -2845
rect -17 -3437 17 -2845
rect 2041 -3437 2075 -2845
<< metal1 >>
rect -2081 3437 -2035 3449
rect -2081 2845 -2075 3437
rect -2041 2845 -2035 3437
rect -2081 2833 -2035 2845
rect -23 3437 23 3449
rect -23 2845 -17 3437
rect 17 2845 23 3437
rect -23 2833 23 2845
rect 2035 3437 2081 3449
rect 2035 2845 2041 3437
rect 2075 2845 2081 3437
rect 2035 2833 2081 2845
rect -2081 1343 -2035 1355
rect -2081 751 -2075 1343
rect -2041 751 -2035 1343
rect -2081 739 -2035 751
rect -23 1343 23 1355
rect -23 751 -17 1343
rect 17 751 23 1343
rect -23 739 23 751
rect 2035 1343 2081 1355
rect 2035 751 2041 1343
rect 2075 751 2081 1343
rect 2035 739 2081 751
rect -2081 -751 -2035 -739
rect -2081 -1343 -2075 -751
rect -2041 -1343 -2035 -751
rect -2081 -1355 -2035 -1343
rect -23 -751 23 -739
rect -23 -1343 -17 -751
rect 17 -1343 23 -751
rect -23 -1355 23 -1343
rect 2035 -751 2081 -739
rect 2035 -1343 2041 -751
rect 2075 -1343 2081 -751
rect 2035 -1355 2081 -1343
rect -2081 -2845 -2035 -2833
rect -2081 -3437 -2075 -2845
rect -2041 -3437 -2035 -2845
rect -2081 -3449 -2035 -3437
rect -23 -2845 23 -2833
rect -23 -3437 -17 -2845
rect 17 -3437 23 -2845
rect -23 -3449 23 -3437
rect 2035 -2845 2081 -2833
rect 2035 -3437 2041 -2845
rect 2075 -3437 2081 -2845
rect 2035 -3449 2081 -3437
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string parameters w 10 l 10 m 4 nf 2 diffcov 30 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 30 viadrn 30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
