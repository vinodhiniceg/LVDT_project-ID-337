magic
tech sky130A
timestamp 1634301196
<< error_s >>
rect 1587 2201 1616 2701
rect 2116 2201 2145 2701
rect 2645 2201 2674 2701
rect 1587 1654 1616 2154
rect 2116 1654 2145 2154
rect 2645 1654 2674 2154
rect 1587 1107 1616 1607
rect 2116 1107 2145 1607
rect 2645 1107 2674 1607
rect 1587 560 1616 1060
rect 2116 560 2145 1060
rect 2645 560 2674 1060
rect 1587 13 1616 513
rect 2116 13 2145 513
rect 2645 13 2674 513
<< pwell >>
rect -376 -69 2845 2828
<< mvpsubdiff >>
rect -333 1757 -229 1838
rect -333 1159 -310 1757
rect -263 1159 -229 1757
rect -333 977 -229 1159
<< mvpsubdiffcont >>
rect -310 1159 -263 1757
<< poly >>
rect 254 2711 2567 2735
rect 155 2164 422 2196
rect 674 2163 941 2195
rect 1233 2162 1500 2194
rect 1741 2160 2008 2192
rect 2274 2162 2541 2194
rect 173 1614 440 1646
rect 651 1615 918 1647
rect 1205 1614 1472 1646
rect 1758 1614 2025 1646
rect 2273 1614 2540 1646
rect 141 1068 408 1100
rect 668 1067 935 1099
rect 1194 1066 1461 1098
rect 1748 1067 2015 1099
rect 2276 1070 2543 1102
rect 155 522 422 554
rect 704 521 971 553
rect 1218 522 1485 554
rect 1700 521 1967 553
rect 2250 522 2517 554
<< locali >>
rect -1 2663 33 2668
rect 1051 2663 1085 2671
rect 2113 2663 2147 2679
rect -1 2658 2147 2663
rect -70 2636 2147 2658
rect -70 2618 2151 2636
rect -70 2613 2075 2618
rect -1 2473 33 2613
rect 1051 2506 1085 2613
rect 1051 2480 1088 2506
rect -321 1757 -246 1820
rect -321 1159 -310 1757
rect -263 1159 -246 1757
rect -321 997 -246 1159
rect -1 307 22 2473
rect 533 296 556 2477
rect 1059 307 1082 2480
rect 1593 299 1616 2480
rect 2109 2478 2151 2618
rect 2119 321 2142 2478
rect 2647 307 2670 2488
rect 525 135 566 240
rect 1588 135 1629 226
rect 2639 135 2680 237
rect 525 90 2750 135
rect 531 87 2750 90
rect 1588 76 1629 87
<< viali >>
rect -310 1159 -263 1757
<< metal1 >>
rect -321 1757 -246 1820
rect -321 1159 -310 1757
rect -263 1159 -246 1757
rect -321 997 -246 1159
use sky130_fd_pr__nfet_g5v0d10v5_7MG9ZH  sky130_fd_pr__nfet_g5v0d10v5_7MG9ZH_0
timestamp 1634301196
transform 1 0 1337 0 1 1357
box -1337 -1357 1337 1357
<< labels >>
flabel locali 2706 104 2706 104 0 FreeSans 800 0 0 0 d
flabel locali -45 2630 -45 2630 0 FreeSans 800 0 0 0 s
flabel poly 2061 2725 2061 2725 0 FreeSans 800 0 0 0 g
<< end >>
