magic
tech sky130A
magscale 1 2
timestamp 1634272161
<< error_p >>
rect -1411 1750 1411 1754
rect -1411 -1750 -1381 1750
rect -1345 1684 1345 1688
rect -1345 1088 -1315 1684
rect 1315 1088 1345 1684
rect -1345 394 -1315 994
rect 1315 394 1345 994
rect -1345 -300 -1315 300
rect 1315 -300 1345 300
rect -1345 -994 -1315 -394
rect 1315 -994 1345 -394
rect -1345 -1684 -1315 -1088
rect 1315 -1684 1345 -1088
rect -1345 -1688 1345 -1684
rect 1381 -1750 1411 1750
rect -1411 -1754 1411 -1750
<< nwell >>
rect -1381 -1750 1381 1750
<< mvpmos >>
rect -1287 1088 -687 1688
rect -629 1088 -29 1688
rect 29 1088 629 1688
rect 687 1088 1287 1688
rect -1287 394 -687 994
rect -629 394 -29 994
rect 29 394 629 994
rect 687 394 1287 994
rect -1287 -300 -687 300
rect -629 -300 -29 300
rect 29 -300 629 300
rect 687 -300 1287 300
rect -1287 -994 -687 -394
rect -629 -994 -29 -394
rect 29 -994 629 -394
rect 687 -994 1287 -394
rect -1287 -1688 -687 -1088
rect -629 -1688 -29 -1088
rect 29 -1688 629 -1088
rect 687 -1688 1287 -1088
<< mvpdiff >>
rect -1345 1474 -1287 1688
rect -1345 1302 -1333 1474
rect -1299 1302 -1287 1474
rect -1345 1088 -1287 1302
rect -687 1474 -629 1688
rect -687 1302 -675 1474
rect -641 1302 -629 1474
rect -687 1088 -629 1302
rect -29 1474 29 1688
rect -29 1302 -17 1474
rect 17 1302 29 1474
rect -29 1088 29 1302
rect 629 1474 687 1688
rect 629 1302 641 1474
rect 675 1302 687 1474
rect 629 1088 687 1302
rect 1287 1474 1345 1688
rect 1287 1302 1299 1474
rect 1333 1302 1345 1474
rect 1287 1088 1345 1302
rect -1345 780 -1287 994
rect -1345 608 -1333 780
rect -1299 608 -1287 780
rect -1345 394 -1287 608
rect -687 780 -629 994
rect -687 608 -675 780
rect -641 608 -629 780
rect -687 394 -629 608
rect -29 780 29 994
rect -29 608 -17 780
rect 17 608 29 780
rect -29 394 29 608
rect 629 780 687 994
rect 629 608 641 780
rect 675 608 687 780
rect 629 394 687 608
rect 1287 780 1345 994
rect 1287 608 1299 780
rect 1333 608 1345 780
rect 1287 394 1345 608
rect -1345 86 -1287 300
rect -1345 -86 -1333 86
rect -1299 -86 -1287 86
rect -1345 -300 -1287 -86
rect -687 86 -629 300
rect -687 -86 -675 86
rect -641 -86 -629 86
rect -687 -300 -629 -86
rect -29 86 29 300
rect -29 -86 -17 86
rect 17 -86 29 86
rect -29 -300 29 -86
rect 629 86 687 300
rect 629 -86 641 86
rect 675 -86 687 86
rect 629 -300 687 -86
rect 1287 86 1345 300
rect 1287 -86 1299 86
rect 1333 -86 1345 86
rect 1287 -300 1345 -86
rect -1345 -608 -1287 -394
rect -1345 -780 -1333 -608
rect -1299 -780 -1287 -608
rect -1345 -994 -1287 -780
rect -687 -608 -629 -394
rect -687 -780 -675 -608
rect -641 -780 -629 -608
rect -687 -994 -629 -780
rect -29 -608 29 -394
rect -29 -780 -17 -608
rect 17 -780 29 -608
rect -29 -994 29 -780
rect 629 -608 687 -394
rect 629 -780 641 -608
rect 675 -780 687 -608
rect 629 -994 687 -780
rect 1287 -608 1345 -394
rect 1287 -780 1299 -608
rect 1333 -780 1345 -608
rect 1287 -994 1345 -780
rect -1345 -1302 -1287 -1088
rect -1345 -1474 -1333 -1302
rect -1299 -1474 -1287 -1302
rect -1345 -1688 -1287 -1474
rect -687 -1302 -629 -1088
rect -687 -1474 -675 -1302
rect -641 -1474 -629 -1302
rect -687 -1688 -629 -1474
rect -29 -1302 29 -1088
rect -29 -1474 -17 -1302
rect 17 -1474 29 -1302
rect -29 -1688 29 -1474
rect 629 -1302 687 -1088
rect 629 -1474 641 -1302
rect 675 -1474 687 -1302
rect 629 -1688 687 -1474
rect 1287 -1302 1345 -1088
rect 1287 -1474 1299 -1302
rect 1333 -1474 1345 -1302
rect 1287 -1688 1345 -1474
<< mvpdiffc >>
rect -1333 1302 -1299 1474
rect -675 1302 -641 1474
rect -17 1302 17 1474
rect 641 1302 675 1474
rect 1299 1302 1333 1474
rect -1333 608 -1299 780
rect -675 608 -641 780
rect -17 608 17 780
rect 641 608 675 780
rect 1299 608 1333 780
rect -1333 -86 -1299 86
rect -675 -86 -641 86
rect -17 -86 17 86
rect 641 -86 675 86
rect 1299 -86 1333 86
rect -1333 -780 -1299 -608
rect -675 -780 -641 -608
rect -17 -780 17 -608
rect 641 -780 675 -608
rect 1299 -780 1333 -608
rect -1333 -1474 -1299 -1302
rect -675 -1474 -641 -1302
rect -17 -1474 17 -1302
rect 641 -1474 675 -1302
rect 1299 -1474 1333 -1302
<< poly >>
rect -1287 1688 -687 1714
rect -629 1688 -29 1714
rect 29 1688 629 1714
rect 687 1688 1287 1714
rect -1287 1062 -687 1088
rect -629 1062 -29 1088
rect 29 1062 629 1088
rect 687 1062 1287 1088
rect -1287 994 -687 1020
rect -629 994 -29 1020
rect 29 994 629 1020
rect 687 994 1287 1020
rect -1287 368 -687 394
rect -629 368 -29 394
rect 29 368 629 394
rect 687 368 1287 394
rect -1287 300 -687 326
rect -629 300 -29 326
rect 29 300 629 326
rect 687 300 1287 326
rect -1287 -326 -687 -300
rect -629 -326 -29 -300
rect 29 -326 629 -300
rect 687 -326 1287 -300
rect -1287 -394 -687 -368
rect -629 -394 -29 -368
rect 29 -394 629 -368
rect 687 -394 1287 -368
rect -1287 -1020 -687 -994
rect -629 -1020 -29 -994
rect 29 -1020 629 -994
rect 687 -1020 1287 -994
rect -1287 -1088 -687 -1062
rect -629 -1088 -29 -1062
rect 29 -1088 629 -1062
rect 687 -1088 1287 -1062
rect -1287 -1714 -687 -1688
rect -629 -1714 -29 -1688
rect 29 -1714 629 -1688
rect 687 -1714 1287 -1688
<< locali >>
rect -1333 1474 -1299 1490
rect -1333 1286 -1299 1302
rect -675 1474 -641 1490
rect -675 1286 -641 1302
rect -17 1474 17 1490
rect -17 1286 17 1302
rect 641 1474 675 1490
rect 641 1286 675 1302
rect 1299 1474 1333 1490
rect 1299 1286 1333 1302
rect -1333 780 -1299 796
rect -1333 592 -1299 608
rect -675 780 -641 796
rect -675 592 -641 608
rect -17 780 17 796
rect -17 592 17 608
rect 641 780 675 796
rect 641 592 675 608
rect 1299 780 1333 796
rect 1299 592 1333 608
rect -1333 86 -1299 102
rect -1333 -102 -1299 -86
rect -675 86 -641 102
rect -675 -102 -641 -86
rect -17 86 17 102
rect -17 -102 17 -86
rect 641 86 675 102
rect 641 -102 675 -86
rect 1299 86 1333 102
rect 1299 -102 1333 -86
rect -1333 -608 -1299 -592
rect -1333 -796 -1299 -780
rect -675 -608 -641 -592
rect -675 -796 -641 -780
rect -17 -608 17 -592
rect -17 -796 17 -780
rect 641 -608 675 -592
rect 641 -796 675 -780
rect 1299 -608 1333 -592
rect 1299 -796 1333 -780
rect -1333 -1302 -1299 -1286
rect -1333 -1490 -1299 -1474
rect -675 -1302 -641 -1286
rect -675 -1490 -641 -1474
rect -17 -1302 17 -1286
rect -17 -1490 17 -1474
rect 641 -1302 675 -1286
rect 641 -1490 675 -1474
rect 1299 -1302 1333 -1286
rect 1299 -1490 1333 -1474
<< viali >>
rect -1333 1302 -1299 1474
rect -675 1302 -641 1474
rect -17 1302 17 1474
rect 641 1302 675 1474
rect 1299 1302 1333 1474
rect -1333 608 -1299 780
rect -675 608 -641 780
rect -17 608 17 780
rect 641 608 675 780
rect 1299 608 1333 780
rect -1333 -86 -1299 86
rect -675 -86 -641 86
rect -17 -86 17 86
rect 641 -86 675 86
rect 1299 -86 1333 86
rect -1333 -780 -1299 -608
rect -675 -780 -641 -608
rect -17 -780 17 -608
rect 641 -780 675 -608
rect 1299 -780 1333 -608
rect -1333 -1474 -1299 -1302
rect -675 -1474 -641 -1302
rect -17 -1474 17 -1302
rect 641 -1474 675 -1302
rect 1299 -1474 1333 -1302
<< metal1 >>
rect -1339 1474 -1293 1486
rect -1339 1302 -1333 1474
rect -1299 1302 -1293 1474
rect -1339 1290 -1293 1302
rect -681 1474 -635 1486
rect -681 1302 -675 1474
rect -641 1302 -635 1474
rect -681 1290 -635 1302
rect -23 1474 23 1486
rect -23 1302 -17 1474
rect 17 1302 23 1474
rect -23 1290 23 1302
rect 635 1474 681 1486
rect 635 1302 641 1474
rect 675 1302 681 1474
rect 635 1290 681 1302
rect 1293 1474 1339 1486
rect 1293 1302 1299 1474
rect 1333 1302 1339 1474
rect 1293 1290 1339 1302
rect -1339 780 -1293 792
rect -1339 608 -1333 780
rect -1299 608 -1293 780
rect -1339 596 -1293 608
rect -681 780 -635 792
rect -681 608 -675 780
rect -641 608 -635 780
rect -681 596 -635 608
rect -23 780 23 792
rect -23 608 -17 780
rect 17 608 23 780
rect -23 596 23 608
rect 635 780 681 792
rect 635 608 641 780
rect 675 608 681 780
rect 635 596 681 608
rect 1293 780 1339 792
rect 1293 608 1299 780
rect 1333 608 1339 780
rect 1293 596 1339 608
rect -1339 86 -1293 98
rect -1339 -86 -1333 86
rect -1299 -86 -1293 86
rect -1339 -98 -1293 -86
rect -681 86 -635 98
rect -681 -86 -675 86
rect -641 -86 -635 86
rect -681 -98 -635 -86
rect -23 86 23 98
rect -23 -86 -17 86
rect 17 -86 23 86
rect -23 -98 23 -86
rect 635 86 681 98
rect 635 -86 641 86
rect 675 -86 681 86
rect 635 -98 681 -86
rect 1293 86 1339 98
rect 1293 -86 1299 86
rect 1333 -86 1339 86
rect 1293 -98 1339 -86
rect -1339 -608 -1293 -596
rect -1339 -780 -1333 -608
rect -1299 -780 -1293 -608
rect -1339 -792 -1293 -780
rect -681 -608 -635 -596
rect -681 -780 -675 -608
rect -641 -780 -635 -608
rect -681 -792 -635 -780
rect -23 -608 23 -596
rect -23 -780 -17 -608
rect 17 -780 23 -608
rect -23 -792 23 -780
rect 635 -608 681 -596
rect 635 -780 641 -608
rect 675 -780 681 -608
rect 635 -792 681 -780
rect 1293 -608 1339 -596
rect 1293 -780 1299 -608
rect 1333 -780 1339 -608
rect 1293 -792 1339 -780
rect -1339 -1302 -1293 -1290
rect -1339 -1474 -1333 -1302
rect -1299 -1474 -1293 -1302
rect -1339 -1486 -1293 -1474
rect -681 -1302 -635 -1290
rect -681 -1474 -675 -1302
rect -641 -1474 -635 -1302
rect -681 -1486 -635 -1474
rect -23 -1302 23 -1290
rect -23 -1474 -17 -1302
rect 17 -1474 23 -1302
rect -23 -1486 23 -1474
rect 635 -1302 681 -1290
rect 635 -1474 641 -1302
rect 675 -1474 681 -1302
rect 635 -1486 681 -1474
rect 1293 -1302 1339 -1290
rect 1293 -1474 1299 -1302
rect 1333 -1474 1339 -1302
rect 1293 -1486 1339 -1474
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string parameters w 3 l 3 m 5 nf 4 diffcov 30 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 30 viadrn 30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
