magic
tech sky130A
timestamp 1634178975
<< error_s >>
rect 1663 1419 1692 1719
rect 1663 1072 1692 1372
rect 1663 725 1692 1025
rect 1663 378 1692 678
rect 1663 31 1692 331
<< nwell >>
rect -281 -180 1875 1835
<< mvnsubdiff >>
rect -241 1585 -40 1620
rect -241 385 -228 1585
rect -62 385 -40 1585
rect -241 297 -40 385
<< mvnsubdiffcont >>
rect -228 385 -62 1585
<< poly >>
rect 170 1728 1503 1763
rect 90 1379 313 1412
rect 411 1374 631 1417
rect 778 1376 998 1419
rect 1070 1375 1290 1418
rect 1389 1375 1609 1418
rect 80 1029 300 1072
rect 417 1025 637 1068
rect 764 1023 984 1066
rect 1064 1026 1284 1069
rect 1402 1026 1622 1069
rect 87 680 307 723
rect 409 676 629 719
rect 753 679 973 722
rect 1064 680 1284 723
rect 1408 681 1628 724
rect 86 331 306 374
rect 421 332 641 375
rect 759 335 979 378
rect 1075 334 1295 377
rect 1429 334 1649 377
<< locali >>
rect 9 1696 47 1708
rect 673 1696 711 1726
rect 1330 1696 1368 1711
rect 9 1669 1369 1696
rect -246 1585 -45 1633
rect -246 385 -228 1585
rect -62 385 -45 1585
rect 9 1576 47 1669
rect -246 310 -45 385
rect 18 175 45 1576
rect 347 192 374 1617
rect 673 1594 711 1669
rect 676 199 703 1594
rect 1005 207 1032 1621
rect 1330 1579 1368 1669
rect 340 90 378 192
rect 1001 90 1039 207
rect 1337 198 1364 1579
rect 1664 197 1691 1618
rect 1654 188 1691 197
rect 1654 90 1692 188
rect 340 49 1693 90
rect 1001 47 1039 49
rect 1654 47 1692 49
<< viali >>
rect -202 459 -101 1546
<< metal1 >>
rect -246 1546 -45 1633
rect -246 459 -202 1546
rect -101 459 -45 1546
rect -246 310 -45 459
use sky130_fd_pr__pfet_g5v0d10v5_TA684Z  sky130_fd_pr__pfet_g5v0d10v5_TA684Z_0
timestamp 1634178975
transform 1 0 855 0 1 875
box -870 -877 870 877
<< end >>
