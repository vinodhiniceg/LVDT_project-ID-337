magic
tech sky130A
timestamp 1634226173
<< pwell >>
rect -47 2462 5313 2470
rect -99 2344 5313 2462
rect -99 2240 5320 2344
rect -87 -218 5320 2240
<< mvpsubdiff >>
rect -47 2277 5261 2470
rect -55 2248 5261 2277
rect -55 -10 189 2248
rect 4994 2092 5238 2248
rect 4994 130 5054 2092
rect 5172 130 5238 2092
rect 4994 42 5238 130
rect -55 -62 175 -10
rect 4972 -25 5238 42
rect 4972 -62 5231 -25
rect -55 -210 5231 -62
rect -10 -218 5231 -210
rect 4972 -232 5231 -218
<< mvpsubdiffcont >>
rect 5054 130 5172 2092
<< poly >>
rect 879 2205 1135 2221
rect 879 2153 951 2205
rect 1081 2153 1135 2205
rect 879 2136 1135 2153
rect 4160 2212 4423 2234
rect 4160 2156 4213 2212
rect 4341 2156 4423 2212
rect 4160 2136 4423 2156
<< polycont >>
rect 951 2153 1081 2205
rect 4213 2156 4341 2212
<< locali >>
rect 931 2205 1100 2214
rect 931 2153 951 2205
rect 1081 2153 1100 2205
rect 931 2143 1100 2153
rect 4197 2212 4369 2221
rect 4197 2156 4213 2212
rect 4341 2156 4369 2212
rect 4197 2151 4369 2156
rect 970 2047 1036 2143
rect 1233 1949 1299 2097
rect 4230 2043 4310 2151
rect 5031 2092 5187 2144
rect 4557 1958 4618 2080
rect 5031 1908 5054 2092
rect 4898 1872 5054 1908
rect 1580 1785 1784 1833
rect 5031 130 5054 1872
rect 5172 130 5187 2092
rect 5031 71 5187 130
<< viali >>
rect 968 2158 1070 2203
rect 4225 2160 4325 2208
rect 5076 278 5135 1944
<< metal1 >>
rect 931 2203 1100 2214
rect 931 2158 968 2203
rect 1070 2158 1100 2203
rect 931 2143 1100 2158
rect 4197 2208 4369 2221
rect 4197 2160 4225 2208
rect 4325 2160 4369 2208
rect 4197 2151 4369 2160
rect 5031 1944 5187 2144
rect 5031 278 5076 1944
rect 5135 278 5187 1944
rect 5031 71 5187 278
use nmos3346  nmos3346_1 ~/layout test
timestamp 1634225045
transform 1 0 1925 0 1 53
box -262 -56 1351 2101
use nmos3346  nmos3346_0
timestamp 1634225045
transform 1 0 262 0 1 56
box -262 -56 1351 2101
use nmos3346  nmos3346_2
timestamp 1634225045
transform 1 0 3580 0 1 53
box -262 -56 1351 2101
<< end >>
