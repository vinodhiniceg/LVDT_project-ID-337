magic
tech sky130A
magscale 1 2
timestamp 1634638746
<< nwell >>
rect -1430 -253 -1010 267
rect -352 -250 5832 960
rect 6548 -163 6968 357
rect 7386 -145 7806 375
rect 8206 -149 8626 371
rect -356 -444 5832 -250
rect -356 -1500 538 -444
rect 4940 -726 5832 -444
rect 4940 -1376 5854 -726
rect 4940 -1490 5832 -1376
<< pwell >>
rect -1360 -587 -1094 -347
rect -1390 -673 -1050 -587
rect 608 -1524 4866 -482
rect 6632 -497 6898 -257
rect 7470 -479 7736 -239
rect 6588 -583 6928 -497
rect 7426 -565 7766 -479
rect 8290 -483 8556 -243
rect 8246 -569 8586 -483
<< mvnmos >>
rect -1277 -523 -1177 -373
rect 6715 -433 6815 -283
rect 7553 -415 7653 -265
rect 8373 -419 8473 -269
rect 1688 -866 1788 -666
rect 1846 -866 1946 -666
rect 2004 -866 2104 -666
rect 2162 -866 2262 -666
rect 3206 -872 3306 -672
rect 3364 -872 3464 -672
rect 3522 -872 3622 -672
rect 3680 -872 3780 -672
rect 1688 -1160 1788 -960
rect 1846 -1160 1946 -960
rect 2004 -1160 2104 -960
rect 2162 -1160 2262 -960
rect 2454 -1170 2554 -970
rect 2612 -1170 2712 -970
rect 2770 -1170 2870 -970
rect 2928 -1170 3028 -970
rect 3206 -1166 3306 -966
rect 3364 -1166 3464 -966
rect 3522 -1166 3622 -966
rect 3680 -1166 3780 -966
rect 938 -1464 1038 -1264
rect 1096 -1464 1196 -1264
rect 1254 -1464 1354 -1264
rect 1412 -1464 1512 -1264
rect 1688 -1454 1788 -1254
rect 1846 -1454 1946 -1254
rect 2004 -1454 2104 -1254
rect 2162 -1454 2262 -1254
rect 2454 -1464 2554 -1264
rect 2612 -1464 2712 -1264
rect 2770 -1464 2870 -1264
rect 2928 -1464 3028 -1264
rect 3206 -1460 3306 -1260
rect 3364 -1460 3464 -1260
rect 3522 -1460 3622 -1260
rect 3680 -1460 3780 -1260
rect 3956 -1464 4056 -1264
rect 4114 -1464 4214 -1264
rect 4272 -1464 4372 -1264
rect 4430 -1464 4530 -1264
rect 7524 -1348 7624 -1148
rect 8334 -1338 8434 -1138
<< mvpmos >>
rect 134 380 234 580
rect 292 380 392 580
rect 450 380 550 580
rect 608 380 708 580
rect 1038 382 1138 582
rect 1196 382 1296 582
rect 1354 382 1454 582
rect 1512 382 1612 582
rect 1942 382 2042 582
rect 2100 382 2200 582
rect 2258 382 2358 582
rect 2416 382 2516 582
rect 2828 378 2928 578
rect 2986 378 3086 578
rect 3144 378 3244 578
rect 3302 378 3402 578
rect 3704 380 3804 580
rect 3862 380 3962 580
rect 4020 380 4120 580
rect 4178 380 4278 580
rect 4568 378 4668 578
rect 4726 378 4826 578
rect 4884 378 4984 578
rect 5042 378 5142 578
rect -1273 -187 -1173 113
rect 134 86 234 286
rect 292 86 392 286
rect 450 86 550 286
rect 608 86 708 286
rect 1038 88 1138 288
rect 1196 88 1296 288
rect 1354 88 1454 288
rect 1512 88 1612 288
rect 1942 88 2042 288
rect 2100 88 2200 288
rect 2258 88 2358 288
rect 2416 88 2516 288
rect 2828 84 2928 284
rect 2986 84 3086 284
rect 3144 84 3244 284
rect 3302 84 3402 284
rect 3704 86 3804 286
rect 3862 86 3962 286
rect 4020 86 4120 286
rect 4178 86 4278 286
rect 4568 84 4668 284
rect 4726 84 4826 284
rect 4884 84 4984 284
rect 5042 84 5142 284
rect 6711 -97 6811 203
rect 7549 -79 7649 221
rect 8369 -83 8469 217
rect -202 -1022 -102 -822
rect -44 -1022 56 -822
rect 114 -1022 214 -822
rect 272 -1022 372 -822
rect -202 -1316 -102 -1116
rect -44 -1316 56 -1116
rect 114 -1316 214 -1116
rect 272 -1316 372 -1116
rect 5154 -996 5254 -796
rect 5312 -996 5412 -796
rect 5470 -996 5570 -796
rect 5628 -996 5728 -796
rect 5154 -1290 5254 -1090
rect 5312 -1290 5412 -1090
rect 5470 -1290 5570 -1090
rect 5628 -1290 5728 -1090
<< mvndiff >>
rect 7496 -273 7553 -265
rect 6658 -291 6715 -283
rect 6658 -325 6670 -291
rect 6704 -325 6715 -291
rect -1334 -381 -1277 -373
rect -1334 -415 -1322 -381
rect -1288 -415 -1277 -381
rect -1334 -481 -1277 -415
rect -1334 -515 -1322 -481
rect -1288 -515 -1277 -481
rect -1334 -523 -1277 -515
rect -1177 -381 -1120 -373
rect -1177 -415 -1166 -381
rect -1132 -415 -1120 -381
rect -1177 -481 -1120 -415
rect 6658 -391 6715 -325
rect 6658 -425 6670 -391
rect 6704 -425 6715 -391
rect 6658 -433 6715 -425
rect 6815 -291 6872 -283
rect 6815 -325 6826 -291
rect 6860 -325 6872 -291
rect 6815 -391 6872 -325
rect 6815 -425 6826 -391
rect 6860 -425 6872 -391
rect 7496 -307 7508 -273
rect 7542 -307 7553 -273
rect 7496 -373 7553 -307
rect 7496 -407 7508 -373
rect 7542 -407 7553 -373
rect 7496 -415 7553 -407
rect 7653 -273 7710 -265
rect 7653 -307 7664 -273
rect 7698 -307 7710 -273
rect 7653 -373 7710 -307
rect 7653 -407 7664 -373
rect 7698 -407 7710 -373
rect 7653 -415 7710 -407
rect 8316 -277 8373 -269
rect 8316 -311 8328 -277
rect 8362 -311 8373 -277
rect 8316 -377 8373 -311
rect 8316 -411 8328 -377
rect 8362 -411 8373 -377
rect 6815 -433 6872 -425
rect 8316 -419 8373 -411
rect 8473 -277 8530 -269
rect 8473 -311 8484 -277
rect 8518 -311 8530 -277
rect 8473 -377 8530 -311
rect 8473 -411 8484 -377
rect 8518 -411 8530 -377
rect 8473 -419 8530 -411
rect -1177 -515 -1166 -481
rect -1132 -515 -1120 -481
rect -1177 -523 -1120 -515
rect 1630 -740 1688 -666
rect 1630 -792 1642 -740
rect 1676 -792 1688 -740
rect 1630 -866 1688 -792
rect 1788 -740 1846 -666
rect 1788 -792 1800 -740
rect 1834 -792 1846 -740
rect 1788 -866 1846 -792
rect 1946 -740 2004 -666
rect 1946 -792 1958 -740
rect 1992 -792 2004 -740
rect 1946 -866 2004 -792
rect 2104 -740 2162 -666
rect 2104 -792 2116 -740
rect 2150 -792 2162 -740
rect 2104 -866 2162 -792
rect 2262 -740 2320 -666
rect 2262 -792 2274 -740
rect 2308 -792 2320 -740
rect 2262 -866 2320 -792
rect 3148 -746 3206 -672
rect 3148 -798 3160 -746
rect 3194 -798 3206 -746
rect 3148 -872 3206 -798
rect 3306 -746 3364 -672
rect 3306 -798 3318 -746
rect 3352 -798 3364 -746
rect 3306 -872 3364 -798
rect 3464 -746 3522 -672
rect 3464 -798 3476 -746
rect 3510 -798 3522 -746
rect 3464 -872 3522 -798
rect 3622 -746 3680 -672
rect 3622 -798 3634 -746
rect 3668 -798 3680 -746
rect 3622 -872 3680 -798
rect 3780 -746 3838 -672
rect 3780 -798 3792 -746
rect 3826 -798 3838 -746
rect 3780 -872 3838 -798
rect 1630 -1034 1688 -960
rect 1630 -1086 1642 -1034
rect 1676 -1086 1688 -1034
rect 1630 -1160 1688 -1086
rect 1788 -1034 1846 -960
rect 1788 -1086 1800 -1034
rect 1834 -1086 1846 -1034
rect 1788 -1160 1846 -1086
rect 1946 -1034 2004 -960
rect 1946 -1086 1958 -1034
rect 1992 -1086 2004 -1034
rect 1946 -1160 2004 -1086
rect 2104 -1034 2162 -960
rect 2104 -1086 2116 -1034
rect 2150 -1086 2162 -1034
rect 2104 -1160 2162 -1086
rect 2262 -1034 2320 -960
rect 2262 -1086 2274 -1034
rect 2308 -1086 2320 -1034
rect 2262 -1160 2320 -1086
rect 2396 -1044 2454 -970
rect 2396 -1096 2408 -1044
rect 2442 -1096 2454 -1044
rect 2396 -1170 2454 -1096
rect 2554 -1044 2612 -970
rect 2554 -1096 2566 -1044
rect 2600 -1096 2612 -1044
rect 2554 -1170 2612 -1096
rect 2712 -1044 2770 -970
rect 2712 -1096 2724 -1044
rect 2758 -1096 2770 -1044
rect 2712 -1170 2770 -1096
rect 2870 -1044 2928 -970
rect 2870 -1096 2882 -1044
rect 2916 -1096 2928 -1044
rect 2870 -1170 2928 -1096
rect 3028 -1044 3086 -970
rect 3028 -1096 3040 -1044
rect 3074 -1096 3086 -1044
rect 3028 -1170 3086 -1096
rect 3148 -1040 3206 -966
rect 3148 -1092 3160 -1040
rect 3194 -1092 3206 -1040
rect 3148 -1166 3206 -1092
rect 3306 -1040 3364 -966
rect 3306 -1092 3318 -1040
rect 3352 -1092 3364 -1040
rect 3306 -1166 3364 -1092
rect 3464 -1040 3522 -966
rect 3464 -1092 3476 -1040
rect 3510 -1092 3522 -1040
rect 3464 -1166 3522 -1092
rect 3622 -1040 3680 -966
rect 3622 -1092 3634 -1040
rect 3668 -1092 3680 -1040
rect 3622 -1166 3680 -1092
rect 3780 -1040 3838 -966
rect 3780 -1092 3792 -1040
rect 3826 -1092 3838 -1040
rect 3780 -1166 3838 -1092
rect 880 -1338 938 -1264
rect 880 -1390 892 -1338
rect 926 -1390 938 -1338
rect 880 -1464 938 -1390
rect 1038 -1338 1096 -1264
rect 1038 -1390 1050 -1338
rect 1084 -1390 1096 -1338
rect 1038 -1464 1096 -1390
rect 1196 -1338 1254 -1264
rect 1196 -1390 1208 -1338
rect 1242 -1390 1254 -1338
rect 1196 -1464 1254 -1390
rect 1354 -1338 1412 -1264
rect 1354 -1390 1366 -1338
rect 1400 -1390 1412 -1338
rect 1354 -1464 1412 -1390
rect 1512 -1338 1570 -1264
rect 1512 -1390 1524 -1338
rect 1558 -1390 1570 -1338
rect 1512 -1464 1570 -1390
rect 1630 -1328 1688 -1254
rect 1630 -1380 1642 -1328
rect 1676 -1380 1688 -1328
rect 1630 -1454 1688 -1380
rect 1788 -1328 1846 -1254
rect 1788 -1380 1800 -1328
rect 1834 -1380 1846 -1328
rect 1788 -1454 1846 -1380
rect 1946 -1328 2004 -1254
rect 1946 -1380 1958 -1328
rect 1992 -1380 2004 -1328
rect 1946 -1454 2004 -1380
rect 2104 -1328 2162 -1254
rect 2104 -1380 2116 -1328
rect 2150 -1380 2162 -1328
rect 2104 -1454 2162 -1380
rect 2262 -1328 2320 -1254
rect 2262 -1380 2274 -1328
rect 2308 -1380 2320 -1328
rect 2262 -1454 2320 -1380
rect 2396 -1338 2454 -1264
rect 2396 -1390 2408 -1338
rect 2442 -1390 2454 -1338
rect 2396 -1464 2454 -1390
rect 2554 -1338 2612 -1264
rect 2554 -1390 2566 -1338
rect 2600 -1390 2612 -1338
rect 2554 -1464 2612 -1390
rect 2712 -1338 2770 -1264
rect 2712 -1390 2724 -1338
rect 2758 -1390 2770 -1338
rect 2712 -1464 2770 -1390
rect 2870 -1338 2928 -1264
rect 2870 -1390 2882 -1338
rect 2916 -1390 2928 -1338
rect 2870 -1464 2928 -1390
rect 3028 -1338 3086 -1264
rect 3028 -1390 3040 -1338
rect 3074 -1390 3086 -1338
rect 3028 -1464 3086 -1390
rect 3148 -1334 3206 -1260
rect 3148 -1386 3160 -1334
rect 3194 -1386 3206 -1334
rect 3148 -1460 3206 -1386
rect 3306 -1334 3364 -1260
rect 3306 -1386 3318 -1334
rect 3352 -1386 3364 -1334
rect 3306 -1460 3364 -1386
rect 3464 -1334 3522 -1260
rect 3464 -1386 3476 -1334
rect 3510 -1386 3522 -1334
rect 3464 -1460 3522 -1386
rect 3622 -1334 3680 -1260
rect 3622 -1386 3634 -1334
rect 3668 -1386 3680 -1334
rect 3622 -1460 3680 -1386
rect 3780 -1334 3838 -1260
rect 3780 -1386 3792 -1334
rect 3826 -1386 3838 -1334
rect 3780 -1460 3838 -1386
rect 3898 -1338 3956 -1264
rect 3898 -1390 3910 -1338
rect 3944 -1390 3956 -1338
rect 3898 -1464 3956 -1390
rect 4056 -1338 4114 -1264
rect 4056 -1390 4068 -1338
rect 4102 -1390 4114 -1338
rect 4056 -1464 4114 -1390
rect 4214 -1338 4272 -1264
rect 4214 -1390 4226 -1338
rect 4260 -1390 4272 -1338
rect 4214 -1464 4272 -1390
rect 4372 -1338 4430 -1264
rect 4372 -1390 4384 -1338
rect 4418 -1390 4430 -1338
rect 4372 -1464 4430 -1390
rect 4530 -1338 4588 -1264
rect 4530 -1390 4542 -1338
rect 4576 -1390 4588 -1338
rect 4530 -1464 4588 -1390
rect 7466 -1222 7524 -1148
rect 7466 -1274 7478 -1222
rect 7512 -1274 7524 -1222
rect 7466 -1348 7524 -1274
rect 7624 -1222 7682 -1148
rect 7624 -1274 7636 -1222
rect 7670 -1274 7682 -1222
rect 7624 -1348 7682 -1274
rect 8276 -1212 8334 -1138
rect 8276 -1264 8288 -1212
rect 8322 -1264 8334 -1212
rect 8276 -1338 8334 -1264
rect 8434 -1212 8492 -1138
rect 8434 -1264 8446 -1212
rect 8480 -1264 8492 -1212
rect 8434 -1338 8492 -1264
<< mvpdiff >>
rect 76 506 134 580
rect 76 454 88 506
rect 122 454 134 506
rect 76 380 134 454
rect 234 506 292 580
rect 234 454 246 506
rect 280 454 292 506
rect 234 380 292 454
rect 392 506 450 580
rect 392 454 404 506
rect 438 454 450 506
rect 392 380 450 454
rect 550 506 608 580
rect 550 454 562 506
rect 596 454 608 506
rect 550 380 608 454
rect 708 506 766 580
rect 708 454 720 506
rect 754 454 766 506
rect 708 380 766 454
rect 980 508 1038 582
rect 980 456 992 508
rect 1026 456 1038 508
rect 980 382 1038 456
rect 1138 508 1196 582
rect 1138 456 1150 508
rect 1184 456 1196 508
rect 1138 382 1196 456
rect 1296 508 1354 582
rect 1296 456 1308 508
rect 1342 456 1354 508
rect 1296 382 1354 456
rect 1454 508 1512 582
rect 1454 456 1466 508
rect 1500 456 1512 508
rect 1454 382 1512 456
rect 1612 508 1670 582
rect 1612 456 1624 508
rect 1658 456 1670 508
rect 1612 382 1670 456
rect 1884 508 1942 582
rect 1884 456 1896 508
rect 1930 456 1942 508
rect 1884 382 1942 456
rect 2042 508 2100 582
rect 2042 456 2054 508
rect 2088 456 2100 508
rect 2042 382 2100 456
rect 2200 508 2258 582
rect 2200 456 2212 508
rect 2246 456 2258 508
rect 2200 382 2258 456
rect 2358 508 2416 582
rect 2358 456 2370 508
rect 2404 456 2416 508
rect 2358 382 2416 456
rect 2516 508 2574 582
rect 2516 456 2528 508
rect 2562 456 2574 508
rect 2516 382 2574 456
rect 2770 504 2828 578
rect 2770 452 2782 504
rect 2816 452 2828 504
rect 2770 378 2828 452
rect 2928 504 2986 578
rect 2928 452 2940 504
rect 2974 452 2986 504
rect 2928 378 2986 452
rect 3086 504 3144 578
rect 3086 452 3098 504
rect 3132 452 3144 504
rect 3086 378 3144 452
rect 3244 504 3302 578
rect 3244 452 3256 504
rect 3290 452 3302 504
rect 3244 378 3302 452
rect 3402 504 3460 578
rect 3402 452 3414 504
rect 3448 452 3460 504
rect 3402 378 3460 452
rect 3646 506 3704 580
rect 3646 454 3658 506
rect 3692 454 3704 506
rect 3646 380 3704 454
rect 3804 506 3862 580
rect 3804 454 3816 506
rect 3850 454 3862 506
rect 3804 380 3862 454
rect 3962 506 4020 580
rect 3962 454 3974 506
rect 4008 454 4020 506
rect 3962 380 4020 454
rect 4120 506 4178 580
rect 4120 454 4132 506
rect 4166 454 4178 506
rect 4120 380 4178 454
rect 4278 506 4336 580
rect 4278 454 4290 506
rect 4324 454 4336 506
rect 4278 380 4336 454
rect 4510 504 4568 578
rect 4510 452 4522 504
rect 4556 452 4568 504
rect 4510 378 4568 452
rect 4668 504 4726 578
rect 4668 452 4680 504
rect 4714 452 4726 504
rect 4668 378 4726 452
rect 4826 504 4884 578
rect 4826 452 4838 504
rect 4872 452 4884 504
rect 4826 378 4884 452
rect 4984 504 5042 578
rect 4984 452 4996 504
rect 5030 452 5042 504
rect 4984 378 5042 452
rect 5142 504 5200 578
rect 5142 452 5154 504
rect 5188 452 5200 504
rect 5142 378 5200 452
rect -1330 105 -1273 113
rect -1330 71 -1318 105
rect -1284 71 -1273 105
rect -1330 22 -1273 71
rect -1330 -12 -1318 22
rect -1284 -12 -1273 22
rect -1330 -62 -1273 -12
rect -1330 -96 -1318 -62
rect -1284 -96 -1273 -62
rect -1330 -145 -1273 -96
rect -1330 -179 -1318 -145
rect -1284 -179 -1273 -145
rect -1330 -187 -1273 -179
rect -1173 105 -1116 113
rect -1173 71 -1162 105
rect -1128 71 -1116 105
rect -1173 22 -1116 71
rect 76 212 134 286
rect 76 160 88 212
rect 122 160 134 212
rect 76 86 134 160
rect 234 212 292 286
rect 234 160 246 212
rect 280 160 292 212
rect 234 86 292 160
rect 392 212 450 286
rect 392 160 404 212
rect 438 160 450 212
rect 392 86 450 160
rect 550 212 608 286
rect 550 160 562 212
rect 596 160 608 212
rect 550 86 608 160
rect 708 212 766 286
rect 708 160 720 212
rect 754 160 766 212
rect 708 86 766 160
rect 980 214 1038 288
rect 980 162 992 214
rect 1026 162 1038 214
rect 980 88 1038 162
rect 1138 214 1196 288
rect 1138 162 1150 214
rect 1184 162 1196 214
rect 1138 88 1196 162
rect 1296 214 1354 288
rect 1296 162 1308 214
rect 1342 162 1354 214
rect 1296 88 1354 162
rect 1454 214 1512 288
rect 1454 162 1466 214
rect 1500 162 1512 214
rect 1454 88 1512 162
rect 1612 214 1670 288
rect 1612 162 1624 214
rect 1658 162 1670 214
rect 1612 88 1670 162
rect 1884 214 1942 288
rect 1884 162 1896 214
rect 1930 162 1942 214
rect 1884 88 1942 162
rect 2042 214 2100 288
rect 2042 162 2054 214
rect 2088 162 2100 214
rect 2042 88 2100 162
rect 2200 214 2258 288
rect 2200 162 2212 214
rect 2246 162 2258 214
rect 2200 88 2258 162
rect 2358 214 2416 288
rect 2358 162 2370 214
rect 2404 162 2416 214
rect 2358 88 2416 162
rect 2516 214 2574 288
rect 2516 162 2528 214
rect 2562 162 2574 214
rect 2516 88 2574 162
rect 2770 210 2828 284
rect 2770 158 2782 210
rect 2816 158 2828 210
rect 2770 84 2828 158
rect 2928 210 2986 284
rect 2928 158 2940 210
rect 2974 158 2986 210
rect 2928 84 2986 158
rect 3086 210 3144 284
rect 3086 158 3098 210
rect 3132 158 3144 210
rect 3086 84 3144 158
rect 3244 210 3302 284
rect 3244 158 3256 210
rect 3290 158 3302 210
rect 3244 84 3302 158
rect 3402 210 3460 284
rect 3402 158 3414 210
rect 3448 158 3460 210
rect 3402 84 3460 158
rect 3646 212 3704 286
rect 3646 160 3658 212
rect 3692 160 3704 212
rect 3646 86 3704 160
rect 3804 212 3862 286
rect 3804 160 3816 212
rect 3850 160 3862 212
rect 3804 86 3862 160
rect 3962 212 4020 286
rect 3962 160 3974 212
rect 4008 160 4020 212
rect 3962 86 4020 160
rect 4120 212 4178 286
rect 4120 160 4132 212
rect 4166 160 4178 212
rect 4120 86 4178 160
rect 4278 212 4336 286
rect 4278 160 4290 212
rect 4324 160 4336 212
rect 4278 86 4336 160
rect 4510 210 4568 284
rect 4510 158 4522 210
rect 4556 158 4568 210
rect -1173 -12 -1162 22
rect -1128 -12 -1116 22
rect -1173 -62 -1116 -12
rect -1173 -96 -1162 -62
rect -1128 -96 -1116 -62
rect 4510 84 4568 158
rect 4668 210 4726 284
rect 4668 158 4680 210
rect 4714 158 4726 210
rect 4668 84 4726 158
rect 4826 210 4884 284
rect 4826 158 4838 210
rect 4872 158 4884 210
rect 4826 84 4884 158
rect 4984 210 5042 284
rect 4984 158 4996 210
rect 5030 158 5042 210
rect 4984 84 5042 158
rect 5142 210 5200 284
rect 5142 158 5154 210
rect 5188 158 5200 210
rect 5142 84 5200 158
rect 7492 213 7549 221
rect 6654 195 6711 203
rect 6654 161 6666 195
rect 6700 161 6711 195
rect 6654 112 6711 161
rect 6654 78 6666 112
rect 6700 78 6711 112
rect 6654 28 6711 78
rect 6654 -6 6666 28
rect 6700 -6 6711 28
rect 6654 -55 6711 -6
rect -1173 -145 -1116 -96
rect 6654 -89 6666 -55
rect 6700 -89 6711 -55
rect 6654 -97 6711 -89
rect 6811 195 6868 203
rect 6811 161 6822 195
rect 6856 161 6868 195
rect 6811 112 6868 161
rect 6811 78 6822 112
rect 6856 78 6868 112
rect 6811 28 6868 78
rect 6811 -6 6822 28
rect 6856 -6 6868 28
rect 6811 -55 6868 -6
rect 6811 -89 6822 -55
rect 6856 -89 6868 -55
rect 7492 179 7504 213
rect 7538 179 7549 213
rect 7492 130 7549 179
rect 7492 96 7504 130
rect 7538 96 7549 130
rect 7492 46 7549 96
rect 7492 12 7504 46
rect 7538 12 7549 46
rect 7492 -37 7549 12
rect 7492 -71 7504 -37
rect 7538 -71 7549 -37
rect 7492 -79 7549 -71
rect 7649 213 7706 221
rect 7649 179 7660 213
rect 7694 179 7706 213
rect 7649 130 7706 179
rect 7649 96 7660 130
rect 7694 96 7706 130
rect 7649 46 7706 96
rect 7649 12 7660 46
rect 7694 12 7706 46
rect 7649 -37 7706 12
rect 7649 -71 7660 -37
rect 7694 -71 7706 -37
rect 7649 -79 7706 -71
rect 8312 209 8369 217
rect 8312 175 8324 209
rect 8358 175 8369 209
rect 8312 126 8369 175
rect 8312 92 8324 126
rect 8358 92 8369 126
rect 8312 42 8369 92
rect 8312 8 8324 42
rect 8358 8 8369 42
rect 8312 -41 8369 8
rect 8312 -75 8324 -41
rect 8358 -75 8369 -41
rect 6811 -97 6868 -89
rect -1173 -179 -1162 -145
rect -1128 -179 -1116 -145
rect -1173 -187 -1116 -179
rect 8312 -83 8369 -75
rect 8469 209 8526 217
rect 8469 175 8480 209
rect 8514 175 8526 209
rect 8469 126 8526 175
rect 8469 92 8480 126
rect 8514 92 8526 126
rect 8469 42 8526 92
rect 8469 8 8480 42
rect 8514 8 8526 42
rect 8469 -41 8526 8
rect 8469 -75 8480 -41
rect 8514 -75 8526 -41
rect 8469 -83 8526 -75
rect -260 -896 -202 -822
rect -260 -948 -248 -896
rect -214 -948 -202 -896
rect -260 -1022 -202 -948
rect -102 -896 -44 -822
rect -102 -948 -90 -896
rect -56 -948 -44 -896
rect -102 -1022 -44 -948
rect 56 -896 114 -822
rect 56 -948 68 -896
rect 102 -948 114 -896
rect 56 -1022 114 -948
rect 214 -896 272 -822
rect 214 -948 226 -896
rect 260 -948 272 -896
rect 214 -1022 272 -948
rect 372 -896 430 -822
rect 372 -948 384 -896
rect 418 -948 430 -896
rect 372 -1022 430 -948
rect -260 -1190 -202 -1116
rect -260 -1242 -248 -1190
rect -214 -1242 -202 -1190
rect -260 -1316 -202 -1242
rect -102 -1190 -44 -1116
rect -102 -1242 -90 -1190
rect -56 -1242 -44 -1190
rect -102 -1316 -44 -1242
rect 56 -1190 114 -1116
rect 56 -1242 68 -1190
rect 102 -1242 114 -1190
rect 56 -1316 114 -1242
rect 214 -1190 272 -1116
rect 214 -1242 226 -1190
rect 260 -1242 272 -1190
rect 214 -1316 272 -1242
rect 372 -1190 430 -1116
rect 372 -1242 384 -1190
rect 418 -1242 430 -1190
rect 372 -1316 430 -1242
rect 5096 -870 5154 -796
rect 5096 -922 5108 -870
rect 5142 -922 5154 -870
rect 5096 -996 5154 -922
rect 5254 -870 5312 -796
rect 5254 -922 5266 -870
rect 5300 -922 5312 -870
rect 5254 -996 5312 -922
rect 5412 -870 5470 -796
rect 5412 -922 5424 -870
rect 5458 -922 5470 -870
rect 5412 -996 5470 -922
rect 5570 -870 5628 -796
rect 5570 -922 5582 -870
rect 5616 -922 5628 -870
rect 5570 -996 5628 -922
rect 5728 -870 5786 -796
rect 5728 -922 5740 -870
rect 5774 -922 5786 -870
rect 5728 -996 5786 -922
rect 5096 -1164 5154 -1090
rect 5096 -1216 5108 -1164
rect 5142 -1216 5154 -1164
rect 5096 -1290 5154 -1216
rect 5254 -1164 5312 -1090
rect 5254 -1216 5266 -1164
rect 5300 -1216 5312 -1164
rect 5254 -1290 5312 -1216
rect 5412 -1164 5470 -1090
rect 5412 -1216 5424 -1164
rect 5458 -1216 5470 -1164
rect 5412 -1290 5470 -1216
rect 5570 -1164 5628 -1090
rect 5570 -1216 5582 -1164
rect 5616 -1216 5628 -1164
rect 5570 -1290 5628 -1216
rect 5728 -1164 5786 -1090
rect 5728 -1216 5740 -1164
rect 5774 -1216 5786 -1164
rect 5728 -1290 5786 -1216
<< mvndiffc >>
rect 6670 -325 6704 -291
rect -1322 -415 -1288 -381
rect -1322 -515 -1288 -481
rect -1166 -415 -1132 -381
rect 6670 -425 6704 -391
rect 6826 -325 6860 -291
rect 6826 -425 6860 -391
rect 7508 -307 7542 -273
rect 7508 -407 7542 -373
rect 7664 -307 7698 -273
rect 7664 -407 7698 -373
rect 8328 -311 8362 -277
rect 8328 -411 8362 -377
rect 8484 -311 8518 -277
rect 8484 -411 8518 -377
rect -1166 -515 -1132 -481
rect 1642 -792 1676 -740
rect 1800 -792 1834 -740
rect 1958 -792 1992 -740
rect 2116 -792 2150 -740
rect 2274 -792 2308 -740
rect 3160 -798 3194 -746
rect 3318 -798 3352 -746
rect 3476 -798 3510 -746
rect 3634 -798 3668 -746
rect 3792 -798 3826 -746
rect 1642 -1086 1676 -1034
rect 1800 -1086 1834 -1034
rect 1958 -1086 1992 -1034
rect 2116 -1086 2150 -1034
rect 2274 -1086 2308 -1034
rect 2408 -1096 2442 -1044
rect 2566 -1096 2600 -1044
rect 2724 -1096 2758 -1044
rect 2882 -1096 2916 -1044
rect 3040 -1096 3074 -1044
rect 3160 -1092 3194 -1040
rect 3318 -1092 3352 -1040
rect 3476 -1092 3510 -1040
rect 3634 -1092 3668 -1040
rect 3792 -1092 3826 -1040
rect 892 -1390 926 -1338
rect 1050 -1390 1084 -1338
rect 1208 -1390 1242 -1338
rect 1366 -1390 1400 -1338
rect 1524 -1390 1558 -1338
rect 1642 -1380 1676 -1328
rect 1800 -1380 1834 -1328
rect 1958 -1380 1992 -1328
rect 2116 -1380 2150 -1328
rect 2274 -1380 2308 -1328
rect 2408 -1390 2442 -1338
rect 2566 -1390 2600 -1338
rect 2724 -1390 2758 -1338
rect 2882 -1390 2916 -1338
rect 3040 -1390 3074 -1338
rect 3160 -1386 3194 -1334
rect 3318 -1386 3352 -1334
rect 3476 -1386 3510 -1334
rect 3634 -1386 3668 -1334
rect 3792 -1386 3826 -1334
rect 3910 -1390 3944 -1338
rect 4068 -1390 4102 -1338
rect 4226 -1390 4260 -1338
rect 4384 -1390 4418 -1338
rect 4542 -1390 4576 -1338
rect 7478 -1274 7512 -1222
rect 7636 -1274 7670 -1222
rect 8288 -1264 8322 -1212
rect 8446 -1264 8480 -1212
<< mvpdiffc >>
rect 88 454 122 506
rect 246 454 280 506
rect 404 454 438 506
rect 562 454 596 506
rect 720 454 754 506
rect 992 456 1026 508
rect 1150 456 1184 508
rect 1308 456 1342 508
rect 1466 456 1500 508
rect 1624 456 1658 508
rect 1896 456 1930 508
rect 2054 456 2088 508
rect 2212 456 2246 508
rect 2370 456 2404 508
rect 2528 456 2562 508
rect 2782 452 2816 504
rect 2940 452 2974 504
rect 3098 452 3132 504
rect 3256 452 3290 504
rect 3414 452 3448 504
rect 3658 454 3692 506
rect 3816 454 3850 506
rect 3974 454 4008 506
rect 4132 454 4166 506
rect 4290 454 4324 506
rect 4522 452 4556 504
rect 4680 452 4714 504
rect 4838 452 4872 504
rect 4996 452 5030 504
rect 5154 452 5188 504
rect -1318 71 -1284 105
rect -1318 -12 -1284 22
rect -1318 -96 -1284 -62
rect -1318 -179 -1284 -145
rect -1162 71 -1128 105
rect 88 160 122 212
rect 246 160 280 212
rect 404 160 438 212
rect 562 160 596 212
rect 720 160 754 212
rect 992 162 1026 214
rect 1150 162 1184 214
rect 1308 162 1342 214
rect 1466 162 1500 214
rect 1624 162 1658 214
rect 1896 162 1930 214
rect 2054 162 2088 214
rect 2212 162 2246 214
rect 2370 162 2404 214
rect 2528 162 2562 214
rect 2782 158 2816 210
rect 2940 158 2974 210
rect 3098 158 3132 210
rect 3256 158 3290 210
rect 3414 158 3448 210
rect 3658 160 3692 212
rect 3816 160 3850 212
rect 3974 160 4008 212
rect 4132 160 4166 212
rect 4290 160 4324 212
rect 4522 158 4556 210
rect -1162 -12 -1128 22
rect -1162 -96 -1128 -62
rect 4680 158 4714 210
rect 4838 158 4872 210
rect 4996 158 5030 210
rect 5154 158 5188 210
rect 6666 161 6700 195
rect 6666 78 6700 112
rect 6666 -6 6700 28
rect 6666 -89 6700 -55
rect 6822 161 6856 195
rect 6822 78 6856 112
rect 6822 -6 6856 28
rect 6822 -89 6856 -55
rect 7504 179 7538 213
rect 7504 96 7538 130
rect 7504 12 7538 46
rect 7504 -71 7538 -37
rect 7660 179 7694 213
rect 7660 96 7694 130
rect 7660 12 7694 46
rect 7660 -71 7694 -37
rect 8324 175 8358 209
rect 8324 92 8358 126
rect 8324 8 8358 42
rect 8324 -75 8358 -41
rect -1162 -179 -1128 -145
rect 8480 175 8514 209
rect 8480 92 8514 126
rect 8480 8 8514 42
rect 8480 -75 8514 -41
rect -248 -948 -214 -896
rect -90 -948 -56 -896
rect 68 -948 102 -896
rect 226 -948 260 -896
rect 384 -948 418 -896
rect -248 -1242 -214 -1190
rect -90 -1242 -56 -1190
rect 68 -1242 102 -1190
rect 226 -1242 260 -1190
rect 384 -1242 418 -1190
rect 5108 -922 5142 -870
rect 5266 -922 5300 -870
rect 5424 -922 5458 -870
rect 5582 -922 5616 -870
rect 5740 -922 5774 -870
rect 5108 -1216 5142 -1164
rect 5266 -1216 5300 -1164
rect 5424 -1216 5458 -1164
rect 5582 -1216 5616 -1164
rect 5740 -1216 5774 -1164
<< mvpsubdiff >>
rect -1364 -647 -1333 -613
rect -1299 -647 -1237 -613
rect -1203 -647 -1141 -613
rect -1107 -647 -1076 -613
rect 628 -646 806 -562
rect 628 -1392 648 -646
rect 776 -1392 806 -646
rect 4664 -636 4848 -536
rect 628 -1456 806 -1392
rect 4664 -1386 4690 -636
rect 4818 -1386 4848 -636
rect 6614 -557 6645 -523
rect 6679 -557 6741 -523
rect 6775 -557 6837 -523
rect 6871 -557 6902 -523
rect 7452 -539 7483 -505
rect 7517 -539 7579 -505
rect 7613 -539 7675 -505
rect 7709 -539 7740 -505
rect 8272 -543 8303 -509
rect 8337 -543 8399 -509
rect 8433 -543 8495 -509
rect 8529 -543 8560 -509
rect 4664 -1436 4848 -1386
<< mvnsubdiff >>
rect -202 538 -54 600
rect -1364 167 -1333 201
rect -1299 167 -1237 201
rect -1203 167 -1141 201
rect -1107 167 -1076 201
rect -202 116 -178 538
rect -86 116 -54 538
rect 5338 602 5512 658
rect -202 28 -54 116
rect 5338 66 5370 602
rect 5474 66 5512 602
rect 6614 257 6645 291
rect 6679 257 6741 291
rect 6775 257 6837 291
rect 6871 257 6902 291
rect 7452 275 7483 309
rect 7517 275 7579 309
rect 7613 275 7675 309
rect 7709 275 7740 309
rect 8272 271 8303 305
rect 8337 271 8399 305
rect 8433 271 8495 305
rect 8529 271 8560 305
rect 5338 -6 5512 66
<< mvpsubdiffcont >>
rect -1333 -647 -1299 -613
rect -1237 -647 -1203 -613
rect -1141 -647 -1107 -613
rect 648 -1392 776 -646
rect 4690 -1386 4818 -636
rect 6645 -557 6679 -523
rect 6741 -557 6775 -523
rect 6837 -557 6871 -523
rect 7483 -539 7517 -505
rect 7579 -539 7613 -505
rect 7675 -539 7709 -505
rect 8303 -543 8337 -509
rect 8399 -543 8433 -509
rect 8495 -543 8529 -509
<< mvnsubdiffcont >>
rect -1333 167 -1299 201
rect -1237 167 -1203 201
rect -1141 167 -1107 201
rect -178 116 -86 538
rect 5370 66 5474 602
rect 6645 257 6679 291
rect 6741 257 6775 291
rect 6837 257 6871 291
rect 7483 275 7517 309
rect 7579 275 7613 309
rect 7675 275 7709 309
rect 8303 271 8337 305
rect 8399 271 8433 305
rect 8495 271 8529 305
<< poly >>
rect 1256 870 4862 876
rect 320 838 4862 870
rect 316 776 4862 838
rect 316 646 410 776
rect 1256 772 4862 776
rect 1280 648 1362 772
rect 3878 762 4862 772
rect 3878 728 4858 762
rect 174 606 666 646
rect 1078 608 1570 648
rect 1982 608 2474 648
rect 3878 646 3974 728
rect 134 600 708 606
rect 134 580 234 600
rect 292 580 392 600
rect 450 580 550 600
rect 608 580 708 600
rect 1038 602 1612 608
rect 1038 582 1138 602
rect 1196 582 1296 602
rect 1354 582 1454 602
rect 1512 582 1612 602
rect 1942 602 2516 608
rect 2868 604 3360 644
rect 3744 606 4236 646
rect 4764 644 4858 728
rect 1942 582 2042 602
rect 2100 582 2200 602
rect 2258 582 2358 602
rect 2416 582 2516 602
rect 2828 598 3402 604
rect -1273 113 -1173 139
rect 2828 578 2928 598
rect 2986 578 3086 598
rect 3144 578 3244 598
rect 3302 578 3402 598
rect 3704 600 4278 606
rect 4608 604 5100 644
rect 3704 580 3804 600
rect 3862 580 3962 600
rect 4020 580 4120 600
rect 4178 580 4278 600
rect 4568 598 5142 604
rect 134 354 234 380
rect 292 354 392 380
rect 450 354 550 380
rect 608 354 708 380
rect 1038 356 1138 382
rect 1196 356 1296 382
rect 1354 356 1454 382
rect 1512 356 1612 382
rect 1942 356 2042 382
rect 2100 356 2200 382
rect 2258 356 2358 382
rect 2416 356 2516 382
rect 4568 578 4668 598
rect 4726 578 4826 598
rect 4884 578 4984 598
rect 5042 578 5142 598
rect 152 312 202 354
rect 318 312 368 354
rect 478 312 528 354
rect 634 312 684 354
rect 1056 314 1106 356
rect 1222 314 1272 356
rect 1382 314 1432 356
rect 1538 314 1588 356
rect 1960 314 2010 356
rect 2126 314 2176 356
rect 2286 314 2336 356
rect 2442 314 2492 356
rect 2828 352 2928 378
rect 2986 352 3086 378
rect 3144 352 3244 378
rect 3302 352 3402 378
rect 3704 354 3804 380
rect 3862 354 3962 380
rect 4020 354 4120 380
rect 4178 354 4278 380
rect 134 286 234 312
rect 292 286 392 312
rect 450 286 550 312
rect 608 286 708 312
rect 1038 288 1138 314
rect 1196 288 1296 314
rect 1354 288 1454 314
rect 1512 288 1612 314
rect 1942 288 2042 314
rect 2100 288 2200 314
rect 2258 288 2358 314
rect 2416 288 2516 314
rect 2846 310 2896 352
rect 3012 310 3062 352
rect 3172 310 3222 352
rect 3328 310 3378 352
rect 3722 312 3772 354
rect 3888 312 3938 354
rect 4048 312 4098 354
rect 4204 312 4254 354
rect 4568 352 4668 378
rect 4726 352 4826 378
rect 4884 352 4984 378
rect 5042 352 5142 378
rect 2828 284 2928 310
rect 2986 284 3086 310
rect 3144 284 3244 310
rect 3302 284 3402 310
rect 3704 286 3804 312
rect 3862 286 3962 312
rect 4020 286 4120 312
rect 4178 286 4278 312
rect 4586 310 4636 352
rect 4752 310 4802 352
rect 4912 310 4962 352
rect 5068 310 5118 352
rect 134 60 234 86
rect 292 60 392 86
rect 450 60 550 86
rect 608 60 708 86
rect 1038 62 1138 88
rect 1196 62 1296 88
rect 1354 62 1454 88
rect 1512 62 1612 88
rect 1942 62 2042 88
rect 2100 62 2200 88
rect 2258 70 2358 88
rect 2258 62 2360 70
rect 2416 62 2516 88
rect 4568 284 4668 310
rect 4726 284 4826 310
rect 4884 284 4984 310
rect 5042 284 5142 310
rect 2260 20 2360 62
rect 2828 58 2928 84
rect 2986 58 3086 84
rect 3144 58 3244 84
rect 3302 58 3402 84
rect 3704 60 3804 86
rect 3862 60 3962 86
rect 4020 60 4120 86
rect 4178 60 4278 86
rect 2260 -30 2280 20
rect 2334 -30 2360 20
rect 2260 -70 2360 -30
rect 2830 -2 2924 58
rect 2830 -42 2852 -2
rect 2896 -42 2924 -2
rect 3706 38 3800 60
rect 4568 58 4668 84
rect 4726 58 4826 84
rect 4884 58 4984 84
rect 5042 58 5142 84
rect 6711 203 6811 229
rect 7549 221 7649 247
rect 3706 -10 3724 38
rect 3780 -10 3800 38
rect 3706 -34 3800 -10
rect 2830 -86 2924 -42
rect 8369 217 8469 243
rect 6711 -123 6811 -97
rect 7549 -105 7649 -79
rect 6711 -169 6815 -123
rect -1273 -213 -1173 -187
rect -1277 -259 -1173 -213
rect 6711 -203 6731 -169
rect 6765 -203 6815 -169
rect 6711 -257 6815 -203
rect 7549 -151 7653 -105
rect 7549 -185 7569 -151
rect 7603 -185 7653 -151
rect 7549 -239 7653 -185
rect -1277 -293 -1227 -259
rect -1193 -293 -1173 -259
rect 6715 -283 6815 -257
rect 7553 -265 7653 -239
rect 8369 -109 8469 -83
rect 8369 -155 8473 -109
rect 8369 -189 8389 -155
rect 8423 -189 8473 -155
rect 8369 -243 8473 -189
rect -1277 -347 -1173 -293
rect -1277 -373 -1177 -347
rect 8373 -269 8473 -243
rect 6715 -459 6815 -433
rect 7553 -441 7653 -415
rect 8373 -445 8473 -419
rect 3736 -498 5308 -484
rect 1942 -510 5308 -498
rect -1277 -549 -1177 -523
rect 1940 -524 5308 -510
rect 1940 -536 3774 -524
rect 1940 -606 1976 -536
rect 1734 -640 2216 -606
rect -162 -796 330 -756
rect -202 -802 372 -796
rect -202 -822 -102 -802
rect -44 -822 56 -802
rect 114 -822 214 -802
rect 272 -822 372 -802
rect -202 -1048 -102 -1022
rect -44 -1048 56 -1022
rect 114 -1048 214 -1022
rect 272 -1048 372 -1022
rect -184 -1090 -134 -1048
rect -18 -1090 32 -1048
rect 142 -1090 192 -1048
rect 298 -1090 348 -1048
rect -202 -1116 -102 -1090
rect -44 -1116 56 -1090
rect 114 -1116 214 -1090
rect 272 -1116 372 -1090
rect -202 -1342 -102 -1316
rect -44 -1342 56 -1316
rect 114 -1342 214 -1316
rect 272 -1342 372 -1316
rect 120 -1558 176 -1342
rect 1688 -644 2262 -640
rect 1688 -666 1788 -644
rect 1846 -666 1946 -644
rect 2004 -666 2104 -644
rect 2162 -666 2262 -644
rect 3252 -646 3734 -612
rect 3206 -650 3780 -646
rect 3206 -672 3306 -650
rect 3364 -672 3464 -650
rect 3522 -672 3622 -650
rect 3680 -672 3780 -650
rect 2650 -844 2780 -810
rect 1688 -892 1788 -866
rect 1846 -892 1946 -866
rect 2004 -892 2104 -866
rect 2162 -892 2262 -866
rect 1702 -934 1764 -892
rect 1870 -934 1932 -892
rect 2030 -934 2092 -892
rect 2180 -934 2242 -892
rect 2650 -896 2680 -844
rect 2734 -896 2780 -844
rect 2650 -916 2780 -896
rect 3206 -898 3306 -872
rect 3364 -898 3464 -872
rect 3522 -898 3622 -872
rect 3680 -898 3780 -872
rect 1688 -960 1788 -934
rect 1846 -960 1946 -934
rect 2004 -960 2104 -934
rect 2162 -960 2262 -934
rect 2490 -944 2990 -916
rect 3220 -940 3282 -898
rect 3388 -940 3450 -898
rect 3548 -940 3610 -898
rect 3698 -940 3760 -898
rect 2454 -950 3028 -944
rect 1250 -1142 1424 -1118
rect 1250 -1182 1284 -1142
rect 1382 -1182 1424 -1142
rect 2454 -970 2554 -950
rect 2612 -970 2712 -950
rect 2770 -970 2870 -950
rect 2928 -970 3028 -950
rect 3206 -966 3306 -940
rect 3364 -966 3464 -940
rect 3522 -966 3622 -940
rect 3680 -966 3780 -940
rect 1250 -1204 1424 -1182
rect 1688 -1186 1788 -1160
rect 1846 -1186 1946 -1160
rect 2004 -1186 2104 -1160
rect 2162 -1186 2262 -1160
rect 4172 -1122 4334 -1096
rect 982 -1238 1468 -1204
rect 1704 -1228 1766 -1186
rect 1862 -1228 1924 -1186
rect 2018 -1228 2080 -1186
rect 2184 -1228 2246 -1186
rect 2454 -1196 2554 -1170
rect 2612 -1196 2712 -1170
rect 2770 -1196 2870 -1170
rect 2928 -1196 3028 -1170
rect 3206 -1192 3306 -1166
rect 3364 -1192 3464 -1166
rect 3522 -1192 3622 -1166
rect 3680 -1192 3780 -1166
rect 938 -1244 1512 -1238
rect 938 -1264 1038 -1244
rect 1096 -1264 1196 -1244
rect 1254 -1264 1354 -1244
rect 1412 -1264 1512 -1244
rect 1688 -1254 1788 -1228
rect 1846 -1254 1946 -1228
rect 2004 -1254 2104 -1228
rect 2162 -1254 2262 -1228
rect 2470 -1238 2534 -1196
rect 2630 -1238 2694 -1196
rect 2782 -1238 2846 -1196
rect 2950 -1238 3014 -1196
rect 3222 -1234 3284 -1192
rect 3380 -1234 3442 -1192
rect 3536 -1234 3598 -1192
rect 3702 -1234 3764 -1192
rect 4172 -1204 4202 -1122
rect 4304 -1204 4334 -1122
rect 2454 -1264 2554 -1238
rect 2612 -1264 2712 -1238
rect 2770 -1264 2870 -1238
rect 2928 -1264 3028 -1238
rect 3206 -1260 3306 -1234
rect 3364 -1260 3464 -1234
rect 3522 -1260 3622 -1234
rect 3680 -1260 3780 -1234
rect 4000 -1238 4486 -1204
rect 3956 -1244 4530 -1238
rect 938 -1490 1038 -1464
rect 1096 -1490 1196 -1464
rect 1254 -1490 1354 -1464
rect 1412 -1490 1512 -1464
rect 1688 -1480 1788 -1454
rect 1846 -1480 1946 -1454
rect 2004 -1480 2104 -1454
rect 2162 -1480 2262 -1454
rect 3956 -1264 4056 -1244
rect 4114 -1264 4214 -1244
rect 4272 -1264 4372 -1244
rect 4430 -1264 4530 -1244
rect 2454 -1490 2554 -1464
rect 2612 -1490 2712 -1464
rect 2770 -1490 2870 -1464
rect 2928 -1490 3028 -1464
rect 3206 -1486 3306 -1460
rect 3364 -1486 3464 -1460
rect 3522 -1486 3622 -1460
rect 3680 -1486 3780 -1460
rect 5262 -730 5308 -524
rect 5194 -770 5686 -730
rect 5154 -776 5728 -770
rect 5154 -796 5254 -776
rect 5312 -796 5412 -776
rect 5470 -796 5570 -776
rect 5628 -796 5728 -776
rect 5154 -1022 5254 -996
rect 5312 -1022 5412 -996
rect 5470 -1022 5570 -996
rect 5628 -1022 5728 -996
rect 7530 -1010 7620 -992
rect 5172 -1064 5222 -1022
rect 5338 -1064 5388 -1022
rect 5498 -1064 5548 -1022
rect 5654 -1064 5704 -1022
rect 5154 -1090 5254 -1064
rect 5312 -1090 5412 -1064
rect 5470 -1090 5570 -1064
rect 5628 -1090 5728 -1064
rect 7530 -1098 7544 -1010
rect 7604 -1098 7620 -1010
rect 7530 -1122 7620 -1098
rect 8342 -1008 8426 -982
rect 8342 -1080 8358 -1008
rect 8404 -1080 8426 -1008
rect 8342 -1112 8426 -1080
rect 7524 -1148 7624 -1122
rect 8334 -1138 8434 -1112
rect 5154 -1316 5254 -1290
rect 5312 -1316 5412 -1290
rect 5470 -1316 5570 -1290
rect 5628 -1316 5728 -1290
rect 7524 -1374 7624 -1348
rect 8334 -1364 8434 -1338
rect 3394 -1558 3436 -1486
rect 3956 -1490 4056 -1464
rect 4114 -1490 4214 -1464
rect 4272 -1490 4372 -1464
rect 4430 -1490 4530 -1464
rect 120 -1588 3436 -1558
rect 120 -1590 3432 -1588
<< polycont >>
rect 2280 -30 2334 20
rect 2852 -42 2896 -2
rect 3724 -10 3780 38
rect 6731 -203 6765 -169
rect 7569 -185 7603 -151
rect -1227 -293 -1193 -259
rect 8389 -189 8423 -155
rect 2680 -896 2734 -844
rect 1284 -1182 1382 -1142
rect 4202 -1204 4304 -1122
rect 7544 -1098 7604 -1010
rect 8358 -1080 8404 -1008
<< locali >>
rect 5338 602 5512 658
rect -202 538 -54 600
rect -1364 167 -1333 201
rect -1299 167 -1237 201
rect -1203 167 -1141 201
rect -1107 167 -1076 201
rect -1345 105 -1268 121
rect -1345 71 -1318 105
rect -1284 71 -1268 105
rect -1345 22 -1268 71
rect -1345 -12 -1318 22
rect -1284 -12 -1268 22
rect -1345 -62 -1268 -12
rect -1345 -96 -1318 -62
rect -1284 -96 -1268 -62
rect -1345 -145 -1268 -96
rect -1345 -179 -1318 -145
rect -1284 -179 -1268 -145
rect -1345 -195 -1268 -179
rect -1212 105 -1094 121
rect -1212 71 -1206 105
rect -1172 71 -1162 105
rect -1100 71 -1094 105
rect -1212 22 -1094 71
rect -202 116 -178 538
rect -86 116 -54 538
rect 88 506 122 522
rect 88 438 122 454
rect 246 506 280 522
rect 246 438 280 454
rect 404 506 438 522
rect 404 438 438 454
rect 562 506 596 522
rect 562 438 596 454
rect 720 506 754 522
rect 720 438 754 454
rect 992 508 1026 524
rect 992 440 1026 456
rect 1150 508 1184 524
rect 1150 440 1184 456
rect 1308 508 1342 524
rect 1308 440 1342 456
rect 1466 508 1500 524
rect 1466 440 1500 456
rect 1624 508 1658 524
rect 1624 440 1658 456
rect 1896 508 1930 524
rect 1896 440 1930 456
rect 2054 508 2088 524
rect 2054 440 2088 456
rect 2212 508 2246 524
rect 2212 440 2246 456
rect 2370 508 2404 524
rect 2370 440 2404 456
rect 2528 508 2562 524
rect 2528 440 2562 456
rect 2782 504 2816 520
rect 2782 436 2816 452
rect 2940 504 2974 520
rect 2940 436 2974 452
rect 3098 504 3132 520
rect 3098 436 3132 452
rect 3256 504 3290 520
rect 3256 436 3290 452
rect 3414 504 3448 520
rect 3414 436 3448 452
rect 3658 506 3692 522
rect 3658 438 3692 454
rect 3816 506 3850 522
rect 3816 438 3850 454
rect 3974 506 4008 522
rect 3974 438 4008 454
rect 4132 506 4166 522
rect 4132 438 4166 454
rect 4290 506 4324 522
rect 4290 438 4324 454
rect 4522 504 4556 520
rect 4522 436 4556 452
rect 4680 504 4714 520
rect 4680 436 4714 452
rect 4838 504 4872 520
rect 4838 436 4872 452
rect 4996 504 5030 520
rect 4996 436 5030 452
rect 5154 504 5188 520
rect 5154 436 5188 452
rect 88 212 122 228
rect 88 144 122 160
rect 246 212 280 228
rect 246 144 280 160
rect 404 212 438 228
rect 404 144 438 160
rect 562 212 596 228
rect 562 144 596 160
rect 720 212 754 228
rect 720 144 754 160
rect 992 214 1026 230
rect 992 146 1026 162
rect 1150 214 1184 230
rect 1150 146 1184 162
rect 1308 214 1342 230
rect 1308 146 1342 162
rect 1466 214 1500 230
rect 1466 146 1500 162
rect 1624 214 1658 230
rect 1624 146 1658 162
rect 1896 214 1930 230
rect 1896 146 1930 162
rect 2054 214 2088 230
rect 2054 146 2088 162
rect 2212 214 2246 230
rect 2212 146 2246 162
rect 2370 214 2404 230
rect 2370 146 2404 162
rect 2528 214 2562 230
rect 2528 146 2562 162
rect 2782 210 2816 226
rect 2782 142 2816 158
rect 2940 210 2974 226
rect 2940 142 2974 158
rect 3098 210 3132 226
rect 3098 142 3132 158
rect 3256 210 3290 226
rect 3256 142 3290 158
rect 3414 210 3448 226
rect 3414 142 3448 158
rect 3658 212 3692 228
rect 3658 144 3692 160
rect 3816 212 3850 228
rect 3816 144 3850 160
rect 3974 212 4008 228
rect 3974 144 4008 160
rect 4132 212 4166 228
rect 4132 144 4166 160
rect 4290 212 4324 228
rect 4290 144 4324 160
rect 4522 210 4556 226
rect 4522 142 4556 158
rect 4680 210 4714 226
rect 4680 142 4714 158
rect 4838 210 4872 226
rect 4838 142 4872 158
rect 4996 210 5030 226
rect 4996 142 5030 158
rect 5154 210 5188 226
rect 5154 142 5188 158
rect -202 28 -54 116
rect 5338 66 5370 602
rect 5474 66 5512 602
rect 6614 257 6645 291
rect 6679 257 6741 291
rect 6775 257 6837 291
rect 6871 257 6902 291
rect 7452 275 7483 309
rect 7517 275 7579 309
rect 7613 275 7675 309
rect 7709 275 7740 309
rect 8272 271 8303 305
rect 8337 271 8399 305
rect 8433 271 8495 305
rect 8529 271 8560 305
rect 7470 213 7588 229
rect 3714 38 3796 60
rect -1212 -12 -1162 22
rect -1128 -12 -1094 22
rect -1212 -62 -1094 -12
rect 2264 20 2358 30
rect 2264 -30 2280 20
rect 2334 -30 2358 20
rect 2264 -46 2358 -30
rect 2832 -2 2918 10
rect 2832 -42 2852 -2
rect 2896 -42 2918 -2
rect 3714 -10 3724 38
rect 3780 -10 3796 38
rect 5338 -6 5512 66
rect 6632 195 6750 211
rect 6632 161 6638 195
rect 6700 161 6710 195
rect 6744 161 6750 195
rect 6632 112 6750 161
rect 6632 78 6666 112
rect 6700 78 6750 112
rect 6632 28 6750 78
rect 6632 -6 6666 28
rect 6700 -6 6750 28
rect 3714 -26 3796 -10
rect 2832 -54 2918 -42
rect -1212 -96 -1162 -62
rect -1128 -96 -1094 -62
rect -1212 -145 -1094 -96
rect 6632 -55 6750 -6
rect 6632 -89 6666 -55
rect 6700 -89 6750 -55
rect 6632 -105 6750 -89
rect 6806 195 6883 211
rect 6806 161 6822 195
rect 6856 161 6883 195
rect 6806 112 6883 161
rect 6806 78 6822 112
rect 6856 78 6883 112
rect 6806 28 6883 78
rect 6806 -6 6822 28
rect 6856 -6 6883 28
rect 6806 -55 6883 -6
rect 6806 -89 6822 -55
rect 6856 -89 6883 -55
rect 7470 179 7476 213
rect 7538 179 7548 213
rect 7582 179 7588 213
rect 7470 130 7588 179
rect 7470 96 7504 130
rect 7538 96 7588 130
rect 7470 46 7588 96
rect 7470 12 7504 46
rect 7538 12 7588 46
rect 7470 -37 7588 12
rect 7470 -71 7504 -37
rect 7538 -71 7588 -37
rect 7470 -87 7588 -71
rect 7644 213 7721 229
rect 7644 179 7660 213
rect 7694 179 7721 213
rect 7644 130 7721 179
rect 7644 96 7660 130
rect 7694 96 7721 130
rect 7644 46 7721 96
rect 7644 12 7660 46
rect 7694 12 7721 46
rect 7644 -37 7721 12
rect 7644 -71 7660 -37
rect 7694 -71 7721 -37
rect 7644 -87 7721 -71
rect 6806 -105 6883 -89
rect -1212 -179 -1162 -145
rect -1128 -179 -1094 -145
rect 6639 -156 6781 -153
rect -1212 -195 -1094 -179
rect 6410 -169 6781 -156
rect -1345 -262 -1279 -195
rect 6410 -203 6731 -169
rect 6765 -203 6781 -169
rect 6410 -230 6781 -203
rect 6817 -170 6883 -105
rect 6968 -170 7136 -168
rect 6817 -178 7136 -170
rect 6817 -226 7138 -178
rect 7516 -151 7619 -135
rect 7516 -185 7569 -151
rect 7603 -185 7619 -151
rect 7516 -212 7619 -185
rect 7655 -158 7721 -87
rect 8290 209 8408 225
rect 8290 175 8296 209
rect 8358 175 8368 209
rect 8402 175 8408 209
rect 8290 126 8408 175
rect 8290 92 8324 126
rect 8358 92 8408 126
rect 8290 42 8408 92
rect 8290 8 8324 42
rect 8358 8 8408 42
rect 8290 -41 8408 8
rect 8290 -75 8324 -41
rect 8358 -75 8408 -41
rect 8290 -91 8408 -75
rect 8464 209 8541 225
rect 8464 175 8480 209
rect 8514 175 8541 209
rect 8464 126 8541 175
rect 8464 92 8480 126
rect 8514 92 8541 126
rect 8464 42 8541 92
rect 8464 8 8480 42
rect 8514 8 8541 42
rect 8464 -41 8541 8
rect 8464 -75 8480 -41
rect 8514 -75 8541 -41
rect 8464 -91 8541 -75
rect 8297 -155 8439 -139
rect 8297 -158 8389 -155
rect 7655 -189 8389 -158
rect 8423 -189 8439 -155
rect 7655 -200 8439 -189
rect -1408 -310 -1279 -262
rect -1345 -381 -1279 -310
rect -1243 -252 -1101 -243
rect -1243 -259 -1008 -252
rect -1243 -293 -1227 -259
rect -1193 -293 -1008 -259
rect -1243 -320 -1008 -293
rect -1154 -324 -1008 -320
rect -1345 -415 -1322 -381
rect -1288 -415 -1279 -381
rect -1345 -481 -1279 -415
rect -1345 -515 -1322 -481
rect -1288 -515 -1279 -481
rect -1345 -531 -1279 -515
rect -1212 -381 -1094 -365
rect -1212 -415 -1166 -381
rect -1132 -415 -1094 -381
rect 6410 -238 6722 -230
rect 6410 -328 6466 -238
rect 6632 -291 6750 -275
rect 6632 -325 6670 -291
rect 6704 -325 6750 -291
rect -1212 -481 -1094 -415
rect 6632 -391 6750 -325
rect 6632 -425 6670 -391
rect 6704 -425 6750 -391
rect 6632 -427 6750 -425
rect 6632 -461 6638 -427
rect 6672 -461 6710 -427
rect 6744 -461 6750 -427
rect 6817 -291 6883 -226
rect 6817 -325 6826 -291
rect 6860 -325 6883 -291
rect 6817 -391 6883 -325
rect 6817 -425 6826 -391
rect 6860 -425 6883 -391
rect 6817 -441 6883 -425
rect 6632 -467 6750 -461
rect -1212 -515 -1166 -481
rect -1132 -515 -1094 -481
rect -1212 -517 -1094 -515
rect -1212 -551 -1206 -517
rect -1172 -551 -1134 -517
rect -1100 -551 -1094 -517
rect -1212 -557 -1094 -551
rect -1364 -647 -1333 -613
rect -1299 -647 -1237 -613
rect -1203 -647 -1141 -613
rect -1107 -647 -1076 -613
rect 628 -646 806 -562
rect -248 -896 -214 -880
rect -248 -964 -214 -948
rect -90 -896 -56 -880
rect -90 -964 -56 -948
rect 68 -896 102 -880
rect 68 -964 102 -948
rect 226 -896 260 -880
rect 226 -964 260 -948
rect 384 -896 418 -880
rect 384 -964 418 -948
rect -248 -1190 -214 -1174
rect -248 -1258 -214 -1242
rect -90 -1190 -56 -1174
rect -90 -1258 -56 -1242
rect 68 -1190 102 -1174
rect 68 -1258 102 -1242
rect 226 -1190 260 -1174
rect 226 -1258 260 -1242
rect 384 -1190 418 -1174
rect 384 -1258 418 -1242
rect 628 -1302 648 -646
rect 776 -1302 806 -646
rect 4664 -636 4848 -536
rect 6614 -557 6645 -523
rect 6679 -557 6741 -523
rect 6775 -557 6837 -523
rect 6871 -557 6902 -523
rect 1642 -740 1676 -724
rect 1642 -808 1676 -792
rect 1800 -740 1834 -724
rect 1800 -808 1834 -792
rect 1958 -740 1992 -724
rect 1958 -808 1992 -792
rect 2116 -740 2150 -724
rect 2116 -808 2150 -792
rect 2274 -740 2308 -724
rect 2274 -808 2308 -792
rect 3160 -746 3194 -730
rect 3160 -814 3194 -798
rect 3318 -746 3352 -730
rect 3318 -814 3352 -798
rect 3476 -746 3510 -730
rect 3476 -814 3510 -798
rect 3634 -746 3668 -730
rect 3634 -814 3668 -798
rect 3792 -746 3826 -730
rect 3792 -814 3826 -798
rect 2664 -844 2760 -826
rect 2664 -896 2680 -844
rect 2734 -896 2760 -844
rect 2664 -910 2760 -896
rect 1642 -1034 1676 -1018
rect 1642 -1102 1676 -1086
rect 1800 -1034 1834 -1018
rect 1800 -1102 1834 -1086
rect 1958 -1034 1992 -1018
rect 1958 -1102 1992 -1086
rect 2116 -1034 2150 -1018
rect 2116 -1102 2150 -1086
rect 2274 -1034 2308 -1018
rect 2274 -1102 2308 -1086
rect 2408 -1044 2442 -1028
rect 2408 -1112 2442 -1096
rect 2566 -1044 2600 -1028
rect 2566 -1112 2600 -1096
rect 2724 -1044 2758 -1028
rect 2724 -1112 2758 -1096
rect 2882 -1044 2916 -1028
rect 2882 -1112 2916 -1096
rect 3040 -1044 3074 -1028
rect 3040 -1112 3074 -1096
rect 3160 -1040 3194 -1024
rect 3160 -1108 3194 -1092
rect 3318 -1040 3352 -1024
rect 3318 -1108 3352 -1092
rect 3476 -1040 3510 -1024
rect 3476 -1108 3510 -1092
rect 3634 -1040 3668 -1024
rect 3634 -1108 3668 -1092
rect 3792 -1040 3826 -1024
rect 3792 -1108 3826 -1092
rect 4184 -1122 4322 -1108
rect 1266 -1142 1400 -1134
rect 1266 -1182 1284 -1142
rect 1382 -1182 1400 -1142
rect 1266 -1196 1400 -1182
rect 4184 -1204 4202 -1122
rect 4304 -1204 4322 -1122
rect 4184 -1218 4322 -1204
rect 628 -1400 640 -1302
rect 786 -1400 806 -1302
rect 628 -1456 806 -1400
rect 892 -1338 926 -1322
rect 892 -1406 926 -1390
rect 1050 -1338 1084 -1322
rect 1050 -1406 1084 -1390
rect 1208 -1338 1242 -1322
rect 1208 -1406 1242 -1390
rect 1366 -1338 1400 -1322
rect 1366 -1406 1400 -1390
rect 1524 -1338 1558 -1322
rect 1524 -1406 1558 -1390
rect 1642 -1328 1676 -1312
rect 1642 -1396 1676 -1380
rect 1800 -1328 1834 -1312
rect 1800 -1396 1834 -1380
rect 1958 -1328 1992 -1312
rect 1958 -1396 1992 -1380
rect 2116 -1328 2150 -1312
rect 2116 -1396 2150 -1380
rect 2274 -1328 2308 -1312
rect 2274 -1396 2308 -1380
rect 2408 -1338 2442 -1322
rect 2408 -1406 2442 -1390
rect 2566 -1338 2600 -1322
rect 2566 -1406 2600 -1390
rect 2724 -1338 2758 -1322
rect 2724 -1406 2758 -1390
rect 2882 -1338 2916 -1322
rect 2882 -1406 2916 -1390
rect 3040 -1338 3074 -1322
rect 3040 -1406 3074 -1390
rect 3160 -1334 3194 -1318
rect 3160 -1402 3194 -1386
rect 3318 -1334 3352 -1318
rect 3318 -1402 3352 -1386
rect 3476 -1334 3510 -1318
rect 3476 -1402 3510 -1386
rect 3634 -1334 3668 -1318
rect 3634 -1402 3668 -1386
rect 3792 -1334 3826 -1318
rect 3792 -1402 3826 -1386
rect 3910 -1338 3944 -1322
rect 3910 -1406 3944 -1390
rect 4068 -1338 4102 -1322
rect 4068 -1406 4102 -1390
rect 4226 -1338 4260 -1322
rect 4226 -1406 4260 -1390
rect 4384 -1338 4418 -1322
rect 4384 -1406 4418 -1390
rect 4542 -1338 4576 -1322
rect 4542 -1406 4576 -1390
rect 4664 -1386 4690 -636
rect 4818 -1386 4848 -636
rect 5108 -870 5142 -854
rect 5108 -938 5142 -922
rect 5266 -870 5300 -854
rect 5266 -938 5300 -922
rect 5424 -870 5458 -854
rect 5424 -938 5458 -922
rect 5582 -870 5616 -854
rect 5582 -938 5616 -922
rect 5740 -870 5774 -854
rect 5740 -938 5774 -922
rect 7058 -1012 7138 -226
rect 7470 -273 7588 -257
rect 7470 -307 7508 -273
rect 7542 -307 7588 -273
rect 7470 -373 7588 -307
rect 7470 -407 7508 -373
rect 7542 -407 7588 -373
rect 7470 -409 7588 -407
rect 7470 -443 7476 -409
rect 7510 -443 7548 -409
rect 7582 -443 7588 -409
rect 7655 -273 7721 -200
rect 7952 -268 7998 -200
rect 8297 -216 8439 -200
rect 8475 -180 8541 -91
rect 8475 -216 8654 -180
rect 7655 -307 7664 -273
rect 7698 -307 7721 -273
rect 7655 -373 7721 -307
rect 8290 -277 8408 -261
rect 8290 -311 8328 -277
rect 8362 -311 8408 -277
rect 7655 -407 7664 -373
rect 7698 -407 7721 -373
rect 7655 -423 7721 -407
rect 8290 -377 8408 -311
rect 8290 -411 8328 -377
rect 8362 -411 8408 -377
rect 8290 -413 8408 -411
rect 7470 -449 7588 -443
rect 8290 -447 8296 -413
rect 8330 -447 8368 -413
rect 8402 -447 8408 -413
rect 8475 -277 8541 -216
rect 8475 -311 8484 -277
rect 8518 -311 8541 -277
rect 8475 -377 8541 -311
rect 8475 -411 8484 -377
rect 8518 -411 8541 -377
rect 8475 -427 8541 -411
rect 8290 -453 8408 -447
rect 7452 -539 7483 -505
rect 7517 -539 7579 -505
rect 7613 -539 7675 -505
rect 7709 -539 7740 -505
rect 8272 -543 8303 -509
rect 8337 -543 8399 -509
rect 8433 -543 8495 -509
rect 8529 -543 8560 -509
rect 7530 -1010 7620 -992
rect 7530 -1012 7544 -1010
rect 7058 -1050 7544 -1012
rect 7058 -1052 7138 -1050
rect 7530 -1098 7544 -1050
rect 7604 -1098 7620 -1010
rect 7530 -1130 7620 -1098
rect 8342 -1008 8426 -982
rect 8342 -1080 8358 -1008
rect 8404 -1080 8426 -1008
rect 8342 -1118 8426 -1080
rect 5108 -1164 5142 -1148
rect 5108 -1232 5142 -1216
rect 5266 -1164 5300 -1148
rect 5266 -1232 5300 -1216
rect 5424 -1164 5458 -1148
rect 5424 -1232 5458 -1216
rect 5582 -1164 5616 -1148
rect 5582 -1232 5616 -1216
rect 5740 -1164 5774 -1148
rect 5740 -1232 5774 -1216
rect 7478 -1222 7512 -1206
rect 7478 -1290 7512 -1274
rect 7636 -1222 7670 -1206
rect 7636 -1290 7670 -1274
rect 8288 -1212 8322 -1196
rect 8288 -1280 8322 -1264
rect 8446 -1212 8480 -1196
rect 8446 -1280 8480 -1264
rect 4664 -1436 4848 -1386
<< viali >>
rect -1333 167 -1299 201
rect -1237 167 -1203 201
rect -1141 167 -1107 201
rect -1206 71 -1172 105
rect -1134 71 -1128 105
rect -1128 71 -1100 105
rect -170 142 -92 526
rect 88 454 122 506
rect 246 454 280 506
rect 404 454 438 506
rect 562 454 596 506
rect 720 454 754 506
rect 992 456 1026 508
rect 1150 456 1184 508
rect 1308 456 1342 508
rect 1466 456 1500 508
rect 1624 456 1658 508
rect 1896 456 1930 508
rect 2054 456 2088 508
rect 2212 456 2246 508
rect 2370 456 2404 508
rect 2528 456 2562 508
rect 2782 452 2816 504
rect 2940 452 2974 504
rect 3098 452 3132 504
rect 3256 452 3290 504
rect 3414 452 3448 504
rect 3658 454 3692 506
rect 3816 454 3850 506
rect 3974 454 4008 506
rect 4132 454 4166 506
rect 4290 454 4324 506
rect 4522 452 4556 504
rect 4680 452 4714 504
rect 4838 452 4872 504
rect 4996 452 5030 504
rect 5154 452 5188 504
rect 88 160 122 212
rect 246 160 280 212
rect 404 160 438 212
rect 562 160 596 212
rect 720 160 754 212
rect 992 162 1026 214
rect 1150 162 1184 214
rect 1308 162 1342 214
rect 1466 162 1500 214
rect 1624 162 1658 214
rect 1896 162 1930 214
rect 2054 162 2088 214
rect 2212 162 2246 214
rect 2370 162 2404 214
rect 2528 162 2562 214
rect 2782 158 2816 210
rect 2940 158 2974 210
rect 3098 158 3132 210
rect 3256 158 3290 210
rect 3414 158 3448 210
rect 3658 160 3692 212
rect 3816 160 3850 212
rect 3974 160 4008 212
rect 4132 160 4166 212
rect 4290 160 4324 212
rect 4522 158 4556 210
rect 4680 158 4714 210
rect 4838 158 4872 210
rect 4996 158 5030 210
rect 5154 158 5188 210
rect 5386 124 5444 564
rect 6645 257 6679 291
rect 6741 257 6775 291
rect 6837 257 6871 291
rect 7483 275 7517 309
rect 7579 275 7613 309
rect 7675 275 7709 309
rect 8303 271 8337 305
rect 8399 271 8433 305
rect 8495 271 8529 305
rect 2284 -20 2334 16
rect 2856 -36 2894 -2
rect 3724 -10 3780 38
rect 6638 161 6666 195
rect 6666 161 6672 195
rect 6710 161 6744 195
rect 7476 179 7504 213
rect 7504 179 7510 213
rect 7548 179 7582 213
rect -1544 -324 -1408 -244
rect 7442 -220 7516 -130
rect 8296 175 8324 209
rect 8324 175 8330 209
rect 8368 175 8402 209
rect -1008 -400 -882 -230
rect 6366 -464 6508 -328
rect 6638 -461 6672 -427
rect 6710 -461 6744 -427
rect -1206 -551 -1172 -517
rect -1134 -551 -1100 -517
rect -1333 -647 -1299 -613
rect -1237 -647 -1203 -613
rect -1141 -647 -1107 -613
rect -1116 -804 -1002 -744
rect -248 -948 -214 -896
rect -90 -948 -56 -896
rect 68 -948 102 -896
rect 226 -948 260 -896
rect 384 -948 418 -896
rect -248 -1242 -214 -1190
rect -90 -1242 -56 -1190
rect 68 -1242 102 -1190
rect 226 -1242 260 -1190
rect 384 -1242 418 -1190
rect 658 -1302 770 -704
rect 6645 -557 6679 -523
rect 6741 -557 6775 -523
rect 6837 -557 6871 -523
rect 1642 -792 1676 -740
rect 1800 -792 1834 -740
rect 1958 -792 1992 -740
rect 2116 -792 2150 -740
rect 2274 -792 2308 -740
rect 3160 -798 3194 -746
rect 3318 -798 3352 -746
rect 3476 -798 3510 -746
rect 3634 -798 3668 -746
rect 3792 -798 3826 -746
rect 2680 -896 2734 -844
rect 1642 -1086 1676 -1034
rect 1800 -1086 1834 -1034
rect 1958 -1086 1992 -1034
rect 2116 -1086 2150 -1034
rect 2274 -1086 2308 -1034
rect 2408 -1096 2442 -1044
rect 2566 -1096 2600 -1044
rect 2724 -1096 2758 -1044
rect 2882 -1096 2916 -1044
rect 3040 -1096 3074 -1044
rect 3160 -1092 3194 -1040
rect 3318 -1092 3352 -1040
rect 3476 -1092 3510 -1040
rect 3634 -1092 3668 -1040
rect 3792 -1092 3826 -1040
rect 1284 -1182 1382 -1142
rect 4202 -1204 4304 -1122
rect 640 -1392 648 -1302
rect 648 -1392 776 -1302
rect 776 -1392 786 -1302
rect 640 -1400 786 -1392
rect 892 -1390 926 -1338
rect 1050 -1390 1084 -1338
rect 1208 -1390 1242 -1338
rect 1366 -1390 1400 -1338
rect 1524 -1390 1558 -1338
rect 1642 -1380 1676 -1328
rect 1800 -1380 1834 -1328
rect 1958 -1380 1992 -1328
rect 2116 -1380 2150 -1328
rect 2274 -1380 2308 -1328
rect 2408 -1390 2442 -1338
rect 2566 -1390 2600 -1338
rect 2724 -1390 2758 -1338
rect 2882 -1390 2916 -1338
rect 3040 -1390 3074 -1338
rect 3160 -1386 3194 -1334
rect 3318 -1386 3352 -1334
rect 3476 -1386 3510 -1334
rect 3634 -1386 3668 -1334
rect 3792 -1386 3826 -1334
rect 3910 -1390 3944 -1338
rect 4068 -1390 4102 -1338
rect 4226 -1390 4260 -1338
rect 4384 -1390 4418 -1338
rect 4542 -1390 4576 -1338
rect 4714 -1302 4804 -690
rect 5108 -922 5142 -870
rect 5266 -922 5300 -870
rect 5424 -922 5458 -870
rect 5582 -922 5616 -870
rect 5740 -922 5774 -870
rect 7476 -443 7510 -409
rect 7548 -443 7582 -409
rect 7938 -332 8014 -268
rect 8296 -447 8330 -413
rect 8368 -447 8402 -413
rect 8654 -246 8716 -176
rect 7483 -539 7517 -505
rect 7579 -539 7613 -505
rect 7675 -539 7709 -505
rect 8303 -543 8337 -509
rect 8399 -543 8433 -509
rect 8495 -543 8529 -509
rect 7544 -1098 7604 -1010
rect 8358 -1080 8404 -1008
rect 5108 -1216 5142 -1164
rect 5266 -1216 5300 -1164
rect 5424 -1216 5458 -1164
rect 5582 -1216 5616 -1164
rect 5740 -1216 5774 -1164
rect 7478 -1274 7512 -1222
rect 7636 -1274 7670 -1222
rect 8288 -1264 8322 -1212
rect 8446 -1264 8480 -1212
<< metal1 >>
rect -338 1060 5960 1224
rect -202 600 -60 1060
rect -202 526 -54 600
rect -202 242 -170 526
rect -1136 207 -170 242
rect -1364 201 -170 207
rect -1364 167 -1333 201
rect -1299 167 -1237 201
rect -1203 167 -1141 201
rect -1107 172 -170 201
rect -1107 167 -1076 172
rect -1364 161 -1076 167
rect -1140 133 -1112 161
rect -202 142 -170 172
rect -92 142 -54 526
rect 80 584 130 1060
rect 1618 586 1668 1060
rect 80 552 762 584
rect 990 554 1668 586
rect 80 506 130 552
rect 402 518 436 552
rect 722 518 756 552
rect 992 520 1026 554
rect 1306 520 1340 554
rect 80 490 88 506
rect 82 454 88 490
rect 122 490 130 506
rect 240 506 286 518
rect 122 454 128 490
rect 82 442 128 454
rect 240 454 246 506
rect 280 454 286 506
rect 240 442 286 454
rect 398 506 444 518
rect 398 454 404 506
rect 438 454 444 506
rect 398 442 444 454
rect 556 506 602 518
rect 556 454 562 506
rect 596 454 602 506
rect 556 442 602 454
rect 714 506 760 518
rect 714 454 720 506
rect 754 454 760 506
rect 714 442 760 454
rect 986 508 1032 520
rect 986 456 992 508
rect 1026 456 1032 508
rect 986 444 1032 456
rect 1144 508 1190 520
rect 1144 456 1150 508
rect 1184 456 1190 508
rect 1144 444 1190 456
rect 1302 508 1348 520
rect 1302 456 1308 508
rect 1342 456 1348 508
rect 1302 444 1348 456
rect 1460 508 1506 520
rect 1460 456 1466 508
rect 1500 456 1506 508
rect 1460 444 1506 456
rect 1618 508 1668 554
rect 1618 456 1624 508
rect 1658 492 1668 508
rect 1890 586 1940 1060
rect 1890 554 2570 586
rect 3406 582 3454 1060
rect 3650 584 3700 1060
rect 1890 508 1940 554
rect 2210 520 2244 554
rect 2530 520 2564 554
rect 2780 550 3456 582
rect 3650 552 4332 584
rect 5150 582 5200 1060
rect 5366 658 5508 1060
rect 1658 456 1664 492
rect 1618 444 1664 456
rect 1890 456 1896 508
rect 1930 470 1940 508
rect 2048 508 2094 520
rect 1930 456 1936 470
rect 1890 444 1936 456
rect 2048 456 2054 508
rect 2088 456 2094 508
rect 2048 444 2094 456
rect 2206 508 2252 520
rect 2206 456 2212 508
rect 2246 456 2252 508
rect 2206 444 2252 456
rect 2364 508 2410 520
rect 2364 456 2370 508
rect 2404 456 2410 508
rect 2364 444 2410 456
rect 2522 508 2568 520
rect 2782 516 2816 550
rect 3096 516 3130 550
rect 2522 456 2528 508
rect 2562 456 2568 508
rect 2522 444 2568 456
rect 2776 504 2822 516
rect 2776 452 2782 504
rect 2816 452 2822 504
rect 88 224 124 442
rect 244 224 280 442
rect 402 224 438 442
rect 558 224 594 442
rect 716 224 752 442
rect 992 226 1028 444
rect 1148 226 1184 444
rect 1306 226 1342 444
rect 1462 226 1498 444
rect 1620 226 1656 444
rect 1896 226 1932 444
rect 2052 226 2088 444
rect 2210 226 2246 444
rect 2366 226 2402 444
rect 2524 226 2560 444
rect 2776 440 2822 452
rect 2934 504 2980 516
rect 2934 452 2940 504
rect 2974 452 2980 504
rect 2934 440 2980 452
rect 3092 504 3138 516
rect 3092 452 3098 504
rect 3132 452 3138 504
rect 3092 440 3138 452
rect 3250 504 3296 516
rect 3250 452 3256 504
rect 3290 452 3296 504
rect 3406 504 3454 550
rect 3406 480 3414 504
rect 3250 440 3296 452
rect 3408 452 3414 480
rect 3448 452 3454 504
rect 3650 506 3700 552
rect 3972 518 4006 552
rect 4292 518 4326 552
rect 4520 550 5200 582
rect 3650 490 3658 506
rect 3408 440 3454 452
rect 3652 454 3658 490
rect 3692 490 3700 506
rect 3810 506 3856 518
rect 3692 454 3698 490
rect 3652 442 3698 454
rect 3810 454 3816 506
rect 3850 454 3856 506
rect 3810 442 3856 454
rect 3968 506 4014 518
rect 3968 454 3974 506
rect 4008 454 4014 506
rect 3968 442 4014 454
rect 4126 506 4172 518
rect 4126 454 4132 506
rect 4166 454 4172 506
rect 4126 442 4172 454
rect 4284 506 4330 518
rect 4522 516 4556 550
rect 4836 516 4870 550
rect 5150 516 5200 550
rect 4284 454 4290 506
rect 4324 454 4330 506
rect 4284 442 4330 454
rect 4516 504 4562 516
rect 4516 452 4522 504
rect 4556 452 4562 504
rect 82 212 128 224
rect 82 160 88 212
rect 122 160 128 212
rect 240 212 286 224
rect 240 192 246 212
rect 82 148 128 160
rect 230 160 246 192
rect 280 160 286 212
rect -1364 105 -1076 133
rect -1364 71 -1206 105
rect -1172 71 -1134 105
rect -1100 71 -1076 105
rect -1364 59 -1076 71
rect -202 28 -54 142
rect 230 120 286 160
rect 398 212 444 224
rect 398 160 404 212
rect 438 160 444 212
rect 398 148 444 160
rect 556 212 602 224
rect 556 160 562 212
rect 596 160 602 212
rect 556 148 602 160
rect 714 212 760 224
rect 714 160 720 212
rect 754 160 760 212
rect 714 148 760 160
rect 986 214 1032 226
rect 986 162 992 214
rect 1026 162 1032 214
rect 986 150 1032 162
rect 1144 214 1190 226
rect 1144 162 1150 214
rect 1184 162 1190 214
rect 1144 150 1190 162
rect 1302 214 1348 226
rect 1302 162 1308 214
rect 1342 162 1348 214
rect 1302 150 1348 162
rect 1460 214 1506 226
rect 1460 162 1466 214
rect 1500 162 1506 214
rect 1460 150 1506 162
rect 1618 214 1664 226
rect 1618 162 1624 214
rect 1658 162 1664 214
rect 1618 150 1664 162
rect 1890 214 1936 226
rect 1890 162 1896 214
rect 1930 162 1936 214
rect 1890 150 1936 162
rect 2048 214 2094 226
rect 2048 162 2054 214
rect 2088 162 2094 214
rect 2048 150 2094 162
rect 2206 214 2252 226
rect 2206 162 2212 214
rect 2246 162 2252 214
rect 2206 150 2252 162
rect 2364 214 2410 226
rect 2364 162 2370 214
rect 2404 162 2410 214
rect 2364 150 2410 162
rect 2522 214 2568 226
rect 2782 222 2818 440
rect 2938 222 2974 440
rect 3096 222 3132 440
rect 3252 222 3288 440
rect 3410 222 3446 440
rect 3658 224 3694 442
rect 3814 224 3850 442
rect 3972 224 4008 442
rect 4128 224 4164 442
rect 4286 224 4322 442
rect 4516 440 4562 452
rect 4674 504 4720 516
rect 4674 452 4680 504
rect 4714 452 4720 504
rect 4674 440 4720 452
rect 4832 504 4878 516
rect 4832 452 4838 504
rect 4872 452 4878 504
rect 4832 440 4878 452
rect 4990 504 5036 516
rect 4990 452 4996 504
rect 5030 452 5036 504
rect 4990 440 5036 452
rect 5148 504 5200 516
rect 5148 452 5154 504
rect 5188 484 5200 504
rect 5338 564 5512 658
rect 5188 452 5194 484
rect 5148 440 5194 452
rect 2522 162 2528 214
rect 2562 162 2568 214
rect 2522 150 2568 162
rect 2776 210 2822 222
rect 2776 158 2782 210
rect 2816 158 2822 210
rect 562 120 598 148
rect 1148 122 1188 150
rect 1466 122 1502 150
rect 2052 122 2088 150
rect 2370 122 2406 150
rect 2776 146 2822 158
rect 2934 210 2980 222
rect 2934 158 2940 210
rect 2974 158 2980 210
rect 2934 146 2980 158
rect 3092 210 3138 222
rect 3092 158 3098 210
rect 3132 158 3138 210
rect 3092 146 3138 158
rect 3250 210 3296 222
rect 3250 158 3256 210
rect 3290 158 3296 210
rect 3250 146 3296 158
rect 3408 210 3454 222
rect 3408 158 3414 210
rect 3448 158 3454 210
rect 3408 146 3454 158
rect 3652 212 3698 224
rect 3652 160 3658 212
rect 3692 160 3698 212
rect 3652 148 3698 160
rect 3810 212 3856 224
rect 3810 160 3816 212
rect 3850 160 3856 212
rect 3810 148 3856 160
rect 3968 212 4014 224
rect 3968 160 3974 212
rect 4008 160 4014 212
rect 3968 148 4014 160
rect 4126 212 4172 224
rect 4126 160 4132 212
rect 4166 160 4172 212
rect 4126 148 4172 160
rect 4284 212 4330 224
rect 4522 222 4558 440
rect 4678 222 4714 440
rect 4836 222 4872 440
rect 4992 222 5028 440
rect 5150 222 5186 440
rect 4284 160 4290 212
rect 4324 160 4330 212
rect 4284 148 4330 160
rect 4516 210 4562 222
rect 4516 158 4522 210
rect 4556 158 4562 210
rect 230 88 604 120
rect 1140 118 1508 122
rect 2044 118 2412 122
rect 2938 118 2974 146
rect 3256 118 3292 146
rect 3814 120 3850 148
rect 4132 120 4168 148
rect 4516 146 4562 158
rect 4674 210 4720 222
rect 4674 158 4680 210
rect 4714 158 4720 210
rect 4674 146 4720 158
rect 4832 210 4878 222
rect 4832 158 4838 210
rect 4872 158 4878 210
rect 4832 146 4878 158
rect 4990 210 5036 222
rect 4990 158 4996 210
rect 5030 158 5036 210
rect 4990 146 5036 158
rect 5148 210 5194 222
rect 5148 158 5154 210
rect 5188 158 5194 210
rect 5148 146 5194 158
rect 3806 118 4174 120
rect 4678 118 4714 146
rect 4996 118 5032 146
rect 5338 124 5386 564
rect 5444 312 5512 564
rect 6838 315 7536 318
rect 7692 315 8634 326
rect 5444 297 6670 312
rect 6838 309 8634 315
rect 6838 297 7483 309
rect 5444 291 7483 297
rect 5444 257 6645 291
rect 6679 257 6741 291
rect 6775 257 6837 291
rect 6871 276 7483 291
rect 6871 257 6902 276
rect 7452 275 7483 276
rect 7517 275 7579 309
rect 7613 275 7675 309
rect 7709 305 8634 309
rect 7709 284 8303 305
rect 7709 275 7740 284
rect 8180 280 8303 284
rect 7452 269 7740 275
rect 8272 271 8303 280
rect 8337 271 8399 305
rect 8433 271 8495 305
rect 8529 284 8634 305
rect 8529 271 8560 284
rect 5444 256 6902 257
rect 5444 124 5512 256
rect 6614 251 6902 256
rect 6640 223 6676 251
rect 7478 241 7526 269
rect 8272 265 8560 271
rect 6614 195 6902 223
rect 6614 161 6638 195
rect 6672 161 6710 195
rect 6744 161 6902 195
rect 7452 213 7740 241
rect 8496 237 8544 265
rect 7452 179 7476 213
rect 7510 179 7548 213
rect 7582 179 7740 213
rect 7452 167 7740 179
rect 8272 209 8560 237
rect 8272 175 8296 209
rect 8330 175 8368 209
rect 8402 175 8560 209
rect 8272 163 8560 175
rect 6614 149 6902 161
rect 1140 104 2676 118
rect 1140 90 2678 104
rect 230 -184 286 88
rect 1154 -114 1188 90
rect 2348 86 2678 90
rect 2930 90 4174 118
rect 2930 86 3298 90
rect 3806 88 4174 90
rect 2264 16 2358 30
rect 2264 -20 2284 16
rect 2334 -20 2358 16
rect 2264 -46 2358 -20
rect 2636 -4 2678 86
rect 2832 -2 2918 10
rect 2832 -4 2856 -2
rect 2636 -36 2856 -4
rect 2894 -36 2918 -2
rect 2636 -40 2918 -36
rect 1272 -114 1282 -52
rect 1152 -170 1282 -114
rect -1014 -230 -876 -218
rect -1556 -244 -1396 -238
rect -1556 -324 -1544 -244
rect -1408 -324 -1396 -244
rect -1556 -330 -1396 -324
rect -1528 -634 -1472 -330
rect -1018 -400 -1008 -230
rect -882 -400 -872 -230
rect -1014 -412 -876 -400
rect -1364 -517 -1076 -505
rect -1364 -551 -1206 -517
rect -1172 -551 -1134 -517
rect -1100 -551 -1076 -517
rect -1364 -579 -1076 -551
rect -1116 -607 -1088 -579
rect -1364 -613 -1076 -607
rect -1576 -688 -1566 -634
rect -1440 -688 -1430 -634
rect -1364 -647 -1333 -613
rect -1299 -647 -1237 -613
rect -1203 -647 -1141 -613
rect -1107 -647 -1076 -613
rect 228 -638 290 -184
rect 1154 -244 1188 -170
rect 1272 -222 1282 -170
rect 1396 -222 1406 -52
rect 2282 -150 2330 -46
rect 2832 -54 2918 -40
rect 2994 -150 3030 86
rect 3714 38 3796 60
rect 3714 6 3724 38
rect 3704 -10 3724 6
rect 3780 -10 3796 38
rect 3704 -26 3796 -10
rect 3704 -54 3788 -26
rect 2282 -182 3032 -150
rect 1006 -372 1016 -244
rect 1170 -372 1188 -244
rect 2690 -328 2734 -316
rect 3704 -328 3758 -54
rect 348 -638 358 -604
rect -1364 -653 -1076 -647
rect -1116 -738 -1088 -653
rect 216 -694 358 -638
rect -1128 -744 -990 -738
rect -1128 -804 -1116 -744
rect -1002 -804 -990 -744
rect -1128 -810 -990 -804
rect 228 -818 290 -694
rect 348 -716 358 -694
rect 530 -716 540 -604
rect 628 -704 806 -562
rect -250 -850 426 -818
rect -248 -884 -214 -850
rect 66 -884 100 -850
rect 386 -884 420 -850
rect -254 -896 -208 -884
rect -254 -948 -248 -896
rect -214 -948 -208 -896
rect -254 -960 -208 -948
rect -96 -896 -50 -884
rect -96 -948 -90 -896
rect -56 -948 -50 -896
rect -96 -960 -50 -948
rect 62 -896 108 -884
rect 62 -948 68 -896
rect 102 -948 108 -896
rect 62 -960 108 -948
rect 220 -896 266 -884
rect 220 -948 226 -896
rect 260 -948 266 -896
rect 220 -960 266 -948
rect 378 -896 424 -884
rect 378 -948 384 -896
rect 418 -948 424 -896
rect 378 -960 424 -948
rect -248 -1178 -212 -960
rect -92 -1178 -56 -960
rect 66 -1178 102 -960
rect 222 -1178 258 -960
rect 380 -1178 416 -960
rect -254 -1190 -208 -1178
rect -254 -1242 -248 -1190
rect -214 -1242 -208 -1190
rect -254 -1254 -208 -1242
rect -96 -1190 -50 -1178
rect -96 -1242 -90 -1190
rect -56 -1242 -50 -1190
rect -96 -1254 -50 -1242
rect 62 -1190 108 -1178
rect 62 -1242 68 -1190
rect 102 -1242 108 -1190
rect 62 -1254 108 -1242
rect 220 -1190 266 -1178
rect 220 -1242 226 -1190
rect 260 -1242 266 -1190
rect 220 -1254 266 -1242
rect 378 -1190 424 -1178
rect 378 -1242 384 -1190
rect 418 -1242 424 -1190
rect 378 -1254 424 -1242
rect -92 -1282 -56 -1254
rect 226 -1282 262 -1254
rect -100 -1314 268 -1282
rect 628 -1302 658 -704
rect 770 -1302 806 -704
rect 1154 -1264 1188 -372
rect 1268 -424 1278 -340
rect 1386 -424 1396 -340
rect 2690 -374 3758 -328
rect 1302 -1134 1354 -424
rect 1462 -728 1472 -614
rect 1582 -658 1592 -614
rect 1582 -664 1692 -658
rect 1582 -694 2318 -664
rect 1582 -728 1692 -694
rect 1952 -728 1996 -694
rect 2272 -728 2316 -694
rect 1636 -740 1684 -728
rect 1636 -792 1642 -740
rect 1676 -760 1684 -740
rect 1794 -740 1840 -728
rect 1676 -792 1682 -760
rect 1636 -804 1682 -792
rect 1794 -792 1800 -740
rect 1834 -792 1840 -740
rect 1794 -804 1840 -792
rect 1952 -740 1998 -728
rect 1952 -792 1958 -740
rect 1992 -792 1998 -740
rect 1952 -804 1998 -792
rect 2110 -740 2156 -728
rect 2110 -792 2116 -740
rect 2150 -792 2156 -740
rect 2110 -804 2156 -792
rect 2268 -740 2316 -728
rect 2268 -792 2274 -740
rect 2308 -762 2316 -740
rect 2308 -792 2314 -762
rect 2268 -804 2314 -792
rect 1638 -1022 1674 -804
rect 1798 -1022 1834 -804
rect 1958 -1022 1994 -804
rect 2114 -1022 2150 -804
rect 2270 -1022 2306 -804
rect 2690 -826 2734 -374
rect 3804 -414 3814 -356
rect 3896 -366 3906 -356
rect 3938 -358 3980 88
rect 4670 86 5038 118
rect 4178 -166 4188 -78
rect 4338 -166 4348 -78
rect 4870 -154 4914 86
rect 5338 -6 5512 124
rect 7436 -130 7522 -118
rect 5488 -154 5534 -150
rect 4014 -358 4024 -340
rect 3938 -366 4024 -358
rect 3896 -394 4024 -366
rect 3896 -414 3906 -394
rect 3938 -416 4024 -394
rect 3800 -670 3810 -656
rect 3154 -700 3810 -670
rect 3158 -734 3202 -700
rect 3470 -734 3514 -700
rect 3790 -712 3810 -700
rect 3886 -712 3896 -656
rect 3790 -734 3834 -712
rect 3154 -746 3202 -734
rect 3154 -798 3160 -746
rect 3194 -766 3202 -746
rect 3312 -746 3358 -734
rect 3194 -798 3200 -766
rect 3154 -810 3200 -798
rect 3312 -798 3318 -746
rect 3352 -798 3358 -746
rect 3312 -810 3358 -798
rect 3470 -746 3516 -734
rect 3470 -798 3476 -746
rect 3510 -798 3516 -746
rect 3470 -810 3516 -798
rect 3628 -746 3674 -734
rect 3628 -798 3634 -746
rect 3668 -798 3674 -746
rect 3628 -810 3674 -798
rect 3786 -746 3834 -734
rect 3786 -798 3792 -746
rect 3826 -768 3834 -746
rect 3826 -798 3832 -768
rect 3786 -810 3832 -798
rect 2664 -844 2760 -826
rect 2664 -896 2680 -844
rect 2734 -896 2760 -844
rect 2664 -910 2760 -896
rect 2402 -1000 3086 -972
rect 1636 -1034 1682 -1022
rect 1636 -1086 1642 -1034
rect 1676 -1086 1682 -1034
rect 1636 -1098 1682 -1086
rect 1794 -1034 1840 -1022
rect 1794 -1086 1800 -1034
rect 1834 -1086 1840 -1034
rect 1794 -1098 1840 -1086
rect 1952 -1034 1998 -1022
rect 1952 -1086 1958 -1034
rect 1992 -1086 1998 -1034
rect 1952 -1098 1998 -1086
rect 2110 -1034 2156 -1022
rect 2110 -1086 2116 -1034
rect 2150 -1086 2156 -1034
rect 2110 -1098 2156 -1086
rect 2268 -1034 2314 -1022
rect 2408 -1032 2446 -1000
rect 2720 -1032 2758 -1000
rect 3042 -1032 3080 -1000
rect 3156 -1028 3192 -810
rect 3316 -1028 3352 -810
rect 3476 -1028 3512 -810
rect 3632 -1028 3668 -810
rect 3788 -1028 3824 -810
rect 2268 -1086 2274 -1034
rect 2308 -1086 2314 -1034
rect 2268 -1098 2314 -1086
rect 2402 -1044 2448 -1032
rect 2402 -1096 2408 -1044
rect 2442 -1096 2448 -1044
rect 1266 -1142 1400 -1134
rect 1266 -1182 1284 -1142
rect 1382 -1182 1400 -1142
rect 1266 -1196 1400 -1182
rect 1520 -1264 1550 -1262
rect 882 -1292 1568 -1264
rect 236 -1444 266 -1314
rect 628 -1400 640 -1302
rect 786 -1400 806 -1302
rect 890 -1326 920 -1292
rect 1208 -1326 1238 -1292
rect 1520 -1326 1550 -1292
rect 1638 -1316 1674 -1098
rect 1798 -1316 1834 -1098
rect 1958 -1316 1994 -1098
rect 2114 -1316 2150 -1098
rect 2270 -1316 2306 -1098
rect 2402 -1108 2448 -1096
rect 2560 -1044 2606 -1032
rect 2560 -1096 2566 -1044
rect 2600 -1096 2606 -1044
rect 2560 -1108 2606 -1096
rect 2718 -1044 2764 -1032
rect 2718 -1096 2724 -1044
rect 2758 -1096 2764 -1044
rect 2718 -1108 2764 -1096
rect 2876 -1044 2922 -1032
rect 2876 -1096 2882 -1044
rect 2916 -1096 2922 -1044
rect 2876 -1108 2922 -1096
rect 3034 -1044 3080 -1032
rect 3034 -1096 3040 -1044
rect 3074 -1096 3080 -1044
rect 3034 -1108 3080 -1096
rect 3154 -1040 3200 -1028
rect 3154 -1092 3160 -1040
rect 3194 -1092 3200 -1040
rect 3154 -1104 3200 -1092
rect 3312 -1040 3358 -1028
rect 3312 -1092 3318 -1040
rect 3352 -1092 3358 -1040
rect 3312 -1104 3358 -1092
rect 3470 -1040 3516 -1028
rect 3470 -1092 3476 -1040
rect 3510 -1092 3516 -1040
rect 3470 -1104 3516 -1092
rect 3628 -1040 3674 -1028
rect 3628 -1092 3634 -1040
rect 3668 -1092 3674 -1040
rect 3628 -1104 3674 -1092
rect 3786 -1040 3832 -1028
rect 3786 -1092 3792 -1040
rect 3826 -1092 3832 -1040
rect 3786 -1104 3832 -1092
rect 220 -1532 230 -1444
rect 300 -1532 310 -1444
rect 628 -1456 806 -1400
rect 886 -1338 932 -1326
rect 886 -1390 892 -1338
rect 926 -1390 932 -1338
rect 886 -1402 932 -1390
rect 1044 -1338 1090 -1326
rect 1044 -1390 1050 -1338
rect 1084 -1390 1090 -1338
rect 1044 -1402 1090 -1390
rect 1202 -1338 1248 -1326
rect 1202 -1390 1208 -1338
rect 1242 -1390 1248 -1338
rect 1202 -1402 1248 -1390
rect 1360 -1338 1406 -1326
rect 1360 -1390 1366 -1338
rect 1400 -1390 1406 -1338
rect 1360 -1402 1406 -1390
rect 1518 -1338 1564 -1326
rect 1518 -1390 1524 -1338
rect 1558 -1390 1564 -1338
rect 1518 -1402 1564 -1390
rect 1636 -1328 1682 -1316
rect 1636 -1380 1642 -1328
rect 1676 -1380 1682 -1328
rect 1794 -1328 1840 -1316
rect 1794 -1350 1800 -1328
rect 1636 -1392 1682 -1380
rect 1792 -1380 1800 -1350
rect 1834 -1380 1840 -1328
rect 1792 -1392 1840 -1380
rect 1952 -1328 1998 -1316
rect 1952 -1380 1958 -1328
rect 1992 -1380 1998 -1328
rect 1952 -1392 1998 -1380
rect 2110 -1328 2156 -1316
rect 2110 -1380 2116 -1328
rect 2150 -1380 2156 -1328
rect 2110 -1392 2156 -1380
rect 2268 -1328 2314 -1316
rect 2406 -1326 2438 -1108
rect 2564 -1326 2596 -1108
rect 2722 -1326 2754 -1108
rect 2880 -1326 2912 -1108
rect 3038 -1326 3070 -1108
rect 3156 -1322 3192 -1104
rect 3316 -1322 3352 -1104
rect 3476 -1322 3512 -1104
rect 3632 -1322 3668 -1104
rect 3788 -1322 3824 -1104
rect 3938 -1264 3980 -416
rect 4014 -432 4024 -416
rect 4142 -432 4152 -340
rect 4224 -1108 4270 -166
rect 4870 -184 5536 -154
rect 4664 -690 4848 -536
rect 5488 -646 5534 -184
rect 7432 -220 7442 -130
rect 7516 -220 7526 -130
rect 8648 -176 8722 -164
rect 7436 -232 7522 -220
rect 8644 -246 8654 -176
rect 8716 -246 8726 -176
rect 8648 -258 8722 -246
rect 7926 -268 8026 -262
rect 6354 -328 6520 -322
rect 6354 -464 6366 -328
rect 6508 -464 6520 -328
rect 7926 -332 7938 -268
rect 8014 -332 8026 -268
rect 7926 -338 8026 -332
rect 7452 -409 7740 -397
rect 6354 -470 6520 -464
rect 6614 -427 6902 -415
rect 6614 -461 6638 -427
rect 6672 -461 6710 -427
rect 6744 -461 6902 -427
rect 6614 -489 6902 -461
rect 7452 -443 7476 -409
rect 7510 -443 7548 -409
rect 7582 -443 7740 -409
rect 7452 -471 7740 -443
rect 8272 -413 8560 -401
rect 8272 -447 8296 -413
rect 8330 -447 8368 -413
rect 8402 -447 8560 -413
rect 6640 -517 6676 -489
rect 7472 -499 7500 -471
rect 8272 -475 8560 -447
rect 7452 -505 7740 -499
rect 8356 -503 8404 -475
rect 6614 -522 6902 -517
rect 7452 -522 7483 -505
rect 6614 -523 7483 -522
rect 6614 -557 6645 -523
rect 6679 -557 6741 -523
rect 6775 -557 6837 -523
rect 6871 -539 7483 -523
rect 7517 -539 7579 -505
rect 7613 -539 7675 -505
rect 7709 -522 7740 -505
rect 8272 -509 8560 -503
rect 7709 -524 8198 -522
rect 8272 -524 8303 -509
rect 7709 -539 8303 -524
rect 6871 -543 8303 -539
rect 8337 -543 8399 -509
rect 8433 -543 8495 -509
rect 8529 -522 8560 -509
rect 8529 -543 8634 -522
rect 6871 -545 8634 -543
rect 6871 -557 7512 -545
rect 6614 -563 7512 -557
rect 4184 -1122 4322 -1108
rect 4184 -1204 4202 -1122
rect 4304 -1204 4322 -1122
rect 4184 -1218 4322 -1204
rect 4538 -1264 4568 -1262
rect 3900 -1292 4586 -1264
rect 2268 -1380 2274 -1328
rect 2308 -1380 2314 -1328
rect 2268 -1392 2314 -1380
rect 2402 -1338 2448 -1326
rect 2402 -1390 2408 -1338
rect 2442 -1390 2448 -1338
rect 1052 -1432 1082 -1402
rect 1368 -1432 1398 -1402
rect 1644 -1432 1680 -1392
rect 648 -1666 742 -1456
rect 1042 -1462 1680 -1432
rect 1792 -1424 1826 -1392
rect 2112 -1424 2146 -1392
rect 2402 -1402 2448 -1390
rect 2560 -1338 2606 -1326
rect 2560 -1390 2566 -1338
rect 2600 -1390 2606 -1338
rect 2560 -1402 2606 -1390
rect 2718 -1338 2764 -1326
rect 2718 -1390 2724 -1338
rect 2758 -1390 2764 -1338
rect 2718 -1402 2764 -1390
rect 2876 -1338 2922 -1326
rect 2876 -1390 2882 -1338
rect 2916 -1390 2922 -1338
rect 2876 -1402 2922 -1390
rect 3034 -1338 3080 -1326
rect 3034 -1390 3040 -1338
rect 3074 -1390 3080 -1338
rect 3034 -1402 3080 -1390
rect 3154 -1334 3200 -1322
rect 3154 -1386 3160 -1334
rect 3194 -1386 3200 -1334
rect 3312 -1334 3358 -1322
rect 3312 -1356 3318 -1334
rect 3154 -1398 3200 -1386
rect 3310 -1386 3318 -1356
rect 3352 -1386 3358 -1334
rect 3310 -1398 3358 -1386
rect 3470 -1334 3516 -1322
rect 3470 -1386 3476 -1334
rect 3510 -1386 3516 -1334
rect 3470 -1398 3516 -1386
rect 3628 -1334 3674 -1322
rect 3628 -1386 3634 -1334
rect 3668 -1386 3674 -1334
rect 3628 -1398 3674 -1386
rect 3786 -1334 3832 -1322
rect 3908 -1326 3938 -1292
rect 4226 -1326 4256 -1292
rect 4538 -1326 4568 -1292
rect 4664 -1302 4714 -690
rect 4804 -1302 4848 -690
rect 5414 -716 5424 -646
rect 5516 -716 5534 -646
rect 6624 -682 6670 -563
rect 6850 -566 7512 -563
rect 7692 -566 8634 -545
rect 8192 -568 8506 -566
rect 5488 -792 5534 -716
rect 6578 -752 6588 -682
rect 6668 -752 6678 -682
rect 7414 -750 7424 -678
rect 7544 -750 7554 -678
rect 5106 -824 5782 -792
rect 5108 -858 5142 -824
rect 5422 -858 5456 -824
rect 5488 -826 5534 -824
rect 5742 -858 5776 -824
rect 5102 -870 5148 -858
rect 5102 -922 5108 -870
rect 5142 -922 5148 -870
rect 5102 -934 5148 -922
rect 5260 -870 5306 -858
rect 5260 -922 5266 -870
rect 5300 -922 5306 -870
rect 5260 -934 5306 -922
rect 5418 -870 5464 -858
rect 5418 -922 5424 -870
rect 5458 -922 5464 -870
rect 5418 -934 5464 -922
rect 5576 -870 5622 -858
rect 5576 -922 5582 -870
rect 5616 -922 5622 -870
rect 5576 -934 5622 -922
rect 5734 -870 5780 -858
rect 5734 -922 5740 -870
rect 5774 -922 5780 -870
rect 5734 -934 5780 -922
rect 5108 -1152 5144 -934
rect 5264 -1152 5300 -934
rect 5422 -1152 5458 -934
rect 5578 -1152 5614 -934
rect 5736 -1152 5772 -934
rect 5102 -1164 5148 -1152
rect 5102 -1216 5108 -1164
rect 5142 -1216 5148 -1164
rect 5102 -1228 5148 -1216
rect 5260 -1164 5306 -1152
rect 5260 -1216 5266 -1164
rect 5300 -1216 5306 -1164
rect 5260 -1228 5306 -1216
rect 5418 -1164 5464 -1152
rect 5418 -1216 5424 -1164
rect 5458 -1216 5464 -1164
rect 5418 -1228 5464 -1216
rect 5576 -1164 5622 -1152
rect 5576 -1216 5582 -1164
rect 5616 -1216 5622 -1164
rect 5576 -1228 5622 -1216
rect 5734 -1164 5780 -1152
rect 5734 -1216 5740 -1164
rect 5774 -1216 5780 -1164
rect 5734 -1228 5780 -1216
rect 7466 -1210 7502 -750
rect 8234 -774 8244 -638
rect 8338 -774 8348 -638
rect 7530 -1010 7620 -992
rect 7530 -1098 7544 -1010
rect 7604 -1098 7620 -1010
rect 7530 -1130 7620 -1098
rect 8280 -1200 8308 -774
rect 8342 -1008 8426 -982
rect 8342 -1080 8358 -1008
rect 8404 -1022 8426 -1008
rect 8628 -1022 8638 -960
rect 8404 -1064 8638 -1022
rect 8404 -1080 8426 -1064
rect 8342 -1118 8426 -1080
rect 8628 -1116 8638 -1064
rect 8814 -1116 8824 -960
rect 7466 -1222 7518 -1210
rect 5264 -1256 5300 -1228
rect 5582 -1256 5618 -1228
rect 7466 -1232 7478 -1222
rect 5256 -1288 5624 -1256
rect 7472 -1274 7478 -1232
rect 7512 -1274 7518 -1222
rect 7472 -1286 7518 -1274
rect 7630 -1222 7676 -1210
rect 7630 -1274 7636 -1222
rect 7670 -1274 7676 -1222
rect 8280 -1212 8328 -1200
rect 8280 -1234 8288 -1212
rect 7630 -1286 7676 -1274
rect 8282 -1264 8288 -1234
rect 8322 -1264 8328 -1212
rect 8282 -1276 8328 -1264
rect 8440 -1212 8486 -1200
rect 8440 -1264 8446 -1212
rect 8480 -1258 8486 -1212
rect 8480 -1264 8490 -1258
rect 8440 -1276 8490 -1264
rect 3786 -1386 3792 -1334
rect 3826 -1358 3832 -1334
rect 3904 -1338 3950 -1326
rect 3826 -1386 3834 -1358
rect 3786 -1398 3834 -1386
rect 2402 -1424 2442 -1402
rect 1792 -1446 2442 -1424
rect 2564 -1436 2598 -1402
rect 2886 -1436 2920 -1402
rect 3036 -1432 3080 -1402
rect 3310 -1430 3344 -1398
rect 3630 -1430 3664 -1398
rect 3310 -1432 3678 -1430
rect 1396 -1468 1680 -1462
rect 1780 -1514 1790 -1446
rect 1852 -1452 2442 -1446
rect 1852 -1454 2160 -1452
rect 1852 -1514 1862 -1454
rect 2402 -1526 2442 -1452
rect 2552 -1464 2924 -1436
rect 3036 -1448 3678 -1432
rect 3794 -1440 3834 -1398
rect 3904 -1390 3910 -1338
rect 3944 -1390 3950 -1338
rect 3904 -1402 3950 -1390
rect 4062 -1338 4108 -1326
rect 4062 -1390 4068 -1338
rect 4102 -1390 4108 -1338
rect 4062 -1402 4108 -1390
rect 4220 -1338 4266 -1326
rect 4220 -1390 4226 -1338
rect 4260 -1390 4266 -1338
rect 4220 -1402 4266 -1390
rect 4378 -1338 4424 -1326
rect 4378 -1390 4384 -1338
rect 4418 -1390 4424 -1338
rect 4378 -1402 4424 -1390
rect 4536 -1338 4582 -1326
rect 4536 -1390 4542 -1338
rect 4576 -1390 4582 -1338
rect 4536 -1402 4582 -1390
rect 4664 -1362 4848 -1302
rect 4964 -1362 4974 -1344
rect 4070 -1432 4100 -1402
rect 4386 -1432 4416 -1402
rect 4664 -1424 4974 -1362
rect 4060 -1440 4424 -1432
rect 4664 -1436 4848 -1424
rect 3036 -1460 3616 -1448
rect 2702 -1666 2770 -1464
rect 3036 -1466 3388 -1460
rect 3606 -1520 3616 -1460
rect 3676 -1520 3686 -1448
rect 3794 -1462 4424 -1440
rect 3794 -1472 4092 -1462
rect 4702 -1666 4796 -1436
rect 4964 -1452 4974 -1424
rect 5064 -1452 5074 -1344
rect 5404 -1558 5446 -1288
rect 5370 -1628 5380 -1558
rect 5484 -1628 5494 -1558
rect 7638 -1664 7674 -1286
rect 8442 -1664 8490 -1276
rect 5966 -1666 8276 -1664
rect 8324 -1666 8918 -1664
rect -372 -1898 8918 -1666
rect 5966 -1904 8918 -1898
<< via1 >>
rect -1008 -400 -882 -230
rect -1566 -688 -1440 -634
rect 1282 -222 1396 -52
rect 1016 -372 1170 -244
rect -1116 -804 -1002 -744
rect 358 -716 530 -604
rect 1278 -424 1386 -340
rect 1472 -728 1582 -614
rect 3814 -414 3896 -356
rect 4188 -166 4338 -78
rect 3810 -712 3886 -656
rect 640 -1400 786 -1302
rect 230 -1532 300 -1444
rect 4024 -432 4142 -340
rect 7442 -220 7516 -130
rect 8654 -246 8716 -176
rect 6366 -464 6508 -328
rect 7938 -332 8014 -268
rect 5424 -716 5516 -646
rect 6588 -752 6668 -682
rect 7424 -750 7544 -678
rect 8244 -774 8338 -638
rect 8638 -1116 8814 -960
rect 1790 -1514 1852 -1446
rect 3616 -1520 3676 -1448
rect 4974 -1452 5064 -1344
rect 5380 -1628 5484 -1558
<< metal2 >>
rect 1282 -52 1396 -42
rect -1008 -230 -882 -220
rect 4188 -78 4338 -68
rect 1396 -160 4188 -114
rect 4188 -176 4338 -166
rect 7442 -130 7516 -120
rect 1282 -232 1396 -222
rect 7434 -220 7442 -180
rect 7434 -230 7516 -220
rect 8654 -176 8716 -166
rect 1016 -244 1170 -234
rect -882 -342 1016 -268
rect 6366 -328 6508 -318
rect 1016 -382 1170 -372
rect 1278 -340 1386 -330
rect -1008 -410 -882 -400
rect 4024 -340 4142 -330
rect 3814 -356 3896 -346
rect 1386 -406 3814 -372
rect 3814 -424 3896 -414
rect 1278 -434 1386 -424
rect 4142 -420 6366 -358
rect 4024 -442 4142 -432
rect 6366 -474 6508 -464
rect 7434 -580 7482 -230
rect 8654 -256 8716 -246
rect 7938 -268 8014 -258
rect 7938 -342 8014 -332
rect 7434 -590 7520 -580
rect 8660 -588 8704 -256
rect 8102 -590 8704 -588
rect 358 -604 530 -594
rect -1566 -634 -1440 -624
rect -1566 -698 -1440 -688
rect -1540 -1718 -1458 -698
rect 1472 -614 1582 -604
rect 530 -696 1472 -654
rect 358 -726 530 -716
rect 7434 -624 8704 -590
rect 8102 -628 8704 -624
rect 5424 -646 5516 -636
rect 3810 -656 3886 -646
rect 3886 -704 5424 -666
rect 3810 -722 3886 -712
rect 8244 -638 8338 -628
rect 7462 -668 7504 -666
rect 5424 -726 5516 -716
rect 6588 -682 6668 -672
rect -1116 -744 -1002 -734
rect 1472 -738 1582 -728
rect 6588 -762 6668 -752
rect 7424 -678 7544 -668
rect 7932 -672 8018 -662
rect 7544 -736 7932 -694
rect 7424 -760 7544 -750
rect -1116 -814 -1002 -804
rect -1090 -1342 -1052 -814
rect 640 -1302 786 -1292
rect -1090 -1372 640 -1342
rect 640 -1410 786 -1400
rect 4974 -1344 5064 -1334
rect 230 -1444 300 -1434
rect 1790 -1446 1852 -1436
rect 300 -1514 1790 -1480
rect 300 -1516 1852 -1514
rect 1790 -1524 1852 -1516
rect 3616 -1448 3676 -1438
rect 6602 -1374 6646 -762
rect 7932 -768 8018 -758
rect 8244 -784 8338 -774
rect 8638 -960 8814 -950
rect 8638 -1126 8814 -1116
rect 5064 -1416 6646 -1374
rect 6602 -1420 6646 -1416
rect 4974 -1462 5064 -1452
rect 3616 -1530 3676 -1520
rect 230 -1542 300 -1532
rect 3634 -1574 3664 -1530
rect 5380 -1558 5484 -1548
rect 3634 -1614 5380 -1574
rect 5380 -1638 5484 -1628
rect 8686 -1708 8730 -1126
rect 6818 -1712 8732 -1708
rect 2372 -1718 8732 -1712
rect -1540 -1778 8732 -1718
rect -1540 -1794 7014 -1778
rect -1540 -1800 3102 -1794
<< via2 >>
rect 7938 -332 8014 -268
rect 7932 -758 8018 -672
<< metal3 >>
rect 7928 -268 8024 -263
rect 7928 -332 7938 -268
rect 8014 -332 8024 -268
rect 7928 -337 8024 -332
rect 7944 -667 8008 -337
rect 7922 -672 8028 -667
rect 7922 -758 7932 -672
rect 8018 -758 8028 -672
rect 7922 -763 8028 -758
<< labels >>
flabel poly 3270 -518 3270 -518 0 FreeSans 800 0 0 0 vinp
flabel poly 3074 -1576 3074 -1576 0 FreeSans 800 0 0 0 vref
flabel poly 3016 820 3016 820 0 FreeSans 800 0 0 0 clk
flabel metal1 4010 -1810 4010 -1810 0 FreeSans 800 0 0 0 vssa
flabel metal1 2572 1128 2572 1128 0 FreeSans 800 0 0 0 vdda
flabel locali 6904 -200 6904 -200 0 FreeSans 800 0 0 0 vom
flabel locali -1380 -296 -1380 -296 0 FreeSans 800 0 0 0 vop
flabel metal1 7478 -894 7478 -894 0 FreeSans 800 0 0 0 vp
flabel metal1 8284 -1046 8284 -1046 0 FreeSans 800 0 0 0 vm
flabel metal1 2418 -988 2418 -988 0 FreeSans 800 0 0 0 nmos8point5_0/d
flabel metal1 2734 -1450 2734 -1450 0 FreeSans 800 0 0 0 nmos8point5_0/s
rlabel comment 8272 -526 8272 -526 4 sky130_fd_sc_hvl__inv_1_3/inv_1
flabel metal1 8272 -475 8560 -401 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_3/VGND
flabel metal1 8272 -526 8560 -503 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_3/VNB
flabel metal1 8272 163 8560 237 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_3/VPWR
flabel metal1 8272 265 8560 288 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_3/VPB
flabel locali 8303 -210 8337 -176 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_3/A
flabel locali 8399 -210 8433 -176 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_3/A
flabel locali 8495 -358 8529 -324 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_3/Y
flabel locali 8495 -284 8529 -250 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_3/Y
flabel locali 8495 -210 8529 -176 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_3/Y
flabel locali 8495 -136 8529 -102 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_3/Y
flabel locali 8495 -62 8529 -28 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_3/Y
flabel locali 8495 12 8529 46 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_3/Y
flabel locali 8495 86 8529 120 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_3/Y
rlabel comment 7452 -522 7452 -522 4 sky130_fd_sc_hvl__inv_1_2/inv_1
flabel metal1 7452 -471 7740 -397 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_2/VGND
flabel metal1 7452 -522 7740 -499 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_2/VNB
flabel metal1 7452 167 7740 241 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_2/VPWR
flabel metal1 7452 269 7740 292 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_2/VPB
flabel locali 7483 -206 7517 -172 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_2/A
flabel locali 7579 -206 7613 -172 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_2/A
flabel locali 7675 -354 7709 -320 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_2/Y
flabel locali 7675 -280 7709 -246 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_2/Y
flabel locali 7675 -206 7709 -172 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_2/Y
flabel locali 7675 -132 7709 -98 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_2/Y
flabel locali 7675 -58 7709 -24 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_2/Y
flabel locali 7675 16 7709 50 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_2/Y
flabel locali 7675 90 7709 124 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_2/Y
rlabel comment -1076 -630 -1076 -630 6 sky130_fd_sc_hvl__inv_1_1/inv_1
flabel metal1 -1364 -579 -1076 -505 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_1/VGND
flabel metal1 -1364 -630 -1076 -607 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_1/VNB
flabel metal1 -1364 59 -1076 133 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_1/VPWR
flabel metal1 -1364 161 -1076 184 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_1/VPB
flabel locali -1141 -314 -1107 -280 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_1/A
flabel locali -1237 -314 -1203 -280 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_1/A
flabel locali -1333 -462 -1299 -428 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_1/Y
flabel locali -1333 -388 -1299 -354 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_1/Y
flabel locali -1333 -314 -1299 -280 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_1/Y
flabel locali -1333 -240 -1299 -206 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_1/Y
flabel locali -1333 -166 -1299 -132 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_1/Y
flabel locali -1333 -92 -1299 -58 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_1/Y
flabel locali -1333 -18 -1299 16 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_1/Y
rlabel comment 6614 -540 6614 -540 4 sky130_fd_sc_hvl__inv_1_0/inv_1
flabel metal1 6614 -489 6902 -415 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_0/VGND
flabel metal1 6614 -540 6902 -517 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_0/VNB
flabel metal1 6614 149 6902 223 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_0/VPWR
flabel metal1 6614 251 6902 274 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_0/VPB
flabel locali 6645 -224 6679 -190 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_0/A
flabel locali 6741 -224 6775 -190 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_0/A
flabel locali 6837 -372 6871 -338 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_0/Y
flabel locali 6837 -298 6871 -264 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_0/Y
flabel locali 6837 -224 6871 -190 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_0/Y
flabel locali 6837 -150 6871 -116 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_0/Y
flabel locali 6837 -76 6871 -42 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_0/Y
flabel locali 6837 -2 6871 32 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_0/Y
flabel locali 6837 72 6871 106 0 FreeSans 340 0 0 0 sky130_fd_sc_hvl__inv_1_0/Y
<< end >>
