magic
tech sky130A
magscale 1 2
timestamp 1634904824
<< metal1 >>
rect 98 3002 1190 3008
rect 96 2998 1190 3002
rect 96 2962 1198 2998
rect 96 2864 152 2962
rect 620 2868 676 2962
rect 1142 2872 1198 2962
rect 96 228 162 2864
rect 360 220 426 2856
rect 618 232 684 2868
rect 882 236 948 2872
rect 1138 236 1204 2872
rect 366 148 422 220
rect 886 148 942 236
rect 356 108 942 148
use sky130_fd_pr__pfet_g5v0d10v5_TV7D4F  sky130_fd_pr__pfet_g5v0d10v5_TV7D4F_0
timestamp 1634904824
transform 1 0 650 0 1 1554
box -745 -1649 745 1649
<< end >>
