magic
tech sky130A
timestamp 1634018273
<< pwell >>
rect -391 -238 17607 12033
use nmos5555  nmos5555_0
timestamp 1634016467
transform 1 0 376 0 1 69
box -376 -69 3019 2828
use nmos5555  nmos5555_1
timestamp 1634016467
transform 1 0 375 0 1 3025
box -376 -69 3019 2828
use nmos5555  nmos5555_5
timestamp 1634016467
transform 1 0 3879 0 1 63
box -376 -69 3019 2828
use nmos5555  nmos5555_8
timestamp 1634016467
transform 1 0 3877 0 1 3025
box -376 -69 3019 2828
use nmos5555  nmos5555_6
timestamp 1634016467
transform 1 0 7386 0 1 63
box -376 -69 3019 2828
use nmos5555  nmos5555_9
timestamp 1634016467
transform 1 0 7386 0 1 3025
box -376 -69 3019 2828
use nmos5555  nmos5555_10
timestamp 1634016467
transform 1 0 10839 0 1 3026
box -376 -69 3019 2828
use nmos5555  nmos5555_7
timestamp 1634016467
transform 1 0 10840 0 1 68
box -376 -69 3019 2828
use nmos5555  nmos5555_14
timestamp 1634016467
transform 1 0 3875 0 1 8979
box -376 -69 3019 2828
use nmos5555  nmos5555_11
timestamp 1634016467
transform 1 0 3877 0 1 5998
box -376 -69 3019 2828
use nmos5555  nmos5555_2
timestamp 1634016467
transform 1 0 374 0 1 5997
box -376 -69 3019 2828
use nmos5555  nmos5555_3
timestamp 1634016467
transform 1 0 374 0 1 8977
box -376 -69 3019 2828
use nmos5555  nmos5555_15
timestamp 1634016467
transform 1 0 7385 0 1 8981
box -376 -69 3019 2828
use nmos5555  nmos5555_12
timestamp 1634016467
transform 1 0 7386 0 1 5998
box -376 -69 3019 2828
use nmos5555  nmos5555_16
timestamp 1634016467
transform 1 0 10836 0 1 8980
box -376 -69 3019 2828
use nmos5555  nmos5555_13
timestamp 1634016467
transform 1 0 10837 0 1 5998
box -376 -69 3019 2828
use nmos5555  nmos5555_19
timestamp 1634016467
transform 1 0 14301 0 1 8977
box -376 -69 3019 2828
use nmos5555  nmos5555_18
timestamp 1634016467
transform 1 0 14301 0 1 6013
box -376 -69 3019 2828
use nmos5555  nmos5555_17
timestamp 1634016467
transform 1 0 14306 0 1 3027
box -376 -69 3019 2828
use nmos5555  nmos5555_4
timestamp 1634016467
transform 1 0 14306 0 1 69
box -376 -69 3019 2828
<< end >>
