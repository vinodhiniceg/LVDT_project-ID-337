magic
tech sky130A
magscale 1 2
timestamp 1634617818
<< mvnmos >>
rect -287 -100 -187 100
rect -129 -100 -29 100
rect 29 -100 129 100
rect 187 -100 287 100
<< mvndiff >>
rect -345 26 -287 100
rect -345 -26 -333 26
rect -299 -26 -287 26
rect -345 -100 -287 -26
rect -187 26 -129 100
rect -187 -26 -175 26
rect -141 -26 -129 26
rect -187 -100 -129 -26
rect -29 26 29 100
rect -29 -26 -17 26
rect 17 -26 29 26
rect -29 -100 29 -26
rect 129 26 187 100
rect 129 -26 141 26
rect 175 -26 187 26
rect 129 -100 187 -26
rect 287 26 345 100
rect 287 -26 299 26
rect 333 -26 345 26
rect 287 -100 345 -26
<< mvndiffc >>
rect -333 -26 -299 26
rect -175 -26 -141 26
rect -17 -26 17 26
rect 141 -26 175 26
rect 299 -26 333 26
<< poly >>
rect -287 100 -187 126
rect -129 100 -29 126
rect 29 100 129 126
rect 187 100 287 126
rect -287 -126 -187 -100
rect -129 -126 -29 -100
rect 29 -126 129 -100
rect 187 -126 287 -100
<< locali >>
rect -333 26 -299 42
rect -333 -42 -299 -26
rect -175 26 -141 42
rect -175 -42 -141 -26
rect -17 26 17 42
rect -17 -42 17 -26
rect 141 26 175 42
rect 141 -42 175 -26
rect 299 26 333 42
rect 299 -42 333 -26
<< viali >>
rect -333 -26 -299 26
rect -175 -26 -141 26
rect -17 -26 17 26
rect 141 -26 175 26
rect 299 -26 333 26
<< metal1 >>
rect -339 26 -293 38
rect -339 -26 -333 26
rect -299 -26 -293 26
rect -339 -38 -293 -26
rect -181 26 -135 38
rect -181 -26 -175 26
rect -141 -26 -135 26
rect -181 -38 -135 -26
rect -23 26 23 38
rect -23 -26 -17 26
rect 17 -26 23 26
rect -23 -38 23 -26
rect 135 26 181 38
rect 135 -26 141 26
rect 175 -26 181 26
rect 135 -38 181 -26
rect 293 26 339 38
rect 293 -26 299 26
rect 333 -26 339 26
rect 293 -38 339 -26
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string parameters w 1 l 0.5 m 1 nf 4 diffcov 30 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 30 viadrn 30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
