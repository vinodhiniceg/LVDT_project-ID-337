magic
tech sky130A
timestamp 1634044821
<< mvnmos >>
rect -2558 547 -1558 1547
rect -1529 547 -529 1547
rect -500 547 500 1547
rect 529 547 1529 1547
rect 1558 547 2558 1547
rect -2558 -500 -1558 500
rect -1529 -500 -529 500
rect -500 -500 500 500
rect 529 -500 1529 500
rect 1558 -500 2558 500
rect -2558 -1547 -1558 -547
rect -1529 -1547 -529 -547
rect -500 -1547 500 -547
rect 529 -1547 1529 -547
rect 1558 -1547 2558 -547
<< mvndiff >>
rect -2587 1195 -2558 1547
rect -2587 899 -2581 1195
rect -2564 899 -2558 1195
rect -2587 547 -2558 899
rect -1558 1195 -1529 1547
rect -1558 899 -1552 1195
rect -1535 899 -1529 1195
rect -1558 547 -1529 899
rect -529 1195 -500 1547
rect -529 899 -523 1195
rect -506 899 -500 1195
rect -529 547 -500 899
rect 500 1195 529 1547
rect 500 899 506 1195
rect 523 899 529 1195
rect 500 547 529 899
rect 1529 1195 1558 1547
rect 1529 899 1535 1195
rect 1552 899 1558 1195
rect 1529 547 1558 899
rect 2558 1195 2587 1547
rect 2558 899 2564 1195
rect 2581 899 2587 1195
rect 2558 547 2587 899
rect -2587 148 -2558 500
rect -2587 -148 -2581 148
rect -2564 -148 -2558 148
rect -2587 -500 -2558 -148
rect -1558 148 -1529 500
rect -1558 -148 -1552 148
rect -1535 -148 -1529 148
rect -1558 -500 -1529 -148
rect -529 148 -500 500
rect -529 -148 -523 148
rect -506 -148 -500 148
rect -529 -500 -500 -148
rect 500 148 529 500
rect 500 -148 506 148
rect 523 -148 529 148
rect 500 -500 529 -148
rect 1529 148 1558 500
rect 1529 -148 1535 148
rect 1552 -148 1558 148
rect 1529 -500 1558 -148
rect 2558 148 2587 500
rect 2558 -148 2564 148
rect 2581 -148 2587 148
rect 2558 -500 2587 -148
rect -2587 -899 -2558 -547
rect -2587 -1195 -2581 -899
rect -2564 -1195 -2558 -899
rect -2587 -1547 -2558 -1195
rect -1558 -899 -1529 -547
rect -1558 -1195 -1552 -899
rect -1535 -1195 -1529 -899
rect -1558 -1547 -1529 -1195
rect -529 -899 -500 -547
rect -529 -1195 -523 -899
rect -506 -1195 -500 -899
rect -529 -1547 -500 -1195
rect 500 -899 529 -547
rect 500 -1195 506 -899
rect 523 -1195 529 -899
rect 500 -1547 529 -1195
rect 1529 -899 1558 -547
rect 1529 -1195 1535 -899
rect 1552 -1195 1558 -899
rect 1529 -1547 1558 -1195
rect 2558 -899 2587 -547
rect 2558 -1195 2564 -899
rect 2581 -1195 2587 -899
rect 2558 -1547 2587 -1195
<< mvndiffc >>
rect -2581 899 -2564 1195
rect -1552 899 -1535 1195
rect -523 899 -506 1195
rect 506 899 523 1195
rect 1535 899 1552 1195
rect 2564 899 2581 1195
rect -2581 -148 -2564 148
rect -1552 -148 -1535 148
rect -523 -148 -506 148
rect 506 -148 523 148
rect 1535 -148 1552 148
rect 2564 -148 2581 148
rect -2581 -1195 -2564 -899
rect -1552 -1195 -1535 -899
rect -523 -1195 -506 -899
rect 506 -1195 523 -899
rect 1535 -1195 1552 -899
rect 2564 -1195 2581 -899
<< poly >>
rect -2558 1547 -1558 1560
rect -1529 1547 -529 1560
rect -500 1547 500 1560
rect 529 1547 1529 1560
rect 1558 1547 2558 1560
rect -2558 534 -1558 547
rect -1529 534 -529 547
rect -500 534 500 547
rect 529 534 1529 547
rect 1558 534 2558 547
rect -2558 500 -1558 513
rect -1529 500 -529 513
rect -500 500 500 513
rect 529 500 1529 513
rect 1558 500 2558 513
rect -2558 -513 -1558 -500
rect -1529 -513 -529 -500
rect -500 -513 500 -500
rect 529 -513 1529 -500
rect 1558 -513 2558 -500
rect -2558 -547 -1558 -534
rect -1529 -547 -529 -534
rect -500 -547 500 -534
rect 529 -547 1529 -534
rect 1558 -547 2558 -534
rect -2558 -1560 -1558 -1547
rect -1529 -1560 -529 -1547
rect -500 -1560 500 -1547
rect 529 -1560 1529 -1547
rect 1558 -1560 2558 -1547
<< locali >>
rect -2581 1195 -2564 1203
rect -2581 891 -2564 899
rect -1552 1195 -1535 1203
rect -1552 891 -1535 899
rect -523 1195 -506 1203
rect -523 891 -506 899
rect 506 1195 523 1203
rect 506 891 523 899
rect 1535 1195 1552 1203
rect 1535 891 1552 899
rect 2564 1195 2581 1203
rect 2564 891 2581 899
rect -2581 148 -2564 156
rect -2581 -156 -2564 -148
rect -1552 148 -1535 156
rect -1552 -156 -1535 -148
rect -523 148 -506 156
rect -523 -156 -506 -148
rect 506 148 523 156
rect 506 -156 523 -148
rect 1535 148 1552 156
rect 1535 -156 1552 -148
rect 2564 148 2581 156
rect 2564 -156 2581 -148
rect -2581 -899 -2564 -891
rect -2581 -1203 -2564 -1195
rect -1552 -899 -1535 -891
rect -1552 -1203 -1535 -1195
rect -523 -899 -506 -891
rect -523 -1203 -506 -1195
rect 506 -899 523 -891
rect 506 -1203 523 -1195
rect 1535 -899 1552 -891
rect 1535 -1203 1552 -1195
rect 2564 -899 2581 -891
rect 2564 -1203 2581 -1195
<< viali >>
rect -2581 899 -2564 1195
rect -1552 899 -1535 1195
rect -523 899 -506 1195
rect 506 899 523 1195
rect 1535 899 1552 1195
rect 2564 899 2581 1195
rect -2581 -148 -2564 148
rect -1552 -148 -1535 148
rect -523 -148 -506 148
rect 506 -148 523 148
rect 1535 -148 1552 148
rect 2564 -148 2581 148
rect -2581 -1195 -2564 -899
rect -1552 -1195 -1535 -899
rect -523 -1195 -506 -899
rect 506 -1195 523 -899
rect 1535 -1195 1552 -899
rect 2564 -1195 2581 -899
<< metal1 >>
rect -2584 1195 -2561 1201
rect -2584 899 -2581 1195
rect -2564 899 -2561 1195
rect -2584 893 -2561 899
rect -1555 1195 -1532 1201
rect -1555 899 -1552 1195
rect -1535 899 -1532 1195
rect -1555 893 -1532 899
rect -526 1195 -503 1201
rect -526 899 -523 1195
rect -506 899 -503 1195
rect -526 893 -503 899
rect 503 1195 526 1201
rect 503 899 506 1195
rect 523 899 526 1195
rect 503 893 526 899
rect 1532 1195 1555 1201
rect 1532 899 1535 1195
rect 1552 899 1555 1195
rect 1532 893 1555 899
rect 2561 1195 2584 1201
rect 2561 899 2564 1195
rect 2581 899 2584 1195
rect 2561 893 2584 899
rect -2584 148 -2561 154
rect -2584 -148 -2581 148
rect -2564 -148 -2561 148
rect -2584 -154 -2561 -148
rect -1555 148 -1532 154
rect -1555 -148 -1552 148
rect -1535 -148 -1532 148
rect -1555 -154 -1532 -148
rect -526 148 -503 154
rect -526 -148 -523 148
rect -506 -148 -503 148
rect -526 -154 -503 -148
rect 503 148 526 154
rect 503 -148 506 148
rect 523 -148 526 148
rect 503 -154 526 -148
rect 1532 148 1555 154
rect 1532 -148 1535 148
rect 1552 -148 1555 148
rect 1532 -154 1555 -148
rect 2561 148 2584 154
rect 2561 -148 2564 148
rect 2581 -148 2584 148
rect 2561 -154 2584 -148
rect -2584 -899 -2561 -893
rect -2584 -1195 -2581 -899
rect -2564 -1195 -2561 -899
rect -2584 -1201 -2561 -1195
rect -1555 -899 -1532 -893
rect -1555 -1195 -1552 -899
rect -1535 -1195 -1532 -899
rect -1555 -1201 -1532 -1195
rect -526 -899 -503 -893
rect -526 -1195 -523 -899
rect -506 -1195 -503 -899
rect -526 -1201 -503 -1195
rect 503 -899 526 -893
rect 503 -1195 506 -899
rect 523 -1195 526 -899
rect 503 -1201 526 -1195
rect 1532 -899 1555 -893
rect 1532 -1195 1535 -899
rect 1552 -1195 1555 -899
rect 1532 -1201 1555 -1195
rect 2561 -899 2584 -893
rect 2561 -1195 2564 -899
rect 2581 -1195 2584 -899
rect 2561 -1201 2584 -1195
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string parameters w 10 l 10 m 3 nf 5 diffcov 30 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 30 viadrn 30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
