magic
tech sky130A
magscale 1 2
timestamp 1634365921
<< error_p >>
rect -70 -2600 -10 2600
rect 10 -2600 70 2600
<< metal3 >>
rect -4309 2572 -10 2600
rect -4309 -2572 -94 2572
rect -30 -2572 -10 2572
rect -4309 -2600 -10 -2572
rect 10 2572 4309 2600
rect 10 -2572 4225 2572
rect 4289 -2572 4309 2572
rect 10 -2600 4309 -2572
<< via3 >>
rect -94 -2572 -30 2572
rect 4225 -2572 4289 2572
<< mimcap >>
rect -4209 2460 -209 2500
rect -4209 -2460 -4169 2460
rect -249 -2460 -209 2460
rect -4209 -2500 -209 -2460
rect 110 2460 4110 2500
rect 110 -2460 150 2460
rect 4070 -2460 4110 2460
rect 110 -2500 4110 -2460
<< mimcapcontact >>
rect -4169 -2460 -249 2460
rect 150 -2460 4070 2460
<< metal4 >>
rect -110 2572 -14 2588
rect -4170 2460 -248 2461
rect -4170 -2460 -4169 2460
rect -249 -2460 -248 2460
rect -4170 -2461 -248 -2460
rect -110 -2572 -94 2572
rect -30 -2572 -14 2572
rect 4209 2572 4305 2588
rect 149 2460 4071 2461
rect 149 -2460 150 2460
rect 4070 -2460 4071 2460
rect 149 -2461 4071 -2460
rect -110 -2588 -14 -2572
rect 4209 -2572 4225 2572
rect 4289 -2572 4305 2572
rect 4209 -2588 4305 -2572
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX 10 -2600 4210 2600
string parameters w 20.00 l 25.00 val 1.017k carea 2.00 cperi 0.19 nx 2 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>
