magic
tech sky130A
magscale 1 2
timestamp 1634128943
<< pwell >>
rect -56 7558 8420 7632
rect -160 7313 8568 7558
rect -160 7308 6787 7313
rect 7017 7308 8568 7313
rect -160 7290 8568 7308
rect -160 7284 1582 7290
rect -160 7270 1222 7284
rect -160 7258 1206 7270
rect 1650 7260 8568 7290
rect -160 7118 1200 7258
rect 1650 7166 3128 7260
rect 1650 7146 1736 7166
rect -160 7086 1206 7118
rect 1614 7086 1736 7146
rect -160 7084 1306 7086
rect 1512 7084 1736 7086
rect 2100 7084 3128 7166
rect -160 7026 422 7084
rect 2508 7048 3128 7084
rect 3356 7052 8568 7260
rect 3356 7048 5074 7052
rect 2508 7026 5074 7048
rect -160 6836 5074 7026
rect 5248 6836 8568 7052
rect -160 -374 8568 6836
<< mvpsubdiff >>
rect -56 7454 8420 7632
rect -56 7313 8436 7454
rect -56 7308 6787 7313
rect 7017 7308 8436 7313
rect -56 24 298 7308
rect 8082 24 8436 7308
rect -56 -270 8464 24
rect -12 -300 8464 -270
<< poly >>
rect 2262 7216 2420 7242
rect 2262 7154 2290 7216
rect 2396 7154 2420 7216
rect 2262 7134 2420 7154
rect 3934 7138 4494 7278
rect 6720 7266 7094 7288
rect 6720 7178 6834 7266
rect 6970 7178 7094 7266
rect 6720 7146 7094 7178
<< polycont >>
rect 2290 7154 2396 7216
rect 6834 7178 6970 7266
<< locali >>
rect 6812 7266 6988 7278
rect 2274 7216 2412 7230
rect 2274 7154 2290 7216
rect 2396 7154 2412 7216
rect 2274 7140 2412 7154
rect 2300 7026 2372 7140
rect 3176 7048 3244 7226
rect 6812 7178 6834 7266
rect 6970 7178 6988 7266
rect 6812 7168 6988 7178
rect 1350 7004 1432 7026
rect 1850 6988 2472 7026
rect 3176 6992 3276 7048
rect 6840 7026 6940 7168
rect 7816 7026 7876 7028
rect 2422 6926 2472 6988
rect 2422 6856 2844 6926
rect 5156 6822 5238 7020
rect 6840 6960 7876 7026
rect 7816 6854 7876 6960
rect 5534 2826 5876 2910
<< viali >>
rect 2306 7164 2378 7206
rect 6856 7190 6944 7254
<< metal1 >>
rect 6812 7254 6988 7278
rect 2274 7206 2412 7230
rect 2274 7164 2306 7206
rect 2378 7164 2412 7206
rect 6812 7190 6856 7254
rect 6944 7190 6988 7254
rect 6812 7168 6988 7190
rect 2274 7140 2412 7164
use nmos33310  nmos33310_2
timestamp 1634127866
transform 1 0 5842 0 1 216
box -444 -236 2354 7116
use nmos33310  nmos33310_1
timestamp 1634127866
transform 1 0 3188 0 1 230
box -444 -236 2354 7116
use nmos33310  nmos33310_0
timestamp 1634127866
transform 1 0 444 0 1 236
box -444 -236 2354 7116
<< labels >>
flabel pwell 2820 6956 2820 6956 0 FreeSans 1600 0 0 0 sub
flabel poly 4160 7200 4160 7200 0 FreeSans 1600 0 0 0 g
flabel locali 3210 7160 3210 7160 0 FreeSans 1600 0 0 0 s
flabel locali 5194 6942 5194 6942 0 FreeSans 1600 0 0 0 d
<< end >>
