magic
tech sky130A
magscale 1 2
timestamp 1634272161
<< nwell >>
rect -266 3580 2936 3588
rect -450 -184 2936 3580
rect -450 -192 -180 -184
<< mvnsubdiff >>
rect -250 3164 -34 3224
rect -250 418 -220 3164
rect -80 418 -34 3164
rect -250 364 -34 418
<< mvnsubdiffcont >>
rect -220 418 -80 3164
<< poly >>
rect 440 3460 2530 3530
rect 154 2760 578 2828
rect 892 2754 1316 2822
rect 1474 2760 1898 2828
rect 2146 2760 2570 2828
rect 148 2064 572 2132
rect 860 2064 1284 2132
rect 1470 2062 1894 2130
rect 2186 2060 2610 2128
rect 134 1366 558 1434
rect 880 1372 1304 1440
rect 1508 1366 1932 1434
rect 2144 1372 2568 1440
rect 130 676 554 744
rect 910 676 1334 744
rect 1460 670 1884 738
rect 2178 674 2602 742
<< locali >>
rect 2670 3380 2848 3390
rect 34 3372 90 3378
rect 2662 3372 2848 3380
rect 30 3330 2848 3372
rect -250 3164 -34 3224
rect -250 418 -220 3164
rect -80 418 -34 3164
rect -250 364 -34 418
rect 34 376 90 3330
rect 696 408 752 3208
rect 1352 3204 1408 3330
rect 686 364 752 408
rect 1350 3172 1408 3204
rect 2662 3320 2848 3330
rect 686 166 746 364
rect 1350 360 1406 3172
rect 2010 406 2066 3162
rect 2662 3142 2738 3320
rect 2010 318 2074 406
rect 2664 322 2720 3142
rect 2014 170 2074 318
rect 2014 166 2172 170
rect 686 104 2172 166
rect 686 98 746 104
rect 2014 96 2074 104
<< viali >>
rect -196 510 -112 3078
<< metal1 >>
rect -250 3078 -34 3224
rect -250 510 -196 3078
rect -112 510 -34 3078
rect -250 364 -34 510
use sky130_fd_pr__pfet_g5v0d10v5_6CSA4Z  sky130_fd_pr__pfet_g5v0d10v5_6CSA4Z_0
timestamp 1634272161
transform 1 0 1381 0 1 1750
box -1411 -1754 1411 1754
<< labels >>
flabel locali 2784 3354 2784 3354 0 FreeSans 1600 0 0 0 s
flabel locali 2116 134 2116 134 0 FreeSans 1600 0 0 0 d
flabel poly 1116 3484 1116 3484 0 FreeSans 1600 0 0 0 g
<< end >>
