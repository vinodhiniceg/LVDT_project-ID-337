`timescale 1us / 1ns

module adc_logic(
    a,
    y
);

input [4:0] a;
output [4:0] y;

wire [4:0] a;
wire [4:0] y;

// Y0 = A4'*A1*A0 (A3*A2 + A3'*A2')
assign y[0] = ( (~a[4]) & a[1] & a[0] ) & ( (a[3] & a[2]) | ((~a[3]) & (~a[2])) );

// Y1 = A4*A3*A2*A1*A0 + A4'*A3'*A2' (A1*A0 + A1'*A0)
assign y[1] = (a[0] & a[1] & a[2] & a[3] & a[4]) | (( (~a[4]) & (~a[3]) & (~a[2]) ) & ( (a[1] & a[0]) | ((~a[1]) & a[0]) ));

// Y2 = A4'*A3'*A2' (A1*A0 + A1'*A0)
assign y[2] = ( (~a[4]) & (~a[3]) & (~a[2]) ) & ( (a[1] & a[0]) | ((~a[1]) & a[0]) );

// Y3 = A4'*A3'*A2' (A1*A0 + A1'*A0)
assign y[3] = ( (~a[4]) & (~a[3]) & (~a[2]) ) & ( (a[1] & a[0]) | ((~a[1]) & a[0]) );

// Y4 = A4'*A3'*A2' (A1*A0 + A1'*A0)
assign y[4] = ( (~a[4]) & (~a[3]) & (~a[2]) ) & ( (a[1] & a[0]) | ((~a[1]) & a[0]) );


endmodule