magic
tech sky130A
timestamp 1634132563
<< error_s >>
rect 1645 1401 1674 1701
rect 1645 1054 1674 1354
rect 1645 707 1674 1007
rect 1645 360 1674 660
rect 1645 13 1674 313
<< mvpsubdiff >>
rect -174 1355 -68 1390
rect -174 478 -158 1355
rect -84 478 -68 1355
rect -174 435 -68 478
<< mvpsubdiffcont >>
rect -158 478 -84 1355
<< poly >>
rect 182 1711 1596 1760
rect 85 1359 247 1392
rect 418 1362 580 1395
rect 744 1362 906 1395
rect 1099 1362 1261 1395
rect 1390 1362 1552 1395
rect 88 1014 250 1047
rect 399 1014 561 1047
rect 711 1010 873 1043
rect 1087 1012 1249 1045
rect 1372 1013 1534 1046
rect 86 669 248 702
rect 432 670 594 703
rect 747 666 909 699
rect 1091 669 1253 702
rect 1431 664 1593 697
rect 75 322 237 355
rect 409 320 571 353
rect 751 317 913 350
rect 1100 321 1262 354
rect 1413 318 1575 351
<< locali >>
rect 1 1682 32 1687
rect -9 1674 32 1682
rect 660 1676 691 1678
rect 656 1674 691 1676
rect 1307 1674 1354 1676
rect -9 1636 1354 1674
rect -9 1522 32 1636
rect -174 1355 -68 1390
rect -174 478 -158 1355
rect -84 478 -68 1355
rect -174 435 -68 478
rect 1 173 30 1522
rect 330 175 359 1558
rect 656 1516 691 1636
rect 656 175 685 1516
rect 987 193 1016 1576
rect 1307 1485 1354 1636
rect 1314 177 1343 1485
rect 1646 176 1675 1547
rect 331 76 358 175
rect 990 76 1017 174
rect 1644 164 1675 176
rect 1644 76 1671 164
rect 323 27 1675 76
rect 990 25 1017 27
<< viali >>
rect -151 554 -104 1306
<< metal1 >>
rect -174 1306 -68 1390
rect -174 554 -151 1306
rect -104 554 -68 1306
rect -174 435 -68 554
use sky130_fd_pr__nfet_g5v0d10v5_QWH9RS  sky130_fd_pr__nfet_g5v0d10v5_QWH9RS_0
timestamp 1634132563
transform 1 0 837 0 1 857
box -837 -857 837 857
<< end >>
