magic
tech sky130A
magscale 1 2
timestamp 1634908262
<< poly >>
rect 100 4966 444 5088
rect 74 4664 208 4740
rect 350 4672 484 4748
rect 64 4370 198 4446
rect 330 4366 464 4442
rect 68 4072 202 4148
rect 348 4074 482 4150
rect 84 3788 218 3864
rect 350 3780 484 3856
rect 78 3490 212 3566
rect 348 3488 482 3564
rect 78 3194 212 3270
rect 328 3196 462 3272
rect 72 2900 206 2976
rect 326 2904 460 2980
rect 90 2608 224 2684
rect 346 2612 480 2688
rect 84 2312 218 2388
rect 316 2314 450 2390
rect 70 2026 204 2102
rect 358 2024 492 2100
rect 58 1726 192 1802
rect 330 1724 464 1800
rect 76 1440 210 1516
rect 338 1434 472 1510
rect 90 1140 224 1216
rect 336 1142 470 1218
rect 74 852 208 928
rect 350 848 484 924
rect 62 558 196 634
rect 356 550 490 626
rect 66 250 200 326
rect 334 252 468 328
<< metal1 >>
rect -10 130 40 4852
rect 254 146 304 4868
rect 504 144 554 4866
use sky130_fd_pr__nfet_g5v0d10v5_U3KEUB  sky130_fd_pr__nfet_g5v0d10v5_U3KEUB_0
timestamp 1634908262
transform 1 0 273 0 1 2498
box -287 -2478 287 2478
<< end >>
