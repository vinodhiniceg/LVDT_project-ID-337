magic
tech sky130A
timestamp 1634123280
<< nwell >>
rect -137 -172 3296 10404
<< poly >>
rect 461 9139 529 9473
rect 674 9137 742 9471
rect 1010 9141 1078 9475
rect 1351 9143 1419 9477
rect 1662 9141 1730 9475
rect 2015 9141 2083 9475
rect 2322 9135 2390 9469
rect 2694 9146 2762 9480
rect 467 7826 546 8130
rect 680 7830 759 8134
rect 1034 7826 1113 8130
rect 1368 7828 1447 8132
rect 1698 7832 1777 8136
rect 2030 7828 2109 8132
rect 2332 7824 2411 8128
rect 2735 7828 2807 8128
rect 467 6501 556 6821
rect 670 6495 759 6815
rect 1006 6501 1095 6821
rect 1319 6508 1408 6828
rect 1687 6495 1776 6815
rect 1992 6501 2081 6821
rect 2326 6504 2415 6824
rect 2741 6501 2830 6821
rect 357 5193 446 5487
rect 282 5167 481 5193
rect 685 5171 774 5491
rect 1014 5173 1103 5493
rect 1323 5167 1412 5487
rect 1672 5179 1761 5499
rect 1987 5173 2076 5493
rect 2311 5167 2400 5487
rect 2730 5165 2819 5485
rect 458 3868 543 4166
rect 326 3856 543 3868
rect 326 3847 511 3856
rect 708 3854 793 4164
rect 1042 3842 1131 4162
rect 1353 3847 1442 4167
rect 1619 3845 1708 4165
rect 1990 3853 2079 4173
rect 2305 3849 2394 4169
rect 2730 3849 2819 4169
rect 478 2514 550 2838
rect 725 2514 797 2838
rect 1034 2514 1106 2838
rect 1358 2515 1430 2839
rect 1671 2517 1743 2841
rect 2023 2520 2095 2844
rect 2305 2517 2377 2841
rect 2747 2512 2819 2836
rect 477 1186 549 1510
rect 677 1186 749 1510
rect 1050 1183 1122 1507
rect 1403 1177 1475 1501
rect 1692 1186 1764 1510
rect 1979 1184 2051 1508
rect 2291 1181 2363 1505
rect 2734 1175 2806 1499
<< locali >>
rect 200 991 285 10075
rect 2485 9338 2569 9511
rect 2523 8085 2602 8328
rect 2540 6734 2599 7041
rect 2527 5434 2586 5771
rect 2523 4088 2586 4222
rect 2531 2775 2586 2897
rect 2536 1449 2607 1563
<< viali >>
rect 2460 9233 2633 9338
rect 2506 7958 2641 8085
rect 2477 6650 2691 6734
rect 2493 5325 2712 5434
rect 2451 3987 2695 4088
rect 2489 2657 2670 2775
rect 2506 1340 2683 1449
<< metal1 >>
rect 2454 9338 2639 9341
rect 2454 9233 2460 9338
rect 2633 9233 2639 9338
rect 2454 9230 2639 9233
rect 2515 8956 2594 9230
rect 2500 8085 2647 8088
rect 2500 7958 2506 8085
rect 2641 7958 2647 8085
rect 2500 7955 2647 7958
rect 2527 7643 2586 7955
rect 2471 6734 2697 6737
rect 2471 6650 2477 6734
rect 2691 6650 2697 6734
rect 2471 6647 2697 6650
rect 2540 6305 2599 6647
rect 2487 5434 2718 5437
rect 2487 5325 2493 5434
rect 2712 5325 2718 5434
rect 2487 5322 2718 5325
rect 2536 5001 2632 5322
rect 2445 4088 2701 4091
rect 2445 3987 2451 4088
rect 2695 3987 2701 4088
rect 2445 3984 2701 3987
rect 2510 3671 2628 3984
rect 2483 2775 2676 2778
rect 2483 2657 2489 2775
rect 2670 2657 2676 2775
rect 2483 2654 2676 2657
rect 2531 2350 2615 2654
rect 2500 1449 2689 1452
rect 2500 1340 2506 1449
rect 2683 1340 2689 1449
rect 2500 1337 2689 1340
rect 2531 995 2611 1337
use pmos3383  pmos3383_6
timestamp 1634121920
transform 1 0 229 0 1 8103
box -232 -142 2727 1151
use pmos3383  pmos3383_5
timestamp 1634121920
transform 1 0 231 0 1 6790
box -232 -142 2727 1151
use pmos3383  pmos3383_4
timestamp 1634121920
transform 1 0 234 0 1 5463
box -232 -142 2727 1151
use pmos3383  pmos3383_3
timestamp 1634121920
transform 1 0 231 0 1 4136
box -232 -142 2727 1151
use pmos3383  pmos3383_2
timestamp 1634121920
transform 1 0 231 0 1 2813
box -232 -142 2727 1151
use pmos3383  pmos3383_1
timestamp 1634121920
transform 1 0 234 0 1 1476
box -232 -142 2727 1151
use pmos3383  pmos3383_0
timestamp 1634121920
transform 1 0 232 0 1 142
box -232 -142 2727 1151
use pmos3382  pmos3382_0
timestamp 1634120139
transform 1 0 207 0 1 9445
box -213 -180 2742 794
<< end >>
