magic
tech sky130A
magscale 1 2
timestamp 1634046259
<< mvnmos >>
rect -3058 2141 -1058 4141
rect -1000 2141 1000 4141
rect 1058 2141 3058 4141
rect -3058 47 -1058 2047
rect -1000 47 1000 2047
rect 1058 47 3058 2047
rect -3058 -2047 -1058 -47
rect -1000 -2047 1000 -47
rect 1058 -2047 3058 -47
rect -3058 -4141 -1058 -2141
rect -1000 -4141 1000 -2141
rect 1058 -4141 3058 -2141
<< mvndiff >>
rect -3116 3437 -3058 4141
rect -3116 2845 -3104 3437
rect -3070 2845 -3058 3437
rect -3116 2141 -3058 2845
rect -1058 3437 -1000 4141
rect -1058 2845 -1046 3437
rect -1012 2845 -1000 3437
rect -1058 2141 -1000 2845
rect 1000 3437 1058 4141
rect 1000 2845 1012 3437
rect 1046 2845 1058 3437
rect 1000 2141 1058 2845
rect 3058 3437 3116 4141
rect 3058 2845 3070 3437
rect 3104 2845 3116 3437
rect 3058 2141 3116 2845
rect -3116 1343 -3058 2047
rect -3116 751 -3104 1343
rect -3070 751 -3058 1343
rect -3116 47 -3058 751
rect -1058 1343 -1000 2047
rect -1058 751 -1046 1343
rect -1012 751 -1000 1343
rect -1058 47 -1000 751
rect 1000 1343 1058 2047
rect 1000 751 1012 1343
rect 1046 751 1058 1343
rect 1000 47 1058 751
rect 3058 1343 3116 2047
rect 3058 751 3070 1343
rect 3104 751 3116 1343
rect 3058 47 3116 751
rect -3116 -751 -3058 -47
rect -3116 -1343 -3104 -751
rect -3070 -1343 -3058 -751
rect -3116 -2047 -3058 -1343
rect -1058 -751 -1000 -47
rect -1058 -1343 -1046 -751
rect -1012 -1343 -1000 -751
rect -1058 -2047 -1000 -1343
rect 1000 -751 1058 -47
rect 1000 -1343 1012 -751
rect 1046 -1343 1058 -751
rect 1000 -2047 1058 -1343
rect 3058 -751 3116 -47
rect 3058 -1343 3070 -751
rect 3104 -1343 3116 -751
rect 3058 -2047 3116 -1343
rect -3116 -2845 -3058 -2141
rect -3116 -3437 -3104 -2845
rect -3070 -3437 -3058 -2845
rect -3116 -4141 -3058 -3437
rect -1058 -2845 -1000 -2141
rect -1058 -3437 -1046 -2845
rect -1012 -3437 -1000 -2845
rect -1058 -4141 -1000 -3437
rect 1000 -2845 1058 -2141
rect 1000 -3437 1012 -2845
rect 1046 -3437 1058 -2845
rect 1000 -4141 1058 -3437
rect 3058 -2845 3116 -2141
rect 3058 -3437 3070 -2845
rect 3104 -3437 3116 -2845
rect 3058 -4141 3116 -3437
<< mvndiffc >>
rect -3104 2845 -3070 3437
rect -1046 2845 -1012 3437
rect 1012 2845 1046 3437
rect 3070 2845 3104 3437
rect -3104 751 -3070 1343
rect -1046 751 -1012 1343
rect 1012 751 1046 1343
rect 3070 751 3104 1343
rect -3104 -1343 -3070 -751
rect -1046 -1343 -1012 -751
rect 1012 -1343 1046 -751
rect 3070 -1343 3104 -751
rect -3104 -3437 -3070 -2845
rect -1046 -3437 -1012 -2845
rect 1012 -3437 1046 -2845
rect 3070 -3437 3104 -2845
<< poly >>
rect -3058 4141 -1058 4167
rect -1000 4141 1000 4167
rect 1058 4141 3058 4167
rect -3058 2115 -1058 2141
rect -1000 2115 1000 2141
rect 1058 2115 3058 2141
rect -3058 2047 -1058 2073
rect -1000 2047 1000 2073
rect 1058 2047 3058 2073
rect -3058 21 -1058 47
rect -1000 21 1000 47
rect 1058 21 3058 47
rect -3058 -47 -1058 -21
rect -1000 -47 1000 -21
rect 1058 -47 3058 -21
rect -3058 -2073 -1058 -2047
rect -1000 -2073 1000 -2047
rect 1058 -2073 3058 -2047
rect -3058 -2141 -1058 -2115
rect -1000 -2141 1000 -2115
rect 1058 -2141 3058 -2115
rect -3058 -4167 -1058 -4141
rect -1000 -4167 1000 -4141
rect 1058 -4167 3058 -4141
<< locali >>
rect -3104 3437 -3070 3453
rect -3104 2829 -3070 2845
rect -1046 3437 -1012 3453
rect -1046 2829 -1012 2845
rect 1012 3437 1046 3453
rect 1012 2829 1046 2845
rect 3070 3437 3104 3453
rect 3070 2829 3104 2845
rect -3104 1343 -3070 1359
rect -3104 735 -3070 751
rect -1046 1343 -1012 1359
rect -1046 735 -1012 751
rect 1012 1343 1046 1359
rect 1012 735 1046 751
rect 3070 1343 3104 1359
rect 3070 735 3104 751
rect -3104 -751 -3070 -735
rect -3104 -1359 -3070 -1343
rect -1046 -751 -1012 -735
rect -1046 -1359 -1012 -1343
rect 1012 -751 1046 -735
rect 1012 -1359 1046 -1343
rect 3070 -751 3104 -735
rect 3070 -1359 3104 -1343
rect -3104 -2845 -3070 -2829
rect -3104 -3453 -3070 -3437
rect -1046 -2845 -1012 -2829
rect -1046 -3453 -1012 -3437
rect 1012 -2845 1046 -2829
rect 1012 -3453 1046 -3437
rect 3070 -2845 3104 -2829
rect 3070 -3453 3104 -3437
<< viali >>
rect -3104 2845 -3070 3437
rect -1046 2845 -1012 3437
rect 1012 2845 1046 3437
rect 3070 2845 3104 3437
rect -3104 751 -3070 1343
rect -1046 751 -1012 1343
rect 1012 751 1046 1343
rect 3070 751 3104 1343
rect -3104 -1343 -3070 -751
rect -1046 -1343 -1012 -751
rect 1012 -1343 1046 -751
rect 3070 -1343 3104 -751
rect -3104 -3437 -3070 -2845
rect -1046 -3437 -1012 -2845
rect 1012 -3437 1046 -2845
rect 3070 -3437 3104 -2845
<< metal1 >>
rect -3110 3437 -3064 3449
rect -3110 2845 -3104 3437
rect -3070 2845 -3064 3437
rect -3110 2833 -3064 2845
rect -1052 3437 -1006 3449
rect -1052 2845 -1046 3437
rect -1012 2845 -1006 3437
rect -1052 2833 -1006 2845
rect 1006 3437 1052 3449
rect 1006 2845 1012 3437
rect 1046 2845 1052 3437
rect 1006 2833 1052 2845
rect 3064 3437 3110 3449
rect 3064 2845 3070 3437
rect 3104 2845 3110 3437
rect 3064 2833 3110 2845
rect -3110 1343 -3064 1355
rect -3110 751 -3104 1343
rect -3070 751 -3064 1343
rect -3110 739 -3064 751
rect -1052 1343 -1006 1355
rect -1052 751 -1046 1343
rect -1012 751 -1006 1343
rect -1052 739 -1006 751
rect 1006 1343 1052 1355
rect 1006 751 1012 1343
rect 1046 751 1052 1343
rect 1006 739 1052 751
rect 3064 1343 3110 1355
rect 3064 751 3070 1343
rect 3104 751 3110 1343
rect 3064 739 3110 751
rect -3110 -751 -3064 -739
rect -3110 -1343 -3104 -751
rect -3070 -1343 -3064 -751
rect -3110 -1355 -3064 -1343
rect -1052 -751 -1006 -739
rect -1052 -1343 -1046 -751
rect -1012 -1343 -1006 -751
rect -1052 -1355 -1006 -1343
rect 1006 -751 1052 -739
rect 1006 -1343 1012 -751
rect 1046 -1343 1052 -751
rect 1006 -1355 1052 -1343
rect 3064 -751 3110 -739
rect 3064 -1343 3070 -751
rect 3104 -1343 3110 -751
rect 3064 -1355 3110 -1343
rect -3110 -2845 -3064 -2833
rect -3110 -3437 -3104 -2845
rect -3070 -3437 -3064 -2845
rect -3110 -3449 -3064 -3437
rect -1052 -2845 -1006 -2833
rect -1052 -3437 -1046 -2845
rect -1012 -3437 -1006 -2845
rect -1052 -3449 -1006 -3437
rect 1006 -2845 1052 -2833
rect 1006 -3437 1012 -2845
rect 1046 -3437 1052 -2845
rect 1006 -3449 1052 -3437
rect 3064 -2845 3110 -2833
rect 3064 -3437 3070 -2845
rect 3104 -3437 3110 -2845
rect 3064 -3449 3110 -3437
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string parameters w 10 l 10 m 4 nf 3 diffcov 30 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 30 viadrn 30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
