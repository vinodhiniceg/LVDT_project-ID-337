magic
tech sky130A
timestamp 1634305305
<< mvpsubdiff >>
rect 3049 -2167 6505 -1911
rect 3049 -4983 3561 -2167
rect 5929 -4983 6505 -2167
rect 3049 -5239 6505 -4983
rect 12073 -2103 15593 -1783
rect 12073 -4407 12521 -2103
rect 15209 -4407 15593 -2103
rect 12073 -5175 15593 -4407
rect 19817 -2423 23337 -1975
rect 19817 -4983 20265 -2423
rect 23017 -4983 23337 -2423
rect 19817 -5431 23337 -4983
rect 28713 -2231 32233 -2039
rect 28713 -4791 29033 -2231
rect 31785 -4791 32233 -2231
rect 28713 -5495 32233 -4791
rect 36905 -2167 40425 -1847
rect 36905 -4727 37161 -2167
rect 39913 -4727 40425 -2167
rect 36905 -5303 40425 -4727
rect 46313 -2103 49833 -1847
rect 46313 -4663 46633 -2103
rect 49385 -4663 49833 -2103
rect 46313 -5303 49833 -4663
<< mvpsubdiffcont >>
rect 3561 -4983 5929 -2167
rect 12521 -4407 15209 -2103
rect 20265 -4983 23017 -2423
rect 29033 -4791 31785 -2231
rect 37161 -4727 39913 -2167
rect 46633 -4663 49385 -2103
<< poly >>
rect 15051 21976 15615 22035
rect 41800 16228 42206 16354
<< locali >>
rect 19880 16160 20016 16270
rect 31476 15794 31557 16181
rect 44699 15599 45205 15779
rect 44991 14088 45205 15599
rect 4235 -1911 5076 1599
rect 3049 -2167 6505 -1911
rect 3049 -4983 3561 -2167
rect 5929 -4983 6505 -2167
rect 3049 -5239 6505 -4983
rect 12073 -2103 15593 -1783
rect 12073 -4407 12521 -2103
rect 15209 -4407 15593 -2103
rect 12073 -5175 15593 -4407
rect 19817 -2423 23337 -1975
rect 29789 -2039 30031 2810
rect 30924 -2039 31310 1923
rect 37313 -1847 37784 992
rect 48045 -1847 48516 1030
rect 19817 -4983 20265 -2423
rect 23017 -4983 23337 -2423
rect 19817 -5431 23337 -4983
rect 28713 -2231 32233 -2039
rect 28713 -4791 29033 -2231
rect 31785 -4791 32233 -2231
rect 28713 -5495 32233 -4791
rect 36905 -2167 40425 -1847
rect 36905 -4727 37161 -2167
rect 39913 -4727 40425 -2167
rect 36905 -5303 40425 -4727
rect 46313 -2103 49833 -1847
rect 46313 -4663 46633 -2103
rect 49385 -4663 49833 -2103
rect 46313 -5303 49833 -4663
<< viali >>
rect 20016 16102 20162 16286
rect 4009 -4535 5289 -2359
rect 12841 -3959 14889 -2423
rect 20713 -4407 22441 -2743
rect 29417 -4343 31145 -2679
rect 37545 -4151 39273 -2487
rect 47337 -4215 49065 -2551
<< metal1 >>
rect 10692 21473 10820 23216
rect 38462 16456 38631 16469
rect 31809 16430 38644 16456
rect 31783 16299 38644 16430
rect 20013 16286 20165 16292
rect 20013 16102 20016 16286
rect 20162 16260 20165 16286
rect 31783 16260 31939 16299
rect 20162 16169 31939 16260
rect 20162 16166 31926 16169
rect 20162 16102 20165 16166
rect 20013 16096 20165 16102
rect 38462 15464 38631 16299
rect -407 -2359 56361 -1463
rect -407 -4535 4009 -2359
rect 5289 -2423 56361 -2359
rect 5289 -3959 12841 -2423
rect 14889 -2487 56361 -2423
rect 14889 -2679 37545 -2487
rect 14889 -2743 29417 -2679
rect 14889 -3959 20713 -2743
rect 5289 -4407 20713 -3959
rect 22441 -4343 29417 -2743
rect 31145 -4151 37545 -2679
rect 39273 -2551 56361 -2487
rect 39273 -4151 47337 -2551
rect 31145 -4215 47337 -4151
rect 49065 -4215 56361 -2551
rect 31145 -4343 56361 -4215
rect 22441 -4407 56361 -4343
rect 5289 -4535 56361 -4407
rect -407 -6199 56361 -4535
use nmos551535  nmos551535_0 ~/layout test
timestamp 1634301196
transform 1 0 -12764 0 1 1390
box 12764 -1390 42910 21326
use nmos1010514guard  nmos1010514guard_0 ~/layout test
timestamp 1634050450
transform 1 0 30952 0 1 598
box -191 -717 21211 16419
<< labels >>
flabel metal1 745 -4599 745 -4599 0 FreeSans 8000 0 0 0 vssa
flabel poly 41941 16285 41941 16285 0 FreeSans 2400 0 0 0 vin2
flabel poly 15355 22018 15355 22018 0 FreeSans 2400 0 0 0 vin1
flabel metal1 34561 16391 34561 16391 0 FreeSans 800 0 0 0 vcap
flabel metal1 10728 22986 10728 22986 0 FreeSans 800 0 0 0 vout
<< end >>
