magic
tech sky130A
timestamp 1634206023
<< metal3 >>
rect -6477 327 -6409 2605
rect -6577 -147 -6375 327
rect -4331 304 -4263 2605
rect -4417 -147 -4215 304
rect -2185 278 -2117 2606
rect -39 317 29 2601
rect -2270 1 -2068 278
rect -2270 0 -2046 1
rect -2270 -147 -2068 0
rect -133 -147 69 317
rect -6577 -335 78 -147
<< metal4 >>
rect -5539 3058 1190 3060
rect -7633 3047 1190 3058
rect -7634 2837 1190 3047
rect -7634 2316 -7414 2837
rect -5539 2808 1190 2837
rect -5533 2206 -5313 2808
rect -3354 2155 -3134 2808
rect -1208 2181 -988 2808
rect 938 2277 1158 2808
use sky130_fd_pr__cap_mim_m3_1_DCN5A5  sky130_fd_pr__cap_mim_m3_1_DCN5A5_0
timestamp 1634205847
transform 1 0 -3224 0 1 1300
box -5360 -1300 5360 1300
<< labels >>
rlabel metal4 -3432 2937 -3432 2937 5 top
rlabel metal3 -2701 -276 -2701 -276 5 bot
<< end >>
