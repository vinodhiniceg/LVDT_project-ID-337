magic
tech sky130A
magscale 1 2
timestamp 1634118957
<< error_p >>
rect -2727 1056 2727 1060
rect -2727 -1056 -2697 1056
rect -2661 990 2661 994
rect -2661 394 -2631 990
rect 2631 394 2661 990
rect -2661 -300 -2631 300
rect 2631 -300 2661 300
rect -2661 -990 -2631 -394
rect 2631 -990 2661 -394
rect -2661 -994 2661 -990
rect 2697 -1056 2727 1056
rect -2727 -1060 2727 -1056
<< nwell >>
rect -2697 -1056 2697 1056
<< mvpmos >>
rect -2603 394 -2003 994
rect -1945 394 -1345 994
rect -1287 394 -687 994
rect -629 394 -29 994
rect 29 394 629 994
rect 687 394 1287 994
rect 1345 394 1945 994
rect 2003 394 2603 994
rect -2603 -300 -2003 300
rect -1945 -300 -1345 300
rect -1287 -300 -687 300
rect -629 -300 -29 300
rect 29 -300 629 300
rect 687 -300 1287 300
rect 1345 -300 1945 300
rect 2003 -300 2603 300
rect -2603 -994 -2003 -394
rect -1945 -994 -1345 -394
rect -1287 -994 -687 -394
rect -629 -994 -29 -394
rect 29 -994 629 -394
rect 687 -994 1287 -394
rect 1345 -994 1945 -394
rect 2003 -994 2603 -394
<< mvpdiff >>
rect -2661 780 -2603 994
rect -2661 608 -2649 780
rect -2615 608 -2603 780
rect -2661 394 -2603 608
rect -2003 780 -1945 994
rect -2003 608 -1991 780
rect -1957 608 -1945 780
rect -2003 394 -1945 608
rect -1345 780 -1287 994
rect -1345 608 -1333 780
rect -1299 608 -1287 780
rect -1345 394 -1287 608
rect -687 780 -629 994
rect -687 608 -675 780
rect -641 608 -629 780
rect -687 394 -629 608
rect -29 780 29 994
rect -29 608 -17 780
rect 17 608 29 780
rect -29 394 29 608
rect 629 780 687 994
rect 629 608 641 780
rect 675 608 687 780
rect 629 394 687 608
rect 1287 780 1345 994
rect 1287 608 1299 780
rect 1333 608 1345 780
rect 1287 394 1345 608
rect 1945 780 2003 994
rect 1945 608 1957 780
rect 1991 608 2003 780
rect 1945 394 2003 608
rect 2603 780 2661 994
rect 2603 608 2615 780
rect 2649 608 2661 780
rect 2603 394 2661 608
rect -2661 86 -2603 300
rect -2661 -86 -2649 86
rect -2615 -86 -2603 86
rect -2661 -300 -2603 -86
rect -2003 86 -1945 300
rect -2003 -86 -1991 86
rect -1957 -86 -1945 86
rect -2003 -300 -1945 -86
rect -1345 86 -1287 300
rect -1345 -86 -1333 86
rect -1299 -86 -1287 86
rect -1345 -300 -1287 -86
rect -687 86 -629 300
rect -687 -86 -675 86
rect -641 -86 -629 86
rect -687 -300 -629 -86
rect -29 86 29 300
rect -29 -86 -17 86
rect 17 -86 29 86
rect -29 -300 29 -86
rect 629 86 687 300
rect 629 -86 641 86
rect 675 -86 687 86
rect 629 -300 687 -86
rect 1287 86 1345 300
rect 1287 -86 1299 86
rect 1333 -86 1345 86
rect 1287 -300 1345 -86
rect 1945 86 2003 300
rect 1945 -86 1957 86
rect 1991 -86 2003 86
rect 1945 -300 2003 -86
rect 2603 86 2661 300
rect 2603 -86 2615 86
rect 2649 -86 2661 86
rect 2603 -300 2661 -86
rect -2661 -608 -2603 -394
rect -2661 -780 -2649 -608
rect -2615 -780 -2603 -608
rect -2661 -994 -2603 -780
rect -2003 -608 -1945 -394
rect -2003 -780 -1991 -608
rect -1957 -780 -1945 -608
rect -2003 -994 -1945 -780
rect -1345 -608 -1287 -394
rect -1345 -780 -1333 -608
rect -1299 -780 -1287 -608
rect -1345 -994 -1287 -780
rect -687 -608 -629 -394
rect -687 -780 -675 -608
rect -641 -780 -629 -608
rect -687 -994 -629 -780
rect -29 -608 29 -394
rect -29 -780 -17 -608
rect 17 -780 29 -608
rect -29 -994 29 -780
rect 629 -608 687 -394
rect 629 -780 641 -608
rect 675 -780 687 -608
rect 629 -994 687 -780
rect 1287 -608 1345 -394
rect 1287 -780 1299 -608
rect 1333 -780 1345 -608
rect 1287 -994 1345 -780
rect 1945 -608 2003 -394
rect 1945 -780 1957 -608
rect 1991 -780 2003 -608
rect 1945 -994 2003 -780
rect 2603 -608 2661 -394
rect 2603 -780 2615 -608
rect 2649 -780 2661 -608
rect 2603 -994 2661 -780
<< mvpdiffc >>
rect -2649 608 -2615 780
rect -1991 608 -1957 780
rect -1333 608 -1299 780
rect -675 608 -641 780
rect -17 608 17 780
rect 641 608 675 780
rect 1299 608 1333 780
rect 1957 608 1991 780
rect 2615 608 2649 780
rect -2649 -86 -2615 86
rect -1991 -86 -1957 86
rect -1333 -86 -1299 86
rect -675 -86 -641 86
rect -17 -86 17 86
rect 641 -86 675 86
rect 1299 -86 1333 86
rect 1957 -86 1991 86
rect 2615 -86 2649 86
rect -2649 -780 -2615 -608
rect -1991 -780 -1957 -608
rect -1333 -780 -1299 -608
rect -675 -780 -641 -608
rect -17 -780 17 -608
rect 641 -780 675 -608
rect 1299 -780 1333 -608
rect 1957 -780 1991 -608
rect 2615 -780 2649 -608
<< poly >>
rect -2603 994 -2003 1020
rect -1945 994 -1345 1020
rect -1287 994 -687 1020
rect -629 994 -29 1020
rect 29 994 629 1020
rect 687 994 1287 1020
rect 1345 994 1945 1020
rect 2003 994 2603 1020
rect -2603 368 -2003 394
rect -1945 368 -1345 394
rect -1287 368 -687 394
rect -629 368 -29 394
rect 29 368 629 394
rect 687 368 1287 394
rect 1345 368 1945 394
rect 2003 368 2603 394
rect -2603 300 -2003 326
rect -1945 300 -1345 326
rect -1287 300 -687 326
rect -629 300 -29 326
rect 29 300 629 326
rect 687 300 1287 326
rect 1345 300 1945 326
rect 2003 300 2603 326
rect -2603 -326 -2003 -300
rect -1945 -326 -1345 -300
rect -1287 -326 -687 -300
rect -629 -326 -29 -300
rect 29 -326 629 -300
rect 687 -326 1287 -300
rect 1345 -326 1945 -300
rect 2003 -326 2603 -300
rect -2603 -394 -2003 -368
rect -1945 -394 -1345 -368
rect -1287 -394 -687 -368
rect -629 -394 -29 -368
rect 29 -394 629 -368
rect 687 -394 1287 -368
rect 1345 -394 1945 -368
rect 2003 -394 2603 -368
rect -2603 -1020 -2003 -994
rect -1945 -1020 -1345 -994
rect -1287 -1020 -687 -994
rect -629 -1020 -29 -994
rect 29 -1020 629 -994
rect 687 -1020 1287 -994
rect 1345 -1020 1945 -994
rect 2003 -1020 2603 -994
<< locali >>
rect -2649 780 -2615 796
rect -2649 592 -2615 608
rect -1991 780 -1957 796
rect -1991 592 -1957 608
rect -1333 780 -1299 796
rect -1333 592 -1299 608
rect -675 780 -641 796
rect -675 592 -641 608
rect -17 780 17 796
rect -17 592 17 608
rect 641 780 675 796
rect 641 592 675 608
rect 1299 780 1333 796
rect 1299 592 1333 608
rect 1957 780 1991 796
rect 1957 592 1991 608
rect 2615 780 2649 796
rect 2615 592 2649 608
rect -2649 86 -2615 102
rect -2649 -102 -2615 -86
rect -1991 86 -1957 102
rect -1991 -102 -1957 -86
rect -1333 86 -1299 102
rect -1333 -102 -1299 -86
rect -675 86 -641 102
rect -675 -102 -641 -86
rect -17 86 17 102
rect -17 -102 17 -86
rect 641 86 675 102
rect 641 -102 675 -86
rect 1299 86 1333 102
rect 1299 -102 1333 -86
rect 1957 86 1991 102
rect 1957 -102 1991 -86
rect 2615 86 2649 102
rect 2615 -102 2649 -86
rect -2649 -608 -2615 -592
rect -2649 -796 -2615 -780
rect -1991 -608 -1957 -592
rect -1991 -796 -1957 -780
rect -1333 -608 -1299 -592
rect -1333 -796 -1299 -780
rect -675 -608 -641 -592
rect -675 -796 -641 -780
rect -17 -608 17 -592
rect -17 -796 17 -780
rect 641 -608 675 -592
rect 641 -796 675 -780
rect 1299 -608 1333 -592
rect 1299 -796 1333 -780
rect 1957 -608 1991 -592
rect 1957 -796 1991 -780
rect 2615 -608 2649 -592
rect 2615 -796 2649 -780
<< viali >>
rect -2649 608 -2615 780
rect -1991 608 -1957 780
rect -1333 608 -1299 780
rect -675 608 -641 780
rect -17 608 17 780
rect 641 608 675 780
rect 1299 608 1333 780
rect 1957 608 1991 780
rect 2615 608 2649 780
rect -2649 -86 -2615 86
rect -1991 -86 -1957 86
rect -1333 -86 -1299 86
rect -675 -86 -641 86
rect -17 -86 17 86
rect 641 -86 675 86
rect 1299 -86 1333 86
rect 1957 -86 1991 86
rect 2615 -86 2649 86
rect -2649 -780 -2615 -608
rect -1991 -780 -1957 -608
rect -1333 -780 -1299 -608
rect -675 -780 -641 -608
rect -17 -780 17 -608
rect 641 -780 675 -608
rect 1299 -780 1333 -608
rect 1957 -780 1991 -608
rect 2615 -780 2649 -608
<< metal1 >>
rect -2655 780 -2609 792
rect -2655 608 -2649 780
rect -2615 608 -2609 780
rect -2655 596 -2609 608
rect -1997 780 -1951 792
rect -1997 608 -1991 780
rect -1957 608 -1951 780
rect -1997 596 -1951 608
rect -1339 780 -1293 792
rect -1339 608 -1333 780
rect -1299 608 -1293 780
rect -1339 596 -1293 608
rect -681 780 -635 792
rect -681 608 -675 780
rect -641 608 -635 780
rect -681 596 -635 608
rect -23 780 23 792
rect -23 608 -17 780
rect 17 608 23 780
rect -23 596 23 608
rect 635 780 681 792
rect 635 608 641 780
rect 675 608 681 780
rect 635 596 681 608
rect 1293 780 1339 792
rect 1293 608 1299 780
rect 1333 608 1339 780
rect 1293 596 1339 608
rect 1951 780 1997 792
rect 1951 608 1957 780
rect 1991 608 1997 780
rect 1951 596 1997 608
rect 2609 780 2655 792
rect 2609 608 2615 780
rect 2649 608 2655 780
rect 2609 596 2655 608
rect -2655 86 -2609 98
rect -2655 -86 -2649 86
rect -2615 -86 -2609 86
rect -2655 -98 -2609 -86
rect -1997 86 -1951 98
rect -1997 -86 -1991 86
rect -1957 -86 -1951 86
rect -1997 -98 -1951 -86
rect -1339 86 -1293 98
rect -1339 -86 -1333 86
rect -1299 -86 -1293 86
rect -1339 -98 -1293 -86
rect -681 86 -635 98
rect -681 -86 -675 86
rect -641 -86 -635 86
rect -681 -98 -635 -86
rect -23 86 23 98
rect -23 -86 -17 86
rect 17 -86 23 86
rect -23 -98 23 -86
rect 635 86 681 98
rect 635 -86 641 86
rect 675 -86 681 86
rect 635 -98 681 -86
rect 1293 86 1339 98
rect 1293 -86 1299 86
rect 1333 -86 1339 86
rect 1293 -98 1339 -86
rect 1951 86 1997 98
rect 1951 -86 1957 86
rect 1991 -86 1997 86
rect 1951 -98 1997 -86
rect 2609 86 2655 98
rect 2609 -86 2615 86
rect 2649 -86 2655 86
rect 2609 -98 2655 -86
rect -2655 -608 -2609 -596
rect -2655 -780 -2649 -608
rect -2615 -780 -2609 -608
rect -2655 -792 -2609 -780
rect -1997 -608 -1951 -596
rect -1997 -780 -1991 -608
rect -1957 -780 -1951 -608
rect -1997 -792 -1951 -780
rect -1339 -608 -1293 -596
rect -1339 -780 -1333 -608
rect -1299 -780 -1293 -608
rect -1339 -792 -1293 -780
rect -681 -608 -635 -596
rect -681 -780 -675 -608
rect -641 -780 -635 -608
rect -681 -792 -635 -780
rect -23 -608 23 -596
rect -23 -780 -17 -608
rect 17 -780 23 -608
rect -23 -792 23 -780
rect 635 -608 681 -596
rect 635 -780 641 -608
rect 675 -780 681 -608
rect 635 -792 681 -780
rect 1293 -608 1339 -596
rect 1293 -780 1299 -608
rect 1333 -780 1339 -608
rect 1293 -792 1339 -780
rect 1951 -608 1997 -596
rect 1951 -780 1957 -608
rect 1991 -780 1997 -608
rect 1951 -792 1997 -780
rect 2609 -608 2655 -596
rect 2609 -780 2615 -608
rect 2649 -780 2655 -608
rect 2609 -792 2655 -780
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string parameters w 3 l 3 m 3 nf 8 diffcov 30 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 30 viadrn 30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
