magic
tech sky130A
magscale 1 2
timestamp 1634127866
<< pwell >>
rect -126 6886 2354 7116
rect -126 6758 1426 6886
rect 1996 6858 2354 6886
rect -444 6716 1426 6758
rect 2048 6716 2354 6858
rect -444 4182 2354 6716
rect -124 2864 2354 4182
rect -444 532 2354 2864
rect -110 208 2354 532
rect -110 66 1260 208
rect 1882 66 2354 208
rect -110 -236 2354 66
<< mvpsubdiff >>
rect -444 6718 -144 6758
rect -444 4356 -344 6718
rect -250 4356 -144 6718
rect -444 4182 -144 4356
rect -444 2782 -144 2864
rect -444 582 -396 2782
rect -196 582 -144 2782
rect -444 532 -144 582
<< mvpsubdiffcont >>
rect -344 4356 -250 6718
rect -396 582 -196 2782
<< poly >>
rect 242 6892 1836 6944
rect 130 6192 592 6262
rect 814 6190 1276 6260
rect 1486 6192 1948 6262
rect 160 5498 622 5568
rect 800 5492 1262 5562
rect 1462 5496 1924 5566
rect 134 4796 596 4866
rect 800 4802 1262 4872
rect 1454 4800 1916 4870
rect 172 4104 634 4174
rect 818 4106 1280 4176
rect 1466 4106 1928 4176
rect 160 3416 622 3486
rect 808 3412 1270 3482
rect 1446 3416 1908 3486
rect 130 2716 592 2786
rect 814 2714 1276 2784
rect 1456 2720 1918 2790
rect 140 2022 602 2092
rect 796 2022 1258 2092
rect 1460 2026 1922 2096
rect 138 1332 600 1402
rect 792 1334 1254 1404
rect 1436 1328 1898 1398
rect 154 636 616 706
rect 808 636 1270 706
rect 1432 634 1894 704
<< locali >>
rect 1316 6820 1384 6828
rect -400 6718 -194 6758
rect -10 6748 1426 6820
rect -400 4356 -344 6718
rect -250 4356 -194 6718
rect -6 6596 62 6748
rect 1316 6640 1384 6748
rect -400 4190 -194 4356
rect -428 2782 -172 2854
rect -428 582 -396 2782
rect -196 582 -172 2782
rect -428 532 -172 582
rect -4 326 48 6596
rect 664 390 716 6588
rect 1314 6568 1386 6640
rect 648 252 718 390
rect 1314 350 1366 6568
rect 1974 6538 2034 6664
rect 1982 382 2034 6538
rect 658 122 718 252
rect 1308 208 1368 350
rect 1944 128 2058 382
rect 1204 122 2058 128
rect 650 70 2058 122
rect 1204 52 2058 70
rect 1944 48 2058 52
<< viali >>
rect -334 4394 -274 6694
rect -364 694 -244 2694
<< metal1 >>
rect -400 6694 -194 6758
rect -400 4394 -334 6694
rect -274 4394 -194 6694
rect -400 4190 -194 4394
rect -428 2694 -172 2854
rect -428 694 -364 2694
rect -244 694 -172 2694
rect -428 532 -172 694
use sky130_fd_pr__nfet_g5v0d10v5_7Z98EG  sky130_fd_pr__nfet_g5v0d10v5_7Z98EG_0 ~/layout test
timestamp 1634127529
transform 1 0 1016 0 1 3449
box -1016 -3449 1016 3449
<< end >>
