magic
tech sky130A
timestamp 1634297993
<< pwell >>
rect -1422 -1442 1422 1442
<< mvnmos >>
rect -1308 844 -808 1344
rect -779 844 -279 1344
rect -250 844 250 1344
rect 279 844 779 1344
rect 808 844 1308 1344
rect -1308 297 -808 797
rect -779 297 -279 797
rect -250 297 250 797
rect 279 297 779 797
rect 808 297 1308 797
rect -1308 -250 -808 250
rect -779 -250 -279 250
rect -250 -250 250 250
rect 279 -250 779 250
rect 808 -250 1308 250
rect -1308 -797 -808 -297
rect -779 -797 -279 -297
rect -250 -797 250 -297
rect 279 -797 779 -297
rect 808 -797 1308 -297
rect -1308 -1344 -808 -844
rect -779 -1344 -279 -844
rect -250 -1344 250 -844
rect 279 -1344 779 -844
rect 808 -1344 1308 -844
<< mvndiff >>
rect -1337 1167 -1308 1344
rect -1337 1021 -1331 1167
rect -1314 1021 -1308 1167
rect -1337 844 -1308 1021
rect -808 1167 -779 1344
rect -808 1021 -802 1167
rect -785 1021 -779 1167
rect -808 844 -779 1021
rect -279 1167 -250 1344
rect -279 1021 -273 1167
rect -256 1021 -250 1167
rect -279 844 -250 1021
rect 250 1167 279 1344
rect 250 1021 256 1167
rect 273 1021 279 1167
rect 250 844 279 1021
rect 779 1167 808 1344
rect 779 1021 785 1167
rect 802 1021 808 1167
rect 779 844 808 1021
rect 1308 1167 1337 1344
rect 1308 1021 1314 1167
rect 1331 1021 1337 1167
rect 1308 844 1337 1021
rect -1337 620 -1308 797
rect -1337 474 -1331 620
rect -1314 474 -1308 620
rect -1337 297 -1308 474
rect -808 620 -779 797
rect -808 474 -802 620
rect -785 474 -779 620
rect -808 297 -779 474
rect -279 620 -250 797
rect -279 474 -273 620
rect -256 474 -250 620
rect -279 297 -250 474
rect 250 620 279 797
rect 250 474 256 620
rect 273 474 279 620
rect 250 297 279 474
rect 779 620 808 797
rect 779 474 785 620
rect 802 474 808 620
rect 779 297 808 474
rect 1308 620 1337 797
rect 1308 474 1314 620
rect 1331 474 1337 620
rect 1308 297 1337 474
rect -1337 73 -1308 250
rect -1337 -73 -1331 73
rect -1314 -73 -1308 73
rect -1337 -250 -1308 -73
rect -808 73 -779 250
rect -808 -73 -802 73
rect -785 -73 -779 73
rect -808 -250 -779 -73
rect -279 73 -250 250
rect -279 -73 -273 73
rect -256 -73 -250 73
rect -279 -250 -250 -73
rect 250 73 279 250
rect 250 -73 256 73
rect 273 -73 279 73
rect 250 -250 279 -73
rect 779 73 808 250
rect 779 -73 785 73
rect 802 -73 808 73
rect 779 -250 808 -73
rect 1308 73 1337 250
rect 1308 -73 1314 73
rect 1331 -73 1337 73
rect 1308 -250 1337 -73
rect -1337 -474 -1308 -297
rect -1337 -620 -1331 -474
rect -1314 -620 -1308 -474
rect -1337 -797 -1308 -620
rect -808 -474 -779 -297
rect -808 -620 -802 -474
rect -785 -620 -779 -474
rect -808 -797 -779 -620
rect -279 -474 -250 -297
rect -279 -620 -273 -474
rect -256 -620 -250 -474
rect -279 -797 -250 -620
rect 250 -474 279 -297
rect 250 -620 256 -474
rect 273 -620 279 -474
rect 250 -797 279 -620
rect 779 -474 808 -297
rect 779 -620 785 -474
rect 802 -620 808 -474
rect 779 -797 808 -620
rect 1308 -474 1337 -297
rect 1308 -620 1314 -474
rect 1331 -620 1337 -474
rect 1308 -797 1337 -620
rect -1337 -1021 -1308 -844
rect -1337 -1167 -1331 -1021
rect -1314 -1167 -1308 -1021
rect -1337 -1344 -1308 -1167
rect -808 -1021 -779 -844
rect -808 -1167 -802 -1021
rect -785 -1167 -779 -1021
rect -808 -1344 -779 -1167
rect -279 -1021 -250 -844
rect -279 -1167 -273 -1021
rect -256 -1167 -250 -1021
rect -279 -1344 -250 -1167
rect 250 -1021 279 -844
rect 250 -1167 256 -1021
rect 273 -1167 279 -1021
rect 250 -1344 279 -1167
rect 779 -1021 808 -844
rect 779 -1167 785 -1021
rect 802 -1167 808 -1021
rect 779 -1344 808 -1167
rect 1308 -1021 1337 -844
rect 1308 -1167 1314 -1021
rect 1331 -1167 1337 -1021
rect 1308 -1344 1337 -1167
<< mvndiffc >>
rect -1331 1021 -1314 1167
rect -802 1021 -785 1167
rect -273 1021 -256 1167
rect 256 1021 273 1167
rect 785 1021 802 1167
rect 1314 1021 1331 1167
rect -1331 474 -1314 620
rect -802 474 -785 620
rect -273 474 -256 620
rect 256 474 273 620
rect 785 474 802 620
rect 1314 474 1331 620
rect -1331 -73 -1314 73
rect -802 -73 -785 73
rect -273 -73 -256 73
rect 256 -73 273 73
rect 785 -73 802 73
rect 1314 -73 1331 73
rect -1331 -620 -1314 -474
rect -802 -620 -785 -474
rect -273 -620 -256 -474
rect 256 -620 273 -474
rect 785 -620 802 -474
rect 1314 -620 1331 -474
rect -1331 -1167 -1314 -1021
rect -802 -1167 -785 -1021
rect -273 -1167 -256 -1021
rect 256 -1167 273 -1021
rect 785 -1167 802 -1021
rect 1314 -1167 1331 -1021
<< mvpsubdiff >>
rect -1404 1395 1404 1424
rect -1404 685 -1375 1395
rect -1404 -685 -1398 685
rect -1381 -685 -1375 685
rect 1375 685 1404 1395
rect -1404 -1395 -1375 -685
rect 1375 -685 1381 685
rect 1398 -685 1404 685
rect 1375 -1395 1404 -685
rect -1404 -1424 1404 -1395
<< mvpsubdiffcont >>
rect -1398 -685 -1381 685
rect 1381 -685 1398 685
<< poly >>
rect -1308 1344 -808 1357
rect -779 1344 -279 1357
rect -250 1344 250 1357
rect 279 1344 779 1357
rect 808 1344 1308 1357
rect -1308 831 -808 844
rect -779 831 -279 844
rect -250 831 250 844
rect 279 831 779 844
rect 808 831 1308 844
rect -1308 797 -808 810
rect -779 797 -279 810
rect -250 797 250 810
rect 279 797 779 810
rect 808 797 1308 810
rect -1308 284 -808 297
rect -779 284 -279 297
rect -250 284 250 297
rect 279 284 779 297
rect 808 284 1308 297
rect -1308 250 -808 263
rect -779 250 -279 263
rect -250 250 250 263
rect 279 250 779 263
rect 808 250 1308 263
rect -1308 -263 -808 -250
rect -779 -263 -279 -250
rect -250 -263 250 -250
rect 279 -263 779 -250
rect 808 -263 1308 -250
rect -1308 -297 -808 -284
rect -779 -297 -279 -284
rect -250 -297 250 -284
rect 279 -297 779 -284
rect 808 -297 1308 -284
rect -1308 -810 -808 -797
rect -779 -810 -279 -797
rect -250 -810 250 -797
rect 279 -810 779 -797
rect 808 -810 1308 -797
rect -1308 -844 -808 -831
rect -779 -844 -279 -831
rect -250 -844 250 -831
rect 279 -844 779 -831
rect 808 -844 1308 -831
rect -1308 -1357 -808 -1344
rect -779 -1357 -279 -1344
rect -250 -1357 250 -1344
rect 279 -1357 779 -1344
rect 808 -1357 1308 -1344
<< locali >>
rect -1398 1401 1398 1418
rect -1398 685 -1381 1401
rect -1331 1167 -1314 1175
rect -1331 1013 -1314 1021
rect -802 1167 -785 1175
rect -802 1013 -785 1021
rect -273 1167 -256 1175
rect -273 1013 -256 1021
rect 256 1167 273 1175
rect 256 1013 273 1021
rect 785 1167 802 1175
rect 785 1013 802 1021
rect 1314 1167 1331 1175
rect 1314 1013 1331 1021
rect 1381 685 1398 1401
rect -1331 620 -1314 628
rect -1331 466 -1314 474
rect -802 620 -785 628
rect -802 466 -785 474
rect -273 620 -256 628
rect -273 466 -256 474
rect 256 620 273 628
rect 256 466 273 474
rect 785 620 802 628
rect 785 466 802 474
rect 1314 620 1331 628
rect 1314 466 1331 474
rect -1331 73 -1314 81
rect -1331 -81 -1314 -73
rect -802 73 -785 81
rect -802 -81 -785 -73
rect -273 73 -256 81
rect -273 -81 -256 -73
rect 256 73 273 81
rect 256 -81 273 -73
rect 785 73 802 81
rect 785 -81 802 -73
rect 1314 73 1331 81
rect 1314 -81 1331 -73
rect -1331 -474 -1314 -466
rect -1331 -628 -1314 -620
rect -802 -474 -785 -466
rect -802 -628 -785 -620
rect -273 -474 -256 -466
rect -273 -628 -256 -620
rect 256 -474 273 -466
rect 256 -628 273 -620
rect 785 -474 802 -466
rect 785 -628 802 -620
rect 1314 -474 1331 -466
rect 1314 -628 1331 -620
rect -1398 -1401 -1381 -685
rect -1331 -1021 -1314 -1013
rect -1331 -1175 -1314 -1167
rect -802 -1021 -785 -1013
rect -802 -1175 -785 -1167
rect -273 -1021 -256 -1013
rect -273 -1175 -256 -1167
rect 256 -1021 273 -1013
rect 256 -1175 273 -1167
rect 785 -1021 802 -1013
rect 785 -1175 802 -1167
rect 1314 -1021 1331 -1013
rect 1314 -1175 1331 -1167
rect 1381 -1401 1398 -685
rect -1398 -1418 1398 -1401
<< viali >>
rect -1331 1021 -1314 1167
rect -802 1021 -785 1167
rect -273 1021 -256 1167
rect 256 1021 273 1167
rect 785 1021 802 1167
rect 1314 1021 1331 1167
rect -1331 474 -1314 620
rect -802 474 -785 620
rect -273 474 -256 620
rect 256 474 273 620
rect 785 474 802 620
rect 1314 474 1331 620
rect -1331 -73 -1314 73
rect -802 -73 -785 73
rect -273 -73 -256 73
rect 256 -73 273 73
rect 785 -73 802 73
rect 1314 -73 1331 73
rect -1331 -620 -1314 -474
rect -802 -620 -785 -474
rect -273 -620 -256 -474
rect 256 -620 273 -474
rect 785 -620 802 -474
rect 1314 -620 1331 -474
rect -1331 -1167 -1314 -1021
rect -802 -1167 -785 -1021
rect -273 -1167 -256 -1021
rect 256 -1167 273 -1021
rect 785 -1167 802 -1021
rect 1314 -1167 1331 -1021
<< metal1 >>
rect -1334 1167 -1311 1173
rect -1334 1021 -1331 1167
rect -1314 1021 -1311 1167
rect -1334 1015 -1311 1021
rect -805 1167 -782 1173
rect -805 1021 -802 1167
rect -785 1021 -782 1167
rect -805 1015 -782 1021
rect -276 1167 -253 1173
rect -276 1021 -273 1167
rect -256 1021 -253 1167
rect -276 1015 -253 1021
rect 253 1167 276 1173
rect 253 1021 256 1167
rect 273 1021 276 1167
rect 253 1015 276 1021
rect 782 1167 805 1173
rect 782 1021 785 1167
rect 802 1021 805 1167
rect 782 1015 805 1021
rect 1311 1167 1334 1173
rect 1311 1021 1314 1167
rect 1331 1021 1334 1167
rect 1311 1015 1334 1021
rect -1334 620 -1311 626
rect -1334 474 -1331 620
rect -1314 474 -1311 620
rect -1334 468 -1311 474
rect -805 620 -782 626
rect -805 474 -802 620
rect -785 474 -782 620
rect -805 468 -782 474
rect -276 620 -253 626
rect -276 474 -273 620
rect -256 474 -253 620
rect -276 468 -253 474
rect 253 620 276 626
rect 253 474 256 620
rect 273 474 276 620
rect 253 468 276 474
rect 782 620 805 626
rect 782 474 785 620
rect 802 474 805 620
rect 782 468 805 474
rect 1311 620 1334 626
rect 1311 474 1314 620
rect 1331 474 1334 620
rect 1311 468 1334 474
rect -1334 73 -1311 79
rect -1334 -73 -1331 73
rect -1314 -73 -1311 73
rect -1334 -79 -1311 -73
rect -805 73 -782 79
rect -805 -73 -802 73
rect -785 -73 -782 73
rect -805 -79 -782 -73
rect -276 73 -253 79
rect -276 -73 -273 73
rect -256 -73 -253 73
rect -276 -79 -253 -73
rect 253 73 276 79
rect 253 -73 256 73
rect 273 -73 276 73
rect 253 -79 276 -73
rect 782 73 805 79
rect 782 -73 785 73
rect 802 -73 805 73
rect 782 -79 805 -73
rect 1311 73 1334 79
rect 1311 -73 1314 73
rect 1331 -73 1334 73
rect 1311 -79 1334 -73
rect -1334 -474 -1311 -468
rect -1334 -620 -1331 -474
rect -1314 -620 -1311 -474
rect -1334 -626 -1311 -620
rect -805 -474 -782 -468
rect -805 -620 -802 -474
rect -785 -620 -782 -474
rect -805 -626 -782 -620
rect -276 -474 -253 -468
rect -276 -620 -273 -474
rect -256 -620 -253 -474
rect -276 -626 -253 -620
rect 253 -474 276 -468
rect 253 -620 256 -474
rect 273 -620 276 -474
rect 253 -626 276 -620
rect 782 -474 805 -468
rect 782 -620 785 -474
rect 802 -620 805 -474
rect 782 -626 805 -620
rect 1311 -474 1334 -468
rect 1311 -620 1314 -474
rect 1331 -620 1334 -474
rect 1311 -626 1334 -620
rect -1334 -1021 -1311 -1015
rect -1334 -1167 -1331 -1021
rect -1314 -1167 -1311 -1021
rect -1334 -1173 -1311 -1167
rect -805 -1021 -782 -1015
rect -805 -1167 -802 -1021
rect -785 -1167 -782 -1021
rect -805 -1173 -782 -1167
rect -276 -1021 -253 -1015
rect -276 -1167 -273 -1021
rect -256 -1167 -253 -1021
rect -276 -1173 -253 -1167
rect 253 -1021 276 -1015
rect 253 -1167 256 -1021
rect 273 -1167 276 -1021
rect 253 -1173 276 -1167
rect 782 -1021 805 -1015
rect 782 -1167 785 -1021
rect 802 -1167 805 -1021
rect 782 -1173 805 -1167
rect 1311 -1021 1334 -1015
rect 1311 -1167 1314 -1021
rect 1331 -1167 1334 -1021
rect 1311 -1173 1334 -1167
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string FIXED_BBOX -1389 -1409 1389 1409
string parameters w 5 l 5 m 5 nf 5 diffcov 30 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 50 rlcov 50 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 30 viadrn 30 viagate 30 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
