magic
tech sky130A
magscale 1 2
timestamp 1634112475
<< mvpsubdiff >>
rect 1502 6138 1644 6182
rect 1502 5320 1522 6138
rect 1620 5320 1644 6138
rect 1502 5292 1644 5320
rect 1584 1704 1760 1768
rect 1584 974 1624 1704
rect 1726 974 1760 1704
rect 1584 880 1760 974
<< mvpsubdiffcont >>
rect 1522 5320 1620 6138
rect 1624 974 1726 1704
<< poly >>
rect 406 6890 962 6962
rect 214 6190 478 6258
rect 906 6194 1170 6262
rect 236 5492 500 5560
rect 962 5492 1226 5560
rect 220 4804 484 4872
rect 970 4804 1234 4872
rect 234 4112 498 4180
rect 1020 4112 1284 4180
rect 262 3410 526 3478
rect 984 3410 1248 3478
rect 264 2720 528 2788
rect 966 2714 1230 2782
rect 278 2026 542 2094
rect 992 2020 1256 2088
rect 290 1332 554 1400
rect 938 1332 1202 1400
rect 260 638 524 706
rect 960 646 1224 714
<< locali >>
rect 4 6812 60 6814
rect 0 6808 1372 6812
rect 0 6756 1374 6808
rect 4 6646 60 6756
rect 4 6628 68 6646
rect 6 332 68 6628
rect 662 366 724 6648
rect 1312 6626 1374 6756
rect 1312 6600 1378 6626
rect 660 88 728 366
rect 1316 312 1378 6600
rect 1502 6138 1644 6182
rect 1502 5320 1522 6138
rect 1620 5320 1644 6138
rect 1502 5292 1644 5320
rect 1584 1704 1760 1768
rect 1584 974 1624 1704
rect 1726 974 1760 1704
rect 1584 880 1760 974
<< viali >>
rect 1546 5430 1590 6074
rect 1648 1014 1704 1658
<< metal1 >>
rect 1502 6074 1644 6182
rect 1502 5430 1546 6074
rect 1590 5430 1644 6074
rect 1502 5292 1644 5430
rect 1584 1658 1760 1768
rect 1584 1014 1648 1658
rect 1704 1014 1760 1658
rect 1584 880 1760 1014
use sky130_fd_pr__nfet_g5v0d10v5_MZR6RC  sky130_fd_pr__nfet_g5v0d10v5_MZR6RC_0
timestamp 1634112475
transform 1 0 687 0 1 3449
box -687 -3449 687 3449
<< end >>
