magic
tech sky130A
magscale 1 2
timestamp 1634045799
<< mvnmos >>
rect -2029 3188 -29 5188
rect 29 3188 2029 5188
rect -2029 1094 -29 3094
rect 29 1094 2029 3094
rect -2029 -1000 -29 1000
rect 29 -1000 2029 1000
rect -2029 -3094 -29 -1094
rect 29 -3094 2029 -1094
rect -2029 -5188 -29 -3188
rect 29 -5188 2029 -3188
<< mvndiff >>
rect -2087 4484 -2029 5188
rect -2087 3892 -2075 4484
rect -2041 3892 -2029 4484
rect -2087 3188 -2029 3892
rect -29 4484 29 5188
rect -29 3892 -17 4484
rect 17 3892 29 4484
rect -29 3188 29 3892
rect 2029 4484 2087 5188
rect 2029 3892 2041 4484
rect 2075 3892 2087 4484
rect 2029 3188 2087 3892
rect -2087 2390 -2029 3094
rect -2087 1798 -2075 2390
rect -2041 1798 -2029 2390
rect -2087 1094 -2029 1798
rect -29 2390 29 3094
rect -29 1798 -17 2390
rect 17 1798 29 2390
rect -29 1094 29 1798
rect 2029 2390 2087 3094
rect 2029 1798 2041 2390
rect 2075 1798 2087 2390
rect 2029 1094 2087 1798
rect -2087 296 -2029 1000
rect -2087 -296 -2075 296
rect -2041 -296 -2029 296
rect -2087 -1000 -2029 -296
rect -29 296 29 1000
rect -29 -296 -17 296
rect 17 -296 29 296
rect -29 -1000 29 -296
rect 2029 296 2087 1000
rect 2029 -296 2041 296
rect 2075 -296 2087 296
rect 2029 -1000 2087 -296
rect -2087 -1798 -2029 -1094
rect -2087 -2390 -2075 -1798
rect -2041 -2390 -2029 -1798
rect -2087 -3094 -2029 -2390
rect -29 -1798 29 -1094
rect -29 -2390 -17 -1798
rect 17 -2390 29 -1798
rect -29 -3094 29 -2390
rect 2029 -1798 2087 -1094
rect 2029 -2390 2041 -1798
rect 2075 -2390 2087 -1798
rect 2029 -3094 2087 -2390
rect -2087 -3892 -2029 -3188
rect -2087 -4484 -2075 -3892
rect -2041 -4484 -2029 -3892
rect -2087 -5188 -2029 -4484
rect -29 -3892 29 -3188
rect -29 -4484 -17 -3892
rect 17 -4484 29 -3892
rect -29 -5188 29 -4484
rect 2029 -3892 2087 -3188
rect 2029 -4484 2041 -3892
rect 2075 -4484 2087 -3892
rect 2029 -5188 2087 -4484
<< mvndiffc >>
rect -2075 3892 -2041 4484
rect -17 3892 17 4484
rect 2041 3892 2075 4484
rect -2075 1798 -2041 2390
rect -17 1798 17 2390
rect 2041 1798 2075 2390
rect -2075 -296 -2041 296
rect -17 -296 17 296
rect 2041 -296 2075 296
rect -2075 -2390 -2041 -1798
rect -17 -2390 17 -1798
rect 2041 -2390 2075 -1798
rect -2075 -4484 -2041 -3892
rect -17 -4484 17 -3892
rect 2041 -4484 2075 -3892
<< poly >>
rect -2029 5188 -29 5214
rect 29 5188 2029 5214
rect -2029 3162 -29 3188
rect 29 3162 2029 3188
rect -2029 3094 -29 3120
rect 29 3094 2029 3120
rect -2029 1068 -29 1094
rect 29 1068 2029 1094
rect -2029 1000 -29 1026
rect 29 1000 2029 1026
rect -2029 -1026 -29 -1000
rect 29 -1026 2029 -1000
rect -2029 -1094 -29 -1068
rect 29 -1094 2029 -1068
rect -2029 -3120 -29 -3094
rect 29 -3120 2029 -3094
rect -2029 -3188 -29 -3162
rect 29 -3188 2029 -3162
rect -2029 -5214 -29 -5188
rect 29 -5214 2029 -5188
<< locali >>
rect -2075 4484 -2041 4500
rect -2075 3876 -2041 3892
rect -17 4484 17 4500
rect -17 3876 17 3892
rect 2041 4484 2075 4500
rect 2041 3876 2075 3892
rect -2075 2390 -2041 2406
rect -2075 1782 -2041 1798
rect -17 2390 17 2406
rect -17 1782 17 1798
rect 2041 2390 2075 2406
rect 2041 1782 2075 1798
rect -2075 296 -2041 312
rect -2075 -312 -2041 -296
rect -17 296 17 312
rect -17 -312 17 -296
rect 2041 296 2075 312
rect 2041 -312 2075 -296
rect -2075 -1798 -2041 -1782
rect -2075 -2406 -2041 -2390
rect -17 -1798 17 -1782
rect -17 -2406 17 -2390
rect 2041 -1798 2075 -1782
rect 2041 -2406 2075 -2390
rect -2075 -3892 -2041 -3876
rect -2075 -4500 -2041 -4484
rect -17 -3892 17 -3876
rect -17 -4500 17 -4484
rect 2041 -3892 2075 -3876
rect 2041 -4500 2075 -4484
<< viali >>
rect -2075 3892 -2041 4484
rect -17 3892 17 4484
rect 2041 3892 2075 4484
rect -2075 1798 -2041 2390
rect -17 1798 17 2390
rect 2041 1798 2075 2390
rect -2075 -296 -2041 296
rect -17 -296 17 296
rect 2041 -296 2075 296
rect -2075 -2390 -2041 -1798
rect -17 -2390 17 -1798
rect 2041 -2390 2075 -1798
rect -2075 -4484 -2041 -3892
rect -17 -4484 17 -3892
rect 2041 -4484 2075 -3892
<< metal1 >>
rect -2081 4484 -2035 4496
rect -2081 3892 -2075 4484
rect -2041 3892 -2035 4484
rect -2081 3880 -2035 3892
rect -23 4484 23 4496
rect -23 3892 -17 4484
rect 17 3892 23 4484
rect -23 3880 23 3892
rect 2035 4484 2081 4496
rect 2035 3892 2041 4484
rect 2075 3892 2081 4484
rect 2035 3880 2081 3892
rect -2081 2390 -2035 2402
rect -2081 1798 -2075 2390
rect -2041 1798 -2035 2390
rect -2081 1786 -2035 1798
rect -23 2390 23 2402
rect -23 1798 -17 2390
rect 17 1798 23 2390
rect -23 1786 23 1798
rect 2035 2390 2081 2402
rect 2035 1798 2041 2390
rect 2075 1798 2081 2390
rect 2035 1786 2081 1798
rect -2081 296 -2035 308
rect -2081 -296 -2075 296
rect -2041 -296 -2035 296
rect -2081 -308 -2035 -296
rect -23 296 23 308
rect -23 -296 -17 296
rect 17 -296 23 296
rect -23 -308 23 -296
rect 2035 296 2081 308
rect 2035 -296 2041 296
rect 2075 -296 2081 296
rect 2035 -308 2081 -296
rect -2081 -1798 -2035 -1786
rect -2081 -2390 -2075 -1798
rect -2041 -2390 -2035 -1798
rect -2081 -2402 -2035 -2390
rect -23 -1798 23 -1786
rect -23 -2390 -17 -1798
rect 17 -2390 23 -1798
rect -23 -2402 23 -2390
rect 2035 -1798 2081 -1786
rect 2035 -2390 2041 -1798
rect 2075 -2390 2081 -1798
rect 2035 -2402 2081 -2390
rect -2081 -3892 -2035 -3880
rect -2081 -4484 -2075 -3892
rect -2041 -4484 -2035 -3892
rect -2081 -4496 -2035 -4484
rect -23 -3892 23 -3880
rect -23 -4484 -17 -3892
rect 17 -4484 23 -3892
rect -23 -4496 23 -4484
rect 2035 -3892 2081 -3880
rect 2035 -4484 2041 -3892
rect 2075 -4484 2081 -3892
rect 2035 -4496 2081 -4484
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string parameters w 10 l 10 m 5 nf 2 diffcov 30 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 30 viadrn 30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
