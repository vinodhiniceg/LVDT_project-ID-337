magic
tech sky130A
timestamp 1634141228
<< pwell >>
rect -106 -269 6041 2014
rect -42 -289 5878 -269
<< mvpsubdiff >>
rect -64 1912 5900 2060
rect -38 -128 129 1912
rect 5722 1541 5899 1912
rect 5722 1478 5901 1541
rect 5722 525 5749 1478
rect 5864 525 5901 1478
rect 5722 374 5901 525
rect 5722 -128 5899 374
rect -42 -254 5899 -128
rect -42 -289 5878 -254
<< mvpsubdiffcont >>
rect 5749 525 5864 1478
<< poly >>
rect 692 1856 1227 1885
rect 692 1773 831 1856
rect 1026 1773 1227 1856
rect 692 1736 1227 1773
rect 2731 1719 3101 1883
rect 4578 1847 5047 1864
rect 4578 1762 4724 1847
rect 4848 1762 5047 1847
rect 4578 1744 5047 1762
<< polycont >>
rect 831 1773 1026 1856
rect 4724 1762 4848 1847
<< locali >>
rect 822 1856 1045 1866
rect 822 1773 831 1856
rect 1026 1773 1045 1856
rect 4711 1847 4865 1859
rect 822 1762 1045 1773
rect 847 1641 922 1762
rect 1814 1681 1851 1683
rect 1459 1622 1856 1681
rect 1814 1567 1851 1622
rect 2060 1613 2150 1806
rect 1813 1544 1853 1567
rect 1869 1372 2027 1499
rect 3715 1498 3800 1814
rect 4711 1762 4724 1847
rect 4848 1762 4865 1847
rect 4711 1753 4865 1762
rect 4754 1641 4820 1753
rect 5608 1683 5654 1684
rect 5294 1636 5656 1683
rect 5608 1580 5654 1636
rect 5608 1557 5656 1580
rect 5613 1511 5656 1557
rect 5731 1488 5901 1541
rect 5629 1478 5901 1488
rect 5629 1433 5749 1478
rect 1825 1312 2027 1372
rect 1869 1264 2027 1312
rect 5731 525 5749 1433
rect 5864 525 5901 1478
rect 5731 374 5901 525
<< viali >>
rect 849 1786 992 1847
rect 4748 1776 4821 1832
rect 5749 525 5864 1478
<< metal1 >>
rect 822 1847 1045 1866
rect 822 1786 849 1847
rect 992 1786 1045 1847
rect 822 1762 1045 1786
rect 4711 1832 4865 1859
rect 4711 1776 4748 1832
rect 4821 1776 4865 1832
rect 4711 1753 4865 1776
rect 5731 1478 5901 1541
rect 5731 525 5749 1478
rect 5864 525 5901 1478
rect 5731 374 5901 525
use nmos3355  nmos3355_0 ~/layout test
timestamp 1634132563
transform 1 0 174 0 1 0
box -174 0 1675 1760
use nmos3355  nmos3355_1
timestamp 1634132563
transform 1 0 2071 0 1 1
box -174 0 1675 1760
use nmos3355  nmos3355_2
timestamp 1634132563
transform 1 0 3975 0 1 8
box -174 0 1675 1760
<< labels >>
flabel poly 2856 1807 2856 1807 0 FreeSans 800 0 0 0 g
flabel locali 2079 1738 2079 1738 0 FreeSans 800 0 0 0 d
flabel locali 3737 1754 3737 1754 0 FreeSans 800 0 0 0 s
flabel locali 1918 1422 1918 1422 0 FreeSans 800 0 0 0 sub
<< end >>
