magic
tech sky130A
timestamp 1634117422
<< pwell >>
rect -346 3753 2887 3767
rect -346 3591 2901 3753
rect -339 -164 2901 3591
rect -339 -252 2894 -164
<< mvpsubdiff >>
rect -346 3753 2887 3767
rect -346 3591 2901 3753
rect -339 -76 -82 3591
rect 2644 -76 2901 3591
rect -339 -164 2901 -76
rect -339 -252 2894 -164
<< poly >>
rect 2121 3538 2390 3549
rect 203 3500 479 3506
rect 203 3473 319 3500
rect 362 3473 479 3500
rect 1197 3474 1402 3530
rect 2121 3490 2208 3538
rect 2282 3490 2390 3538
rect 2121 3478 2390 3490
rect 203 3464 479 3473
<< polycont >>
rect 319 3473 362 3500
rect 2208 3490 2282 3538
<< locali >>
rect 2193 3538 2300 3558
rect 311 3500 371 3511
rect 311 3473 319 3500
rect 362 3473 371 3500
rect 2193 3490 2208 3538
rect 2282 3490 2300 3538
rect 2193 3483 2300 3490
rect 311 3464 371 3473
rect 330 3418 351 3464
rect 330 3391 352 3418
rect 331 3320 352 3391
rect 920 3380 974 3410
rect 2245 3320 2276 3483
rect 659 3006 822 3070
rect 1699 2962 1757 3229
rect 2573 3045 2735 3082
rect 1259 -39 1324 72
<< viali >>
rect 326 3477 355 3496
rect 2222 3498 2264 3525
<< metal1 >>
rect 2193 3525 2300 3558
rect 311 3496 371 3511
rect 311 3477 326 3496
rect 355 3477 371 3496
rect 2193 3498 2222 3525
rect 2264 3498 2300 3525
rect 2193 3483 2300 3498
rect 311 3464 371 3477
use nmos33210  nmos33210_2
timestamp 1634112475
transform 1 0 1916 0 1 11
box 0 0 880 3481
use nmos33210  nmos33210_1
timestamp 1634112475
transform 1 0 945 0 1 3
box 0 0 880 3481
use nmos33210  nmos33210_0
timestamp 1634112475
transform 1 0 0 0 1 0
box 0 0 880 3481
<< labels >>
flabel locali 926 3392 926 3392 0 FreeSans 800 0 0 0 d
flabel locali 1286 -24 1286 -24 0 FreeSans 800 0 0 0 s
flabel poly 1270 3505 1270 3505 0 FreeSans 800 0 0 0 g
flabel locali 1730 3132 1730 3132 0 FreeSans 800 0 0 0 sub
<< end >>
