magic
tech sky130A
magscale 1 2
timestamp 1634224850
<< mvnmos >>
rect -1287 1435 -687 2035
rect -629 1435 -29 2035
rect 29 1435 629 2035
rect 687 1435 1287 2035
rect -1287 741 -687 1341
rect -629 741 -29 1341
rect 29 741 629 1341
rect 687 741 1287 1341
rect -1287 47 -687 647
rect -629 47 -29 647
rect 29 47 629 647
rect 687 47 1287 647
rect -1287 -647 -687 -47
rect -629 -647 -29 -47
rect 29 -647 629 -47
rect 687 -647 1287 -47
rect -1287 -1341 -687 -741
rect -629 -1341 -29 -741
rect 29 -1341 629 -741
rect 687 -1341 1287 -741
rect -1287 -2035 -687 -1435
rect -629 -2035 -29 -1435
rect 29 -2035 629 -1435
rect 687 -2035 1287 -1435
<< mvndiff >>
rect -1345 1821 -1287 2035
rect -1345 1649 -1333 1821
rect -1299 1649 -1287 1821
rect -1345 1435 -1287 1649
rect -687 1821 -629 2035
rect -687 1649 -675 1821
rect -641 1649 -629 1821
rect -687 1435 -629 1649
rect -29 1821 29 2035
rect -29 1649 -17 1821
rect 17 1649 29 1821
rect -29 1435 29 1649
rect 629 1821 687 2035
rect 629 1649 641 1821
rect 675 1649 687 1821
rect 629 1435 687 1649
rect 1287 1821 1345 2035
rect 1287 1649 1299 1821
rect 1333 1649 1345 1821
rect 1287 1435 1345 1649
rect -1345 1127 -1287 1341
rect -1345 955 -1333 1127
rect -1299 955 -1287 1127
rect -1345 741 -1287 955
rect -687 1127 -629 1341
rect -687 955 -675 1127
rect -641 955 -629 1127
rect -687 741 -629 955
rect -29 1127 29 1341
rect -29 955 -17 1127
rect 17 955 29 1127
rect -29 741 29 955
rect 629 1127 687 1341
rect 629 955 641 1127
rect 675 955 687 1127
rect 629 741 687 955
rect 1287 1127 1345 1341
rect 1287 955 1299 1127
rect 1333 955 1345 1127
rect 1287 741 1345 955
rect -1345 433 -1287 647
rect -1345 261 -1333 433
rect -1299 261 -1287 433
rect -1345 47 -1287 261
rect -687 433 -629 647
rect -687 261 -675 433
rect -641 261 -629 433
rect -687 47 -629 261
rect -29 433 29 647
rect -29 261 -17 433
rect 17 261 29 433
rect -29 47 29 261
rect 629 433 687 647
rect 629 261 641 433
rect 675 261 687 433
rect 629 47 687 261
rect 1287 433 1345 647
rect 1287 261 1299 433
rect 1333 261 1345 433
rect 1287 47 1345 261
rect -1345 -261 -1287 -47
rect -1345 -433 -1333 -261
rect -1299 -433 -1287 -261
rect -1345 -647 -1287 -433
rect -687 -261 -629 -47
rect -687 -433 -675 -261
rect -641 -433 -629 -261
rect -687 -647 -629 -433
rect -29 -261 29 -47
rect -29 -433 -17 -261
rect 17 -433 29 -261
rect -29 -647 29 -433
rect 629 -261 687 -47
rect 629 -433 641 -261
rect 675 -433 687 -261
rect 629 -647 687 -433
rect 1287 -261 1345 -47
rect 1287 -433 1299 -261
rect 1333 -433 1345 -261
rect 1287 -647 1345 -433
rect -1345 -955 -1287 -741
rect -1345 -1127 -1333 -955
rect -1299 -1127 -1287 -955
rect -1345 -1341 -1287 -1127
rect -687 -955 -629 -741
rect -687 -1127 -675 -955
rect -641 -1127 -629 -955
rect -687 -1341 -629 -1127
rect -29 -955 29 -741
rect -29 -1127 -17 -955
rect 17 -1127 29 -955
rect -29 -1341 29 -1127
rect 629 -955 687 -741
rect 629 -1127 641 -955
rect 675 -1127 687 -955
rect 629 -1341 687 -1127
rect 1287 -955 1345 -741
rect 1287 -1127 1299 -955
rect 1333 -1127 1345 -955
rect 1287 -1341 1345 -1127
rect -1345 -1649 -1287 -1435
rect -1345 -1821 -1333 -1649
rect -1299 -1821 -1287 -1649
rect -1345 -2035 -1287 -1821
rect -687 -1649 -629 -1435
rect -687 -1821 -675 -1649
rect -641 -1821 -629 -1649
rect -687 -2035 -629 -1821
rect -29 -1649 29 -1435
rect -29 -1821 -17 -1649
rect 17 -1821 29 -1649
rect -29 -2035 29 -1821
rect 629 -1649 687 -1435
rect 629 -1821 641 -1649
rect 675 -1821 687 -1649
rect 629 -2035 687 -1821
rect 1287 -1649 1345 -1435
rect 1287 -1821 1299 -1649
rect 1333 -1821 1345 -1649
rect 1287 -2035 1345 -1821
<< mvndiffc >>
rect -1333 1649 -1299 1821
rect -675 1649 -641 1821
rect -17 1649 17 1821
rect 641 1649 675 1821
rect 1299 1649 1333 1821
rect -1333 955 -1299 1127
rect -675 955 -641 1127
rect -17 955 17 1127
rect 641 955 675 1127
rect 1299 955 1333 1127
rect -1333 261 -1299 433
rect -675 261 -641 433
rect -17 261 17 433
rect 641 261 675 433
rect 1299 261 1333 433
rect -1333 -433 -1299 -261
rect -675 -433 -641 -261
rect -17 -433 17 -261
rect 641 -433 675 -261
rect 1299 -433 1333 -261
rect -1333 -1127 -1299 -955
rect -675 -1127 -641 -955
rect -17 -1127 17 -955
rect 641 -1127 675 -955
rect 1299 -1127 1333 -955
rect -1333 -1821 -1299 -1649
rect -675 -1821 -641 -1649
rect -17 -1821 17 -1649
rect 641 -1821 675 -1649
rect 1299 -1821 1333 -1649
<< poly >>
rect -1287 2035 -687 2061
rect -629 2035 -29 2061
rect 29 2035 629 2061
rect 687 2035 1287 2061
rect -1287 1409 -687 1435
rect -629 1409 -29 1435
rect 29 1409 629 1435
rect 687 1409 1287 1435
rect -1287 1341 -687 1367
rect -629 1341 -29 1367
rect 29 1341 629 1367
rect 687 1341 1287 1367
rect -1287 715 -687 741
rect -629 715 -29 741
rect 29 715 629 741
rect 687 715 1287 741
rect -1287 647 -687 673
rect -629 647 -29 673
rect 29 647 629 673
rect 687 647 1287 673
rect -1287 21 -687 47
rect -629 21 -29 47
rect 29 21 629 47
rect 687 21 1287 47
rect -1287 -47 -687 -21
rect -629 -47 -29 -21
rect 29 -47 629 -21
rect 687 -47 1287 -21
rect -1287 -673 -687 -647
rect -629 -673 -29 -647
rect 29 -673 629 -647
rect 687 -673 1287 -647
rect -1287 -741 -687 -715
rect -629 -741 -29 -715
rect 29 -741 629 -715
rect 687 -741 1287 -715
rect -1287 -1367 -687 -1341
rect -629 -1367 -29 -1341
rect 29 -1367 629 -1341
rect 687 -1367 1287 -1341
rect -1287 -1435 -687 -1409
rect -629 -1435 -29 -1409
rect 29 -1435 629 -1409
rect 687 -1435 1287 -1409
rect -1287 -2061 -687 -2035
rect -629 -2061 -29 -2035
rect 29 -2061 629 -2035
rect 687 -2061 1287 -2035
<< locali >>
rect -1333 1821 -1299 1837
rect -1333 1633 -1299 1649
rect -675 1821 -641 1837
rect -675 1633 -641 1649
rect -17 1821 17 1837
rect -17 1633 17 1649
rect 641 1821 675 1837
rect 641 1633 675 1649
rect 1299 1821 1333 1837
rect 1299 1633 1333 1649
rect -1333 1127 -1299 1143
rect -1333 939 -1299 955
rect -675 1127 -641 1143
rect -675 939 -641 955
rect -17 1127 17 1143
rect -17 939 17 955
rect 641 1127 675 1143
rect 641 939 675 955
rect 1299 1127 1333 1143
rect 1299 939 1333 955
rect -1333 433 -1299 449
rect -1333 245 -1299 261
rect -675 433 -641 449
rect -675 245 -641 261
rect -17 433 17 449
rect -17 245 17 261
rect 641 433 675 449
rect 641 245 675 261
rect 1299 433 1333 449
rect 1299 245 1333 261
rect -1333 -261 -1299 -245
rect -1333 -449 -1299 -433
rect -675 -261 -641 -245
rect -675 -449 -641 -433
rect -17 -261 17 -245
rect -17 -449 17 -433
rect 641 -261 675 -245
rect 641 -449 675 -433
rect 1299 -261 1333 -245
rect 1299 -449 1333 -433
rect -1333 -955 -1299 -939
rect -1333 -1143 -1299 -1127
rect -675 -955 -641 -939
rect -675 -1143 -641 -1127
rect -17 -955 17 -939
rect -17 -1143 17 -1127
rect 641 -955 675 -939
rect 641 -1143 675 -1127
rect 1299 -955 1333 -939
rect 1299 -1143 1333 -1127
rect -1333 -1649 -1299 -1633
rect -1333 -1837 -1299 -1821
rect -675 -1649 -641 -1633
rect -675 -1837 -641 -1821
rect -17 -1649 17 -1633
rect -17 -1837 17 -1821
rect 641 -1649 675 -1633
rect 641 -1837 675 -1821
rect 1299 -1649 1333 -1633
rect 1299 -1837 1333 -1821
<< viali >>
rect -1333 1649 -1299 1821
rect -675 1649 -641 1821
rect -17 1649 17 1821
rect 641 1649 675 1821
rect 1299 1649 1333 1821
rect -1333 955 -1299 1127
rect -675 955 -641 1127
rect -17 955 17 1127
rect 641 955 675 1127
rect 1299 955 1333 1127
rect -1333 261 -1299 433
rect -675 261 -641 433
rect -17 261 17 433
rect 641 261 675 433
rect 1299 261 1333 433
rect -1333 -433 -1299 -261
rect -675 -433 -641 -261
rect -17 -433 17 -261
rect 641 -433 675 -261
rect 1299 -433 1333 -261
rect -1333 -1127 -1299 -955
rect -675 -1127 -641 -955
rect -17 -1127 17 -955
rect 641 -1127 675 -955
rect 1299 -1127 1333 -955
rect -1333 -1821 -1299 -1649
rect -675 -1821 -641 -1649
rect -17 -1821 17 -1649
rect 641 -1821 675 -1649
rect 1299 -1821 1333 -1649
<< metal1 >>
rect -1339 1821 -1293 1833
rect -1339 1649 -1333 1821
rect -1299 1649 -1293 1821
rect -1339 1637 -1293 1649
rect -681 1821 -635 1833
rect -681 1649 -675 1821
rect -641 1649 -635 1821
rect -681 1637 -635 1649
rect -23 1821 23 1833
rect -23 1649 -17 1821
rect 17 1649 23 1821
rect -23 1637 23 1649
rect 635 1821 681 1833
rect 635 1649 641 1821
rect 675 1649 681 1821
rect 635 1637 681 1649
rect 1293 1821 1339 1833
rect 1293 1649 1299 1821
rect 1333 1649 1339 1821
rect 1293 1637 1339 1649
rect -1339 1127 -1293 1139
rect -1339 955 -1333 1127
rect -1299 955 -1293 1127
rect -1339 943 -1293 955
rect -681 1127 -635 1139
rect -681 955 -675 1127
rect -641 955 -635 1127
rect -681 943 -635 955
rect -23 1127 23 1139
rect -23 955 -17 1127
rect 17 955 23 1127
rect -23 943 23 955
rect 635 1127 681 1139
rect 635 955 641 1127
rect 675 955 681 1127
rect 635 943 681 955
rect 1293 1127 1339 1139
rect 1293 955 1299 1127
rect 1333 955 1339 1127
rect 1293 943 1339 955
rect -1339 433 -1293 445
rect -1339 261 -1333 433
rect -1299 261 -1293 433
rect -1339 249 -1293 261
rect -681 433 -635 445
rect -681 261 -675 433
rect -641 261 -635 433
rect -681 249 -635 261
rect -23 433 23 445
rect -23 261 -17 433
rect 17 261 23 433
rect -23 249 23 261
rect 635 433 681 445
rect 635 261 641 433
rect 675 261 681 433
rect 635 249 681 261
rect 1293 433 1339 445
rect 1293 261 1299 433
rect 1333 261 1339 433
rect 1293 249 1339 261
rect -1339 -261 -1293 -249
rect -1339 -433 -1333 -261
rect -1299 -433 -1293 -261
rect -1339 -445 -1293 -433
rect -681 -261 -635 -249
rect -681 -433 -675 -261
rect -641 -433 -635 -261
rect -681 -445 -635 -433
rect -23 -261 23 -249
rect -23 -433 -17 -261
rect 17 -433 23 -261
rect -23 -445 23 -433
rect 635 -261 681 -249
rect 635 -433 641 -261
rect 675 -433 681 -261
rect 635 -445 681 -433
rect 1293 -261 1339 -249
rect 1293 -433 1299 -261
rect 1333 -433 1339 -261
rect 1293 -445 1339 -433
rect -1339 -955 -1293 -943
rect -1339 -1127 -1333 -955
rect -1299 -1127 -1293 -955
rect -1339 -1139 -1293 -1127
rect -681 -955 -635 -943
rect -681 -1127 -675 -955
rect -641 -1127 -635 -955
rect -681 -1139 -635 -1127
rect -23 -955 23 -943
rect -23 -1127 -17 -955
rect 17 -1127 23 -955
rect -23 -1139 23 -1127
rect 635 -955 681 -943
rect 635 -1127 641 -955
rect 675 -1127 681 -955
rect 635 -1139 681 -1127
rect 1293 -955 1339 -943
rect 1293 -1127 1299 -955
rect 1333 -1127 1339 -955
rect 1293 -1139 1339 -1127
rect -1339 -1649 -1293 -1637
rect -1339 -1821 -1333 -1649
rect -1299 -1821 -1293 -1649
rect -1339 -1833 -1293 -1821
rect -681 -1649 -635 -1637
rect -681 -1821 -675 -1649
rect -641 -1821 -635 -1649
rect -681 -1833 -635 -1821
rect -23 -1649 23 -1637
rect -23 -1821 -17 -1649
rect 17 -1821 23 -1649
rect -23 -1833 23 -1821
rect 635 -1649 681 -1637
rect 635 -1821 641 -1649
rect 675 -1821 681 -1649
rect 635 -1833 681 -1821
rect 1293 -1649 1339 -1637
rect 1293 -1821 1299 -1649
rect 1333 -1821 1339 -1649
rect 1293 -1833 1339 -1821
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string parameters w 3 l 3 m 6 nf 4 diffcov 30 polycov 30 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 30 viadrn 30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
