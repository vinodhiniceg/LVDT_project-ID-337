magic
tech sky130A
timestamp 1634274673
<< nwell >>
rect -26 12197 5807 12361
rect -26 12100 5814 12197
rect -11 11712 5814 12100
rect -18 -573 5814 32
<< mvnsubdiff >>
rect 146 12100 5754 12167
rect 146 11943 5762 12100
rect 161 11591 318 11943
rect 5597 11592 5762 11943
rect 161 11517 321 11591
rect 175 10606 321 11517
rect 179 7120 313 10606
rect 179 7116 317 7120
rect 183 256 317 7116
rect 176 117 317 256
rect 5612 219 5762 11592
rect 176 -102 310 117
rect 5612 -102 5777 219
rect 161 -319 5777 -102
rect 161 -334 5747 -319
<< poly >>
rect 4692 11880 5361 11897
rect 816 11833 1401 11854
rect 816 11770 998 11833
rect 1142 11770 1401 11833
rect 816 11747 1401 11770
rect 4692 11788 4898 11880
rect 5121 11788 5361 11880
rect 4692 11745 5361 11788
<< polycont >>
rect 998 11770 1142 11833
rect 4898 11788 5121 11880
<< locali >>
rect 4860 11880 5160 11889
rect 985 11833 1157 11854
rect 985 11770 998 11833
rect 1142 11770 1157 11833
rect 985 11749 1157 11770
rect 4860 11788 4898 11880
rect 5121 11788 5160 11880
rect 4860 11768 5160 11788
rect 1017 11638 1080 11749
rect 1341 11582 1403 11685
rect 4960 11633 5027 11768
rect 5201 11573 5248 11687
rect 4102 10975 4233 11013
rect 252 10900 361 10947
<< viali >>
rect 1019 11775 1122 11826
rect 4935 11796 5080 11871
<< metal1 >>
rect 4860 11871 5160 11889
rect 985 11826 1157 11854
rect 985 11775 1019 11826
rect 1122 11775 1157 11826
rect 985 11749 1157 11775
rect 4860 11796 4935 11871
rect 5080 11796 5160 11871
rect 4860 11768 5160 11796
use pmos33431  pmos33431_2
timestamp 1634273660
transform 1 0 3966 0 1 8
box -109 -11 1850 11807
use pmos33431  pmos33431_1
timestamp 1634273660
transform 1 0 2041 0 1 1
box -109 -11 1850 11807
use pmos33431  pmos33431_0
timestamp 1634273660
transform 1 0 109 0 1 11
box -109 -11 1850 11807
<< end >>
