magic
tech sky130A
magscale 1 2
timestamp 1634929433
<< nwell >>
rect -1632 3426 738 3622
rect -1642 3382 738 3426
rect -1642 1848 734 3382
rect -1642 -88 1654 1848
<< pwell >>
rect -2456 5006 -1748 5010
rect -2684 4986 -1692 5006
rect -2684 -134 -1674 4986
rect 1022 3556 2004 3562
rect 850 3548 2004 3556
rect 2256 3548 2882 3572
rect 850 1908 2882 3548
rect 1684 -102 2882 1908
rect 2256 -124 2882 -102
rect -2456 -144 -1674 -134
<< mvpsubdiff >>
rect -2584 2594 -2450 2676
rect -2584 450 -2560 2594
rect -2482 450 -2450 2594
rect 2432 1222 2602 1280
rect -2584 328 -2450 450
rect 2432 190 2456 1222
rect 2554 190 2602 1222
rect 2432 116 2602 190
<< mvnsubdiff >>
rect -398 3376 -124 3426
rect -398 3054 -378 3376
rect -196 3054 -124 3376
rect -398 3004 -124 3054
rect 1480 960 1576 994
rect 1480 238 1492 960
rect 1564 238 1576 960
rect 1480 210 1576 238
<< mvpsubdiffcont >>
rect -2560 450 -2482 2594
rect 2456 190 2554 1222
<< mvnsubdiffcont >>
rect -378 3054 -196 3376
rect 1492 238 1564 960
<< poly >>
rect -2262 5024 -1908 5090
rect -2262 4922 -2180 5024
rect -2024 4922 -1908 5024
rect -2262 4914 -1908 4922
rect 1238 3430 1542 3690
rect 190 3312 494 3430
rect -1364 2334 -466 2378
rect -268 1586 -200 1590
rect -268 1584 440 1586
rect -268 1514 1092 1584
rect -268 1496 -200 1514
rect 370 1512 1092 1514
rect -532 1490 -200 1496
rect -536 1452 -200 1490
rect -268 1442 -200 1452
rect 126 -6 282 34
rect 126 -86 160 -6
rect 236 -86 282 -6
rect 126 -122 282 -86
<< polycont >>
rect -2180 4922 -2024 5024
rect 1940 1498 2086 1566
rect 160 -86 236 -6
<< locali >>
rect -2204 5024 -1988 5048
rect -2204 4922 -2180 5024
rect -2024 4922 -1988 5024
rect -2204 4900 -1988 4922
rect -408 3376 -134 3416
rect -408 3054 -378 3376
rect -196 3054 -134 3376
rect -408 3000 -134 3054
rect -2584 2594 -2450 2676
rect -2584 450 -2560 2594
rect -2482 450 -2450 2594
rect 1916 1566 2118 1578
rect 1916 1498 1940 1566
rect 2086 1498 2118 1566
rect 1916 1478 2118 1498
rect 2432 1222 2602 1280
rect -2584 328 -2450 450
rect 1480 960 1576 994
rect 1480 238 1492 960
rect 1564 238 1576 960
rect 1480 210 1576 238
rect 2432 190 2456 1222
rect 2554 190 2602 1222
rect 2432 116 2602 190
rect 144 -6 262 22
rect 144 -86 160 -6
rect 236 -86 262 -6
rect 144 -104 262 -86
<< viali >>
rect -2180 4922 -2024 5024
rect -378 3054 -196 3376
rect -2554 528 -2486 2562
rect 1960 1506 2062 1558
rect 1498 268 1552 922
rect 2456 190 2554 1222
rect 160 -86 236 -6
<< metal1 >>
rect -2204 5024 -1988 5048
rect -1770 5024 -1760 5082
rect -2204 4922 -2180 5024
rect -2024 4958 -1760 5024
rect -2024 4922 -1988 4958
rect -1770 4928 -1760 4958
rect -1590 4928 -1580 5082
rect -2204 4900 -1988 4922
rect -2374 4830 -1792 4844
rect -2642 4686 -2632 4810
rect -2528 4780 -2518 4810
rect -2376 4808 -1792 4830
rect -2376 4780 -2326 4808
rect -2528 4742 -2326 4780
rect -2528 4732 -2330 4742
rect -1858 4734 -1812 4808
rect -1514 4750 2742 5148
rect -1430 4738 2742 4750
rect -2528 4702 -2338 4732
rect -2528 4686 -2518 4702
rect -1430 2872 -1258 4738
rect -328 3416 -250 4738
rect 42 4732 88 4738
rect 956 4732 1004 4738
rect 1048 3814 1058 3954
rect 1208 3814 1218 3954
rect -408 3376 -134 3416
rect -408 3054 -378 3376
rect -196 3054 -134 3376
rect 1092 3220 1146 3814
rect 28 3180 86 3220
rect 28 3114 94 3180
rect 1612 3086 1708 3148
rect -408 3000 -134 3054
rect -410 2774 -374 2866
rect 36 2774 84 2866
rect -2584 2562 -2450 2676
rect -2584 528 -2554 2562
rect -2486 528 -2450 2562
rect -718 2434 -708 2632
rect -606 2434 -596 2632
rect -30 2466 -20 2660
rect 148 2466 158 2660
rect -424 2380 -370 2434
rect 62 2380 104 2434
rect 312 1846 366 1974
rect 1352 1944 1394 2092
rect 1352 1878 2466 1944
rect 1494 1846 1550 1878
rect 312 1792 1558 1846
rect 1494 1784 1550 1792
rect 1676 1486 1686 1600
rect 1758 1550 1768 1600
rect 1916 1558 2118 1578
rect 1916 1550 1960 1558
rect 1758 1506 1960 1550
rect 2062 1506 2118 1558
rect 1758 1504 2118 1506
rect 1758 1486 1768 1504
rect 1916 1478 2118 1504
rect 572 1422 908 1424
rect 1494 1422 1560 1452
rect 554 1390 1560 1422
rect 554 1382 908 1390
rect 572 1378 908 1382
rect 874 1324 908 1378
rect 1466 1360 1560 1390
rect 2012 1386 2042 1478
rect -424 1176 106 1216
rect 1494 994 1560 1360
rect 2432 1222 2602 1280
rect -2584 328 -2450 528
rect 1480 922 1576 994
rect -2558 -214 -2490 328
rect 1480 268 1498 922
rect 1552 268 1576 922
rect 2432 464 2456 1222
rect -2112 -214 -2068 58
rect 144 -2 262 22
rect 308 -2 378 178
rect 144 -6 378 -2
rect 144 -86 160 -6
rect 236 -24 378 -6
rect 1080 60 1182 212
rect 1480 210 1576 268
rect 2426 190 2456 464
rect 2554 190 2602 1222
rect 1720 60 1810 166
rect 1080 -16 1810 60
rect 1720 -18 1810 -16
rect 236 -50 366 -24
rect 236 -86 262 -50
rect 144 -104 262 -86
rect 2000 -214 2052 178
rect 2426 116 2602 190
rect 2426 -214 2588 116
rect -2558 -630 2676 -214
<< via1 >>
rect -1760 4928 -1590 5082
rect -2632 4686 -2528 4810
rect 1058 3814 1208 3954
rect -708 2434 -606 2632
rect -20 2466 148 2660
rect 1686 1486 1758 1600
<< metal2 >>
rect -1760 5082 -1590 5092
rect -1760 4918 -1590 4928
rect -2632 4810 -2528 4820
rect -2632 4676 -2528 4686
rect -1668 1558 -1596 4918
rect 1058 3954 1208 3964
rect 1058 3804 1208 3814
rect -20 2660 148 2670
rect -708 2632 -606 2642
rect -606 2516 -20 2562
rect -20 2456 148 2466
rect -708 2424 -606 2434
rect 1686 1600 1758 1610
rect -1670 1498 1686 1558
rect -1668 1480 -1596 1498
rect 1686 1476 1758 1486
<< via2 >>
rect -2632 4686 -2528 4810
rect 1058 3814 1208 3954
<< metal3 >>
rect -2642 4810 -2518 4815
rect -2642 4686 -2632 4810
rect -2528 4686 -2518 4810
rect -2642 4681 -2518 4686
rect -2588 4598 -2528 4681
rect 114 4598 912 4600
rect 1084 4598 1158 4602
rect -2590 4530 1158 4598
rect 114 4528 912 4530
rect 1084 3959 1158 4530
rect 1048 3954 1218 3959
rect 1048 3814 1058 3954
rect 1208 3814 1218 3954
rect 1048 3809 1218 3814
use nmos1125  nmos1125_0
timestamp 1634907805
transform 1 0 1746 0 1 8
box -16 0 586 1582
use pmos1125  pmos1125_1
timestamp 1634908039
transform 1 0 802 0 1 -16
box -30 -4 680 1566
use pmos1125  pmos1125_0
timestamp 1634908039
transform 1 0 14 0 1 -14
box -30 -4 680 1566
use pmos1125  pmos1125_2
timestamp 1634908039
transform 1 0 14 0 1 1786
box -30 -4 680 1566
use pmos11410  pmos11410_0 ~/Desktop/Layout documents/layout/mag files
timestamp 1634908693
transform 1 0 -1498 0 1 -12
box -42 -38 1212 3002
use nmos1125  nmos1125_1
timestamp 1634907805
transform 1 0 1088 0 1 1932
box -16 0 586 1582
use nmos11217  nmos11217_0 ~/Desktop/Layout documents/layout/mag files
timestamp 1634908262
transform 1 0 -2360 0 1 -112
box -14 20 560 5088
<< labels >>
flabel metal1 -612 4962 -612 4962 0 FreeSans 1600 0 0 0 vdda
flabel metal1 332 4 332 4 0 FreeSans 1600 0 0 0 Iin
flabel metal1 2208 1902 2208 1904 0 FreeSans 1600 0 0 0 vc
flabel poly 1326 3494 1326 3494 0 FreeSans 1600 0 0 0 out2
flabel poly 282 3362 282 3362 0 FreeSans 1600 0 0 0 out1
flabel metal3 448 4556 448 4556 0 FreeSans 1600 0 0 0 nc
flabel metal2 -248 2538 -248 2538 0 FreeSans 1600 0 0 0 pc
flabel metal1 1832 1526 1832 1526 0 FreeSans 1600 0 0 0 dg
flabel metal1 -2098 -144 -2098 -144 0 FreeSans 1600 0 0 0 vssa
<< end >>
