magic
tech sky130A
magscale 1 2
timestamp 1634616517
<< mvnmos >>
rect -287 47 -187 247
rect -129 47 -29 247
rect 29 47 129 247
rect 187 47 287 247
rect -287 -247 -187 -47
rect -129 -247 -29 -47
rect 29 -247 129 -47
rect 187 -247 287 -47
<< mvndiff >>
rect -345 173 -287 247
rect -345 121 -333 173
rect -299 121 -287 173
rect -345 47 -287 121
rect -187 173 -129 247
rect -187 121 -175 173
rect -141 121 -129 173
rect -187 47 -129 121
rect -29 173 29 247
rect -29 121 -17 173
rect 17 121 29 173
rect -29 47 29 121
rect 129 173 187 247
rect 129 121 141 173
rect 175 121 187 173
rect 129 47 187 121
rect 287 173 345 247
rect 287 121 299 173
rect 333 121 345 173
rect 287 47 345 121
rect -345 -121 -287 -47
rect -345 -173 -333 -121
rect -299 -173 -287 -121
rect -345 -247 -287 -173
rect -187 -121 -129 -47
rect -187 -173 -175 -121
rect -141 -173 -129 -121
rect -187 -247 -129 -173
rect -29 -121 29 -47
rect -29 -173 -17 -121
rect 17 -173 29 -121
rect -29 -247 29 -173
rect 129 -121 187 -47
rect 129 -173 141 -121
rect 175 -173 187 -121
rect 129 -247 187 -173
rect 287 -121 345 -47
rect 287 -173 299 -121
rect 333 -173 345 -121
rect 287 -247 345 -173
<< mvndiffc >>
rect -333 121 -299 173
rect -175 121 -141 173
rect -17 121 17 173
rect 141 121 175 173
rect 299 121 333 173
rect -333 -173 -299 -121
rect -175 -173 -141 -121
rect -17 -173 17 -121
rect 141 -173 175 -121
rect 299 -173 333 -121
<< poly >>
rect -287 247 -187 273
rect -129 247 -29 273
rect 29 247 129 273
rect 187 247 287 273
rect -287 21 -187 47
rect -129 21 -29 47
rect 29 21 129 47
rect 187 21 287 47
rect -287 -47 -187 -21
rect -129 -47 -29 -21
rect 29 -47 129 -21
rect 187 -47 287 -21
rect -287 -273 -187 -247
rect -129 -273 -29 -247
rect 29 -273 129 -247
rect 187 -273 287 -247
<< locali >>
rect -333 173 -299 189
rect -333 105 -299 121
rect -175 173 -141 189
rect -175 105 -141 121
rect -17 173 17 189
rect -17 105 17 121
rect 141 173 175 189
rect 141 105 175 121
rect 299 173 333 189
rect 299 105 333 121
rect -333 -121 -299 -105
rect -333 -189 -299 -173
rect -175 -121 -141 -105
rect -175 -189 -141 -173
rect -17 -121 17 -105
rect -17 -189 17 -173
rect 141 -121 175 -105
rect 141 -189 175 -173
rect 299 -121 333 -105
rect 299 -189 333 -173
<< viali >>
rect -333 121 -299 173
rect -175 121 -141 173
rect -17 121 17 173
rect 141 121 175 173
rect 299 121 333 173
rect -333 -173 -299 -121
rect -175 -173 -141 -121
rect -17 -173 17 -121
rect 141 -173 175 -121
rect 299 -173 333 -121
<< metal1 >>
rect -339 173 -293 185
rect -339 121 -333 173
rect -299 121 -293 173
rect -339 109 -293 121
rect -181 173 -135 185
rect -181 121 -175 173
rect -141 121 -135 173
rect -181 109 -135 121
rect -23 173 23 185
rect -23 121 -17 173
rect 17 121 23 173
rect -23 109 23 121
rect 135 173 181 185
rect 135 121 141 173
rect 175 121 181 173
rect 135 109 181 121
rect 293 173 339 185
rect 293 121 299 173
rect 333 121 339 173
rect 293 109 339 121
rect -339 -121 -293 -109
rect -339 -173 -333 -121
rect -299 -173 -293 -121
rect -339 -185 -293 -173
rect -181 -121 -135 -109
rect -181 -173 -175 -121
rect -141 -173 -135 -121
rect -181 -185 -135 -173
rect -23 -121 23 -109
rect -23 -173 -17 -121
rect 17 -173 23 -121
rect -23 -185 23 -173
rect 135 -121 181 -109
rect 135 -173 141 -121
rect 175 -173 181 -121
rect 135 -185 181 -173
rect 293 -121 339 -109
rect 293 -173 299 -121
rect 333 -173 339 -121
rect 293 -185 339 -173
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string parameters w 1 l 0.50 m 2 nf 4 diffcov 30 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 30 viadrn 30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
