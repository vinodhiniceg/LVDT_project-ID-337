magic
tech sky130A
timestamp 1634181701
<< error_s >>
rect 4043 7614 4072 7914
rect 4043 7267 4072 7567
rect 4043 6920 4072 7220
rect 4043 6573 4072 6873
rect 4043 6226 4072 6526
rect 4043 5603 4072 5903
rect 4043 5256 4072 5556
rect 4043 4909 4072 5209
rect 4043 4562 4072 4862
rect 4043 4215 4072 4515
rect 1785 3922 1786 3937
rect 3883 3924 3884 3926
rect 4043 3592 4072 3892
rect 4043 3245 4072 3545
rect 4043 2898 4072 3198
rect 4043 2551 4072 2851
rect 4043 2204 4072 2504
rect 4043 1595 4072 1895
rect 4043 1248 4072 1548
rect 4043 901 4072 1201
rect 4043 554 4072 854
rect 4043 207 4072 507
<< nwell >>
rect -113 7890 4688 8286
rect -113 7841 1644 7890
rect 2391 7841 4688 7890
rect -113 -50 4688 7841
<< poly >>
rect 1607 7952 2666 8053
rect 466 5929 583 6226
rect 695 5927 812 6224
rect 1060 5931 1177 6228
rect 1361 5927 1478 6224
rect 1647 5925 1764 6222
rect 2570 5938 2688 6222
rect 2831 5938 2949 6222
rect 3156 5938 3274 6222
rect 3450 5940 3568 6224
rect 3751 5938 3869 6222
rect 461 3922 578 4219
rect 716 3920 833 4217
rect 1052 3926 1169 4223
rect 1373 3922 1490 4219
rect 1669 3922 1786 4219
rect 2570 3926 2688 4210
rect 2836 3928 2954 4212
rect 3182 3928 3300 4212
rect 3503 3924 3621 4208
rect 3766 3924 3884 4208
rect 463 1914 580 2211
rect 716 1918 833 2215
rect 1055 1916 1172 2213
rect 1356 1918 1473 2215
rect 1657 1912 1774 2209
rect 2568 1917 2686 2201
rect 2816 1923 2934 2207
rect 3156 1915 3274 2199
rect 3503 1917 3621 2201
rect 3758 1917 3876 2201
<< locali >>
rect 1617 7885 2423 7905
rect 1617 7862 2498 7885
rect 1622 7844 1644 7862
rect 2391 7844 2498 7862
rect 297 347 323 7772
rect 1940 325 1966 7750
rect 2398 355 2424 7780
rect 4040 347 4066 7772
rect 1932 220 2808 261
use pmos3355  pmos3355_0 ~/layout test
timestamp 1634178975
transform 1 0 281 0 1 180
box -281 -180 1875 1835
use pmos3355  pmos3355_1
timestamp 1634178975
transform 1 0 282 0 1 2184
box -281 -180 1875 1835
use pmos3355  pmos3355_2
timestamp 1634178975
transform 1 0 282 0 1 4190
box -281 -180 1875 1835
use pmos3355  pmos3355_3
timestamp 1634178975
transform 1 0 282 0 1 6195
box -281 -180 1875 1835
use pmos3355  pmos3355_4
timestamp 1634178975
transform 1 0 2380 0 1 176
box -281 -180 1875 1835
use pmos3355  pmos3355_5
timestamp 1634178975
transform 1 0 2380 0 1 2173
box -281 -180 1875 1835
use pmos3355  pmos3355_6
timestamp 1634178975
transform 1 0 2380 0 1 4184
box -281 -180 1875 1835
use pmos3355  pmos3355_7
timestamp 1634178975
transform 1 0 2380 0 1 6195
box -281 -180 1875 1835
<< end >>
