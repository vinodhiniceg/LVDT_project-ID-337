magic
tech sky130A
magscale 1 2
timestamp 1634629898
<< nwell >>
rect -352 592 5832 960
rect -352 488 2770 592
rect 2820 554 5832 592
rect 2854 514 5832 554
rect 2820 488 5832 514
rect -352 462 2772 488
rect 2776 462 5832 488
rect -352 -250 5832 462
rect -356 -444 5832 -250
rect -356 -1266 538 -444
rect -356 -1280 236 -1266
rect -356 -1380 262 -1280
rect 268 -1380 538 -1266
rect -356 -1500 538 -1380
rect 4940 -1490 5832 -444
<< pwell >>
rect 608 -1524 4866 -482
<< mvpsubdiff >>
rect 628 -646 806 -562
rect 628 -1392 648 -646
rect 776 -1392 806 -646
rect 4664 -636 4848 -536
rect 628 -1456 806 -1392
rect 4664 -1386 4690 -636
rect 4818 -1386 4848 -636
rect 4664 -1436 4848 -1386
<< mvnsubdiff >>
rect 5338 602 5512 658
rect -202 538 -54 600
rect -202 116 -178 538
rect -86 116 -54 538
rect -202 28 -54 116
rect 5338 66 5370 602
rect 5474 66 5512 602
rect 5338 -6 5512 66
<< mvpsubdiffcont >>
rect 648 -1392 776 -646
rect 4690 -1386 4818 -636
<< mvnsubdiffcont >>
rect -178 116 -86 538
rect 5370 66 5474 602
<< poly >>
rect 1256 870 4862 876
rect 320 838 4862 870
rect 316 776 4862 838
rect 316 616 410 776
rect 1256 772 4862 776
rect 1280 608 1362 772
rect 3878 762 4862 772
rect 3878 728 4858 762
rect 3878 624 3974 728
rect 4764 602 4858 728
rect 2260 20 2360 70
rect 2260 -30 2280 20
rect 2334 -30 2360 20
rect 2260 -70 2360 -30
rect 2830 -2 2924 62
rect 2830 -42 2852 -2
rect 2896 -42 2924 -2
rect 3706 38 3800 72
rect 3706 -10 3724 38
rect 3780 -10 3800 38
rect 3706 -34 3800 -10
rect 2830 -86 2924 -42
rect 3736 -498 5308 -484
rect 1942 -510 5308 -498
rect 1940 -524 5308 -510
rect 1940 -536 3774 -524
rect 1940 -618 1976 -536
rect 120 -1558 176 -1318
rect 2650 -844 2780 -810
rect 2650 -896 2680 -844
rect 2734 -896 2780 -844
rect 2650 -930 2780 -896
rect 1250 -1142 1424 -1118
rect 1250 -1182 1284 -1142
rect 1382 -1182 1424 -1142
rect 1250 -1214 1424 -1182
rect 4172 -1122 4334 -1096
rect 4172 -1204 4202 -1122
rect 4304 -1204 4334 -1122
rect 4172 -1230 4334 -1204
rect 5262 -756 5308 -524
rect 7530 -1010 7620 -992
rect 7530 -1098 7544 -1010
rect 7604 -1098 7620 -1010
rect 7530 -1130 7620 -1098
rect 8342 -1008 8426 -982
rect 8342 -1080 8358 -1008
rect 8404 -1080 8426 -1008
rect 8342 -1118 8426 -1080
rect 3394 -1558 3436 -1476
rect 120 -1588 3436 -1558
rect 120 -1590 3432 -1588
<< polycont >>
rect 2280 -30 2334 20
rect 2852 -42 2896 -2
rect 3724 -10 3780 38
rect 2680 -896 2734 -844
rect 1284 -1182 1382 -1142
rect 4202 -1204 4304 -1122
rect 7544 -1098 7604 -1010
rect 8358 -1080 8404 -1008
<< locali >>
rect 5338 602 5512 658
rect -202 538 -54 600
rect -202 116 -178 538
rect -86 116 -54 538
rect -202 28 -54 116
rect 5338 66 5370 602
rect 5474 66 5512 602
rect 3714 38 3796 60
rect 2264 20 2358 30
rect 2264 -30 2280 20
rect 2334 -30 2358 20
rect 2264 -46 2358 -30
rect 2832 -2 2918 10
rect 2832 -42 2852 -2
rect 2896 -42 2918 -2
rect 3714 -10 3724 38
rect 3780 -10 3796 38
rect 5338 -6 5512 66
rect 3714 -26 3796 -10
rect 2832 -54 2918 -42
rect -1408 -310 -1296 -262
rect -1154 -324 -1008 -252
rect 6410 -238 6722 -156
rect 6968 -170 7136 -168
rect 6842 -178 7136 -170
rect 6842 -226 7138 -178
rect 7684 -200 8354 -158
rect 6410 -328 6466 -238
rect 628 -646 806 -562
rect 628 -1302 648 -646
rect 776 -1302 806 -646
rect 4664 -636 4848 -536
rect 2664 -844 2760 -826
rect 2664 -896 2680 -844
rect 2734 -896 2760 -844
rect 2664 -910 2760 -896
rect 4184 -1122 4322 -1108
rect 1266 -1142 1400 -1134
rect 1266 -1182 1284 -1142
rect 1382 -1182 1400 -1142
rect 1266 -1196 1400 -1182
rect 4184 -1204 4202 -1122
rect 4304 -1204 4322 -1122
rect 4184 -1218 4322 -1204
rect 628 -1400 640 -1302
rect 786 -1400 806 -1302
rect 628 -1456 806 -1400
rect 4664 -1386 4690 -636
rect 4818 -1386 4848 -636
rect 7058 -1012 7138 -226
rect 7952 -268 7998 -200
rect 8502 -216 8654 -180
rect 7530 -1010 7620 -992
rect 7530 -1012 7544 -1010
rect 7058 -1050 7544 -1012
rect 7058 -1052 7138 -1050
rect 7530 -1098 7544 -1050
rect 7604 -1098 7620 -1010
rect 7530 -1130 7620 -1098
rect 8342 -1008 8426 -982
rect 8342 -1080 8358 -1008
rect 8404 -1080 8426 -1008
rect 8342 -1118 8426 -1080
rect 4664 -1436 4848 -1386
<< viali >>
rect -170 142 -92 526
rect 5386 124 5444 564
rect 2284 -20 2334 16
rect 2856 -36 2894 -2
rect 3724 -10 3780 38
rect -1544 -324 -1408 -244
rect -1008 -400 -882 -230
rect 7442 -220 7516 -130
rect 6366 -464 6508 -328
rect -1116 -804 -1002 -744
rect 658 -1302 770 -704
rect 2680 -896 2734 -844
rect 1284 -1182 1382 -1142
rect 4202 -1204 4304 -1122
rect 640 -1392 648 -1302
rect 648 -1392 776 -1302
rect 776 -1392 786 -1302
rect 640 -1400 786 -1392
rect 4714 -1302 4804 -690
rect 8654 -246 8716 -176
rect 7938 -332 8014 -268
rect 7544 -1098 7604 -1010
rect 8358 -1080 8404 -1008
<< metal1 >>
rect -338 1060 5960 1224
rect -202 600 -60 1060
rect -202 526 -54 600
rect -202 242 -170 526
rect -1136 188 -170 242
rect -1140 172 -170 188
rect -1140 66 -1112 172
rect -202 142 -170 172
rect -92 142 -54 526
rect 80 490 130 1060
rect 1618 492 1668 1060
rect 1890 470 1940 1060
rect 2820 554 2822 578
rect 2820 488 2822 514
rect 2776 462 2822 488
rect 3406 480 3454 1060
rect 3650 490 3700 1060
rect 5150 484 5200 1060
rect 5366 658 5508 1060
rect 5338 564 5512 658
rect -202 28 -54 142
rect 230 -184 286 192
rect 1154 -114 1188 186
rect 5338 124 5386 564
rect 5444 312 5512 564
rect 5444 276 6670 312
rect 6838 276 7536 318
rect 7692 284 8634 326
rect 8180 280 8544 284
rect 5444 256 6676 276
rect 5444 124 5512 256
rect 6640 168 6676 256
rect 7478 184 7526 276
rect 8496 174 8544 280
rect 1478 90 2102 118
rect 2348 104 2676 118
rect 2348 86 2678 104
rect 2264 16 2358 30
rect 2264 -20 2284 16
rect 2334 -20 2358 16
rect 2264 -46 2358 -20
rect 2636 -4 2678 86
rect 2832 -2 2918 10
rect 2832 -4 2856 -2
rect 2636 -36 2856 -4
rect 2894 -36 2918 -2
rect 2636 -40 2918 -36
rect 1272 -114 1282 -52
rect 1152 -170 1282 -114
rect -1014 -230 -876 -218
rect -1556 -244 -1396 -238
rect -1556 -324 -1544 -244
rect -1408 -324 -1396 -244
rect -1556 -330 -1396 -324
rect -1528 -634 -1472 -330
rect -1018 -400 -1008 -230
rect -882 -400 -872 -230
rect -1014 -412 -876 -400
rect -1576 -688 -1566 -634
rect -1440 -688 -1430 -634
rect -1116 -738 -1088 -538
rect 228 -638 290 -184
rect 1154 -244 1188 -170
rect 1272 -222 1282 -170
rect 1396 -222 1406 -52
rect 2282 -150 2330 -46
rect 2832 -54 2918 -40
rect 2994 -150 3030 110
rect 3290 108 3866 118
rect 3290 90 3888 108
rect 3714 38 3796 60
rect 3714 6 3724 38
rect 3704 -10 3724 6
rect 3780 -10 3796 38
rect 3704 -26 3796 -10
rect 3704 -54 3788 -26
rect 2282 -182 3032 -150
rect 1006 -372 1016 -244
rect 1170 -372 1188 -244
rect 2690 -328 2734 -316
rect 3704 -328 3758 -54
rect 348 -638 358 -604
rect 216 -694 358 -638
rect -1128 -744 -990 -738
rect -1128 -804 -1116 -744
rect -1002 -804 -990 -744
rect -1128 -810 -990 -804
rect 228 -844 290 -694
rect 348 -716 358 -694
rect 530 -716 540 -604
rect 628 -704 806 -562
rect 236 -1302 256 -1232
rect 628 -1302 658 -704
rect 770 -1302 806 -704
rect 1154 -1290 1188 -372
rect 1268 -424 1278 -340
rect 1386 -424 1396 -340
rect 2690 -374 3758 -328
rect 1302 -1134 1354 -424
rect 1462 -728 1472 -614
rect 1582 -658 1592 -614
rect 1582 -728 1692 -658
rect 2690 -826 2734 -374
rect 3804 -414 3814 -356
rect 3896 -366 3906 -356
rect 3938 -358 3980 104
rect 4178 -166 4188 -78
rect 4338 -166 4348 -78
rect 4870 -154 4914 118
rect 5338 -6 5512 124
rect 7436 -130 7522 -118
rect 5488 -154 5534 -150
rect 4014 -358 4024 -340
rect 3938 -366 4024 -358
rect 3896 -394 4024 -366
rect 3896 -414 3906 -394
rect 3938 -416 4024 -394
rect 3800 -712 3810 -656
rect 3886 -712 3896 -656
rect 2664 -844 2760 -826
rect 2664 -896 2680 -844
rect 2734 -896 2760 -844
rect 2664 -910 2760 -896
rect 1266 -1142 1400 -1134
rect 1266 -1182 1284 -1142
rect 1382 -1182 1400 -1142
rect 1266 -1196 1400 -1182
rect 3938 -1290 3980 -416
rect 4014 -432 4024 -416
rect 4142 -432 4152 -340
rect 4224 -1108 4270 -166
rect 4870 -184 5536 -154
rect 4664 -690 4848 -536
rect 5488 -646 5534 -184
rect 7432 -220 7442 -130
rect 7516 -220 7526 -130
rect 8648 -176 8722 -164
rect 7436 -232 7522 -220
rect 8644 -246 8654 -176
rect 8716 -246 8726 -176
rect 8648 -258 8722 -246
rect 7926 -268 8026 -262
rect 6354 -328 6520 -322
rect 6354 -464 6366 -328
rect 6508 -464 6520 -328
rect 7926 -332 7938 -268
rect 8014 -332 8026 -268
rect 7926 -338 8026 -332
rect 6354 -470 6520 -464
rect 6640 -530 6676 -444
rect 7472 -514 7500 -416
rect 4184 -1122 4322 -1108
rect 4184 -1204 4202 -1122
rect 4304 -1204 4322 -1122
rect 4184 -1218 4322 -1204
rect 236 -1444 266 -1302
rect 628 -1400 640 -1302
rect 786 -1400 806 -1302
rect 4664 -1302 4714 -690
rect 4804 -1302 4848 -690
rect 5414 -716 5424 -646
rect 5516 -716 5534 -646
rect 6624 -556 6676 -530
rect 6624 -682 6670 -556
rect 6850 -566 7512 -522
rect 7692 -524 8198 -522
rect 8356 -524 8404 -430
rect 8478 -524 8634 -522
rect 7692 -566 8634 -524
rect 8192 -568 8506 -566
rect 5488 -826 5534 -716
rect 6578 -752 6588 -682
rect 6668 -752 6678 -682
rect 7414 -750 7424 -678
rect 7544 -750 7554 -678
rect 7466 -1232 7502 -750
rect 8234 -774 8244 -638
rect 8338 -774 8348 -638
rect 7530 -1010 7620 -992
rect 7530 -1098 7544 -1010
rect 7604 -1098 7620 -1010
rect 7530 -1130 7620 -1098
rect 8280 -1204 8308 -774
rect 8342 -1008 8426 -982
rect 8342 -1080 8358 -1008
rect 8404 -1022 8426 -1008
rect 8628 -1022 8638 -960
rect 8404 -1064 8638 -1022
rect 8404 -1080 8426 -1064
rect 8342 -1118 8426 -1080
rect 8628 -1116 8638 -1064
rect 8814 -1116 8824 -960
rect 8280 -1230 8306 -1204
rect 8280 -1234 8318 -1230
rect 220 -1532 230 -1444
rect 300 -1532 310 -1444
rect 628 -1456 806 -1400
rect 1644 -1432 1680 -1360
rect 2402 -1424 2442 -1360
rect 2160 -1426 2442 -1424
rect 648 -1666 742 -1456
rect 1396 -1468 1680 -1432
rect 1780 -1514 1790 -1446
rect 1852 -1514 1862 -1446
rect 2138 -1452 2442 -1426
rect 3036 -1432 3080 -1354
rect 2402 -1526 2442 -1452
rect 2702 -1666 2770 -1440
rect 3036 -1466 3388 -1432
rect 3794 -1440 3834 -1358
rect 4664 -1362 4848 -1302
rect 4964 -1362 4974 -1344
rect 4664 -1424 4974 -1362
rect 4664 -1436 4848 -1424
rect 3606 -1520 3616 -1448
rect 3676 -1520 3686 -1448
rect 3794 -1472 4092 -1440
rect 4702 -1666 4796 -1436
rect 4964 -1452 4974 -1424
rect 5064 -1452 5074 -1344
rect 5404 -1558 5446 -1262
rect 5370 -1628 5380 -1558
rect 5484 -1628 5494 -1558
rect 7638 -1664 7674 -1256
rect 8442 -1664 8490 -1258
rect 5966 -1666 8276 -1664
rect 8324 -1666 8918 -1664
rect -372 -1898 8918 -1666
rect 5966 -1904 8918 -1898
<< via1 >>
rect -1008 -400 -882 -230
rect -1566 -688 -1440 -634
rect 1282 -222 1396 -52
rect 1016 -372 1170 -244
rect -1116 -804 -1002 -744
rect 358 -716 530 -604
rect 1278 -424 1386 -340
rect 1472 -728 1582 -614
rect 3814 -414 3896 -356
rect 4188 -166 4338 -78
rect 3810 -712 3886 -656
rect 4024 -432 4142 -340
rect 7442 -220 7516 -130
rect 8654 -246 8716 -176
rect 6366 -464 6508 -328
rect 7938 -332 8014 -268
rect 640 -1400 786 -1302
rect 5424 -716 5516 -646
rect 6588 -752 6668 -682
rect 7424 -750 7544 -678
rect 8244 -774 8338 -638
rect 8638 -1116 8814 -960
rect 230 -1532 300 -1444
rect 1790 -1514 1852 -1446
rect 3616 -1520 3676 -1448
rect 4974 -1452 5064 -1344
rect 5380 -1628 5484 -1558
<< metal2 >>
rect 1282 -52 1396 -42
rect -1008 -230 -882 -220
rect 4188 -78 4338 -68
rect 1396 -160 4188 -114
rect 4188 -176 4338 -166
rect 7442 -130 7516 -120
rect 1282 -232 1396 -222
rect 7434 -220 7442 -180
rect 7434 -230 7516 -220
rect 8654 -176 8716 -166
rect 1016 -244 1170 -234
rect -882 -342 1016 -268
rect 6366 -328 6508 -318
rect 1016 -382 1170 -372
rect 1278 -340 1386 -330
rect -1008 -410 -882 -400
rect 4024 -340 4142 -330
rect 3814 -356 3896 -346
rect 1386 -406 3814 -372
rect 3814 -424 3896 -414
rect 1278 -434 1386 -424
rect 4142 -420 6366 -358
rect 4024 -442 4142 -432
rect 6366 -474 6508 -464
rect 7434 -580 7482 -230
rect 8654 -256 8716 -246
rect 7938 -268 8014 -258
rect 7938 -342 8014 -332
rect 7434 -590 7520 -580
rect 8660 -588 8704 -256
rect 8102 -590 8704 -588
rect 358 -604 530 -594
rect -1566 -634 -1440 -624
rect -1566 -698 -1440 -688
rect -1540 -1718 -1458 -698
rect 1472 -614 1582 -604
rect 530 -696 1472 -654
rect 358 -726 530 -716
rect 7434 -624 8704 -590
rect 8102 -628 8704 -624
rect 5424 -646 5516 -636
rect 3810 -656 3886 -646
rect 3886 -704 5424 -666
rect 3810 -722 3886 -712
rect 8244 -638 8338 -628
rect 7462 -668 7504 -666
rect 5424 -726 5516 -716
rect 6588 -682 6668 -672
rect -1116 -744 -1002 -734
rect 1472 -738 1582 -728
rect 6588 -762 6668 -752
rect 7424 -678 7544 -668
rect 7932 -672 8018 -662
rect 7544 -736 7932 -694
rect 7424 -760 7544 -750
rect -1116 -814 -1002 -804
rect -1090 -1342 -1052 -814
rect 640 -1302 786 -1292
rect -1090 -1372 640 -1342
rect 640 -1410 786 -1400
rect 4974 -1344 5064 -1334
rect 230 -1444 300 -1434
rect 1790 -1446 1852 -1436
rect 300 -1514 1790 -1480
rect 300 -1516 1852 -1514
rect 1790 -1524 1852 -1516
rect 3616 -1448 3676 -1438
rect 6602 -1374 6646 -762
rect 7932 -768 8018 -758
rect 8244 -784 8338 -774
rect 8638 -960 8814 -950
rect 8638 -1126 8814 -1116
rect 5064 -1416 6646 -1374
rect 6602 -1420 6646 -1416
rect 4974 -1462 5064 -1452
rect 3616 -1530 3676 -1520
rect 230 -1542 300 -1532
rect 3634 -1574 3664 -1530
rect 5380 -1558 5484 -1548
rect 3634 -1614 5380 -1574
rect 5380 -1638 5484 -1628
rect 8686 -1708 8730 -1126
rect 6818 -1712 8732 -1708
rect 2372 -1718 8732 -1712
rect -1540 -1778 8732 -1718
rect -1540 -1794 7014 -1778
rect -1540 -1800 3102 -1794
<< via2 >>
rect 7938 -332 8014 -268
rect 7932 -758 8018 -672
<< metal3 >>
rect 7928 -268 8024 -263
rect 7928 -332 7938 -268
rect 8014 -332 8024 -268
rect 7928 -337 8024 -332
rect 7944 -667 8008 -337
rect 7922 -672 8028 -667
rect 7922 -758 7932 -672
rect 8018 -758 8028 -672
rect 7922 -763 8028 -758
use nmos4point5  nmos4point5_0
timestamp 1634617818
transform 1 0 880 0 1 -1490
box 0 0 690 286
use nmos12point5  nmos12point5_0
timestamp 1634616792
transform 1 0 1630 0 1 -1480
box 0 0 690 874
use nmos12point5  nmos12point5_1
timestamp 1634616792
transform 1 0 3148 0 1 -1486
box 0 0 690 874
use nmos8point5  nmos8point5_0
timestamp 1634616517
transform 1 0 2396 0 1 -1490
box 0 0 690 574
use nmos4point5  nmos4point5_1
timestamp 1634617818
transform 1 0 3898 0 1 -1490
box 0 0 690 286
use pmos8point5  pmos8point5_0
timestamp 1634618124
transform 1 0 40 0 1 24
box -40 -24 794 626
use pmos8point5  pmos8point5_1
timestamp 1634618124
transform 1 0 944 0 1 26
box -40 -24 794 626
use pmos8point5  pmos8point5_2
timestamp 1634618124
transform 1 0 1848 0 1 26
box -40 -24 794 626
use pmos8point5  pmos8point5_3
timestamp 1634618124
transform 1 0 2734 0 1 22
box -40 -24 794 626
use pmos8point5  pmos8point5_4
timestamp 1634618124
transform 1 0 3610 0 1 24
box -40 -24 794 626
use pmos8point5  pmos8point5_5
timestamp 1634618124
transform 1 0 4474 0 1 22
box -40 -24 794 626
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_3
timestamp 1632099954
transform 1 0 8272 0 1 -526
box -66 -43 354 897
use sky130_fd_pr__nfet_g5v0d10v5_R5T9XB  sky130_fd_pr__nfet_g5v0d10v5_R5T9XB_1
timestamp 1634629898
transform 1 0 8384 0 1 -1238
box -108 -126 108 126
use sky130_fd_pr__nfet_g5v0d10v5_R5T9XB  sky130_fd_pr__nfet_g5v0d10v5_R5T9XB_0
timestamp 1634629898
transform 1 0 7574 0 1 -1248
box -108 -126 108 126
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_2
timestamp 1632099954
transform 1 0 7452 0 1 -522
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_1
timestamp 1632099954
transform -1 0 -1076 0 1 -630
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_0
timestamp 1632099954
transform 1 0 6614 0 1 -540
box -66 -43 354 897
use pmos8point5  pmos8point5_7
timestamp 1634618124
transform 1 0 5060 0 1 -1352
box -40 -24 794 626
use pmos8point5  pmos8point5_6
timestamp 1634618124
transform 1 0 -296 0 1 -1378
box -40 -24 794 626
<< labels >>
flabel poly 3270 -518 3270 -518 0 FreeSans 800 0 0 0 vinp
flabel poly 3074 -1576 3074 -1576 0 FreeSans 800 0 0 0 vref
flabel poly 3016 820 3016 820 0 FreeSans 800 0 0 0 clk
flabel metal1 4010 -1810 4010 -1810 0 FreeSans 800 0 0 0 vssa
flabel metal1 2572 1128 2572 1128 0 FreeSans 800 0 0 0 vdda
flabel locali 6904 -200 6904 -200 0 FreeSans 800 0 0 0 vom
flabel locali -1380 -296 -1380 -296 0 FreeSans 800 0 0 0 vop
flabel metal1 7478 -894 7478 -894 0 FreeSans 800 0 0 0 vp
flabel metal1 8284 -1046 8284 -1046 0 FreeSans 800 0 0 0 vm
<< end >>
