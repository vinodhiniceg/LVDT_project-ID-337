magic
tech sky130A
magscale 1 2
timestamp 1634908693
<< nwell >>
rect -42 -38 1212 3002
<< poly >>
rect 116 2626 252 2702
rect 394 2622 530 2698
rect 644 2628 780 2704
rect 898 2622 1034 2698
rect 138 2334 274 2410
rect 402 2332 538 2408
rect 628 2334 764 2410
rect 894 2332 1030 2408
rect 114 2036 250 2112
rect 382 2038 518 2114
rect 650 2032 786 2108
rect 916 2042 1052 2118
rect 132 1746 268 1822
rect 384 1744 520 1820
rect 644 1738 780 1814
rect 898 1746 1034 1822
rect 120 1448 256 1524
rect 372 1442 508 1518
rect 638 1444 774 1520
rect 898 1452 1034 1528
rect 120 1154 256 1230
rect 406 1152 542 1228
rect 648 1150 784 1226
rect 894 1148 1030 1224
rect 118 860 254 936
rect 390 856 526 932
rect 638 860 774 936
rect 904 858 1040 934
rect 120 566 256 642
rect 374 556 510 632
rect 652 572 788 648
rect 924 568 1060 644
rect 122 272 258 348
rect 400 270 536 346
rect 638 272 774 348
rect 908 268 1044 344
<< metal1 >>
rect 546 2930 604 2932
rect 38 2918 1120 2930
rect 38 2884 1132 2918
rect 38 2820 96 2884
rect 34 2812 96 2820
rect 34 156 90 2812
rect 298 202 354 2824
rect 546 2820 604 2884
rect 546 2814 610 2820
rect 288 84 354 202
rect 554 156 610 2814
rect 810 196 866 2822
rect 1074 2800 1132 2884
rect 802 84 868 196
rect 1074 166 1130 2800
rect 288 40 876 84
rect 802 34 868 40
use sky130_fd_pr__pfet_g5v0d10v5_TMTL6D  sky130_fd_pr__pfet_g5v0d10v5_TMTL6D_0
timestamp 1634908693
transform 1 0 581 0 1 1485
box -611 -1489 611 1489
<< end >>
