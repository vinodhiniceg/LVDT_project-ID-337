magic
tech sky130A
magscale 1 2
timestamp 1634297993
<< pwell >>
rect -2844 -1243 2844 1243
<< mvnmos >>
rect -2616 47 -1616 1047
rect -1558 47 -558 1047
rect -500 47 500 1047
rect 558 47 1558 1047
rect 1616 47 2616 1047
rect -2616 -1047 -1616 -47
rect -1558 -1047 -558 -47
rect -500 -1047 500 -47
rect 558 -1047 1558 -47
rect 1616 -1047 2616 -47
<< mvndiff >>
rect -2674 693 -2616 1047
rect -2674 401 -2662 693
rect -2628 401 -2616 693
rect -2674 47 -2616 401
rect -1616 693 -1558 1047
rect -1616 401 -1604 693
rect -1570 401 -1558 693
rect -1616 47 -1558 401
rect -558 693 -500 1047
rect -558 401 -546 693
rect -512 401 -500 693
rect -558 47 -500 401
rect 500 693 558 1047
rect 500 401 512 693
rect 546 401 558 693
rect 500 47 558 401
rect 1558 693 1616 1047
rect 1558 401 1570 693
rect 1604 401 1616 693
rect 1558 47 1616 401
rect 2616 693 2674 1047
rect 2616 401 2628 693
rect 2662 401 2674 693
rect 2616 47 2674 401
rect -2674 -401 -2616 -47
rect -2674 -693 -2662 -401
rect -2628 -693 -2616 -401
rect -2674 -1047 -2616 -693
rect -1616 -401 -1558 -47
rect -1616 -693 -1604 -401
rect -1570 -693 -1558 -401
rect -1616 -1047 -1558 -693
rect -558 -401 -500 -47
rect -558 -693 -546 -401
rect -512 -693 -500 -401
rect -558 -1047 -500 -693
rect 500 -401 558 -47
rect 500 -693 512 -401
rect 546 -693 558 -401
rect 500 -1047 558 -693
rect 1558 -401 1616 -47
rect 1558 -693 1570 -401
rect 1604 -693 1616 -401
rect 1558 -1047 1616 -693
rect 2616 -401 2674 -47
rect 2616 -693 2628 -401
rect 2662 -693 2674 -401
rect 2616 -1047 2674 -693
<< mvndiffc >>
rect -2662 401 -2628 693
rect -1604 401 -1570 693
rect -546 401 -512 693
rect 512 401 546 693
rect 1570 401 1604 693
rect 2628 401 2662 693
rect -2662 -693 -2628 -401
rect -1604 -693 -1570 -401
rect -546 -693 -512 -401
rect 512 -693 546 -401
rect 1570 -693 1604 -401
rect 2628 -693 2662 -401
<< mvpsubdiff >>
rect -2808 1149 2808 1207
rect -2808 550 -2750 1149
rect -2808 -550 -2796 550
rect -2762 -550 -2750 550
rect 2750 550 2808 1149
rect -2808 -1149 -2750 -550
rect 2750 -550 2762 550
rect 2796 -550 2808 550
rect 2750 -1149 2808 -550
rect -2808 -1207 2808 -1149
<< mvpsubdiffcont >>
rect -2796 -550 -2762 550
rect 2762 -550 2796 550
<< poly >>
rect -2616 1047 -1616 1073
rect -1558 1047 -558 1073
rect -500 1047 500 1073
rect 558 1047 1558 1073
rect 1616 1047 2616 1073
rect -2616 21 -1616 47
rect -1558 21 -558 47
rect -500 21 500 47
rect 558 21 1558 47
rect 1616 21 2616 47
rect -2616 -47 -1616 -21
rect -1558 -47 -558 -21
rect -500 -47 500 -21
rect 558 -47 1558 -21
rect 1616 -47 2616 -21
rect -2616 -1073 -1616 -1047
rect -1558 -1073 -558 -1047
rect -500 -1073 500 -1047
rect 558 -1073 1558 -1047
rect 1616 -1073 2616 -1047
<< locali >>
rect -2662 693 -2628 709
rect -2796 550 -2762 566
rect -2662 385 -2628 401
rect -1604 693 -1570 709
rect -1604 385 -1570 401
rect -546 693 -512 709
rect -546 385 -512 401
rect 512 693 546 709
rect 512 385 546 401
rect 1570 693 1604 709
rect 1570 385 1604 401
rect 2628 693 2662 709
rect 2628 385 2662 401
rect 2762 550 2796 566
rect -2796 -566 -2762 -550
rect -2662 -401 -2628 -385
rect -2662 -709 -2628 -693
rect -1604 -401 -1570 -385
rect -1604 -709 -1570 -693
rect -546 -401 -512 -385
rect -546 -709 -512 -693
rect 512 -401 546 -385
rect 512 -709 546 -693
rect 1570 -401 1604 -385
rect 1570 -709 1604 -693
rect 2628 -401 2662 -385
rect 2762 -566 2796 -550
rect 2628 -709 2662 -693
<< viali >>
rect -2662 401 -2628 693
rect -1604 401 -1570 693
rect -546 401 -512 693
rect 512 401 546 693
rect 1570 401 1604 693
rect 2628 401 2662 693
rect -2662 -693 -2628 -401
rect -1604 -693 -1570 -401
rect -546 -693 -512 -401
rect 512 -693 546 -401
rect 1570 -693 1604 -401
rect 2628 -693 2662 -401
<< metal1 >>
rect -2668 693 -2622 705
rect -2668 401 -2662 693
rect -2628 401 -2622 693
rect -2668 389 -2622 401
rect -1610 693 -1564 705
rect -1610 401 -1604 693
rect -1570 401 -1564 693
rect -1610 389 -1564 401
rect -552 693 -506 705
rect -552 401 -546 693
rect -512 401 -506 693
rect -552 389 -506 401
rect 506 693 552 705
rect 506 401 512 693
rect 546 401 552 693
rect 506 389 552 401
rect 1564 693 1610 705
rect 1564 401 1570 693
rect 1604 401 1610 693
rect 1564 389 1610 401
rect 2622 693 2668 705
rect 2622 401 2628 693
rect 2662 401 2668 693
rect 2622 389 2668 401
rect -2668 -401 -2622 -389
rect -2668 -693 -2662 -401
rect -2628 -693 -2622 -401
rect -2668 -705 -2622 -693
rect -1610 -401 -1564 -389
rect -1610 -693 -1604 -401
rect -1570 -693 -1564 -401
rect -1610 -705 -1564 -693
rect -552 -401 -506 -389
rect -552 -693 -546 -401
rect -512 -693 -506 -401
rect -552 -705 -506 -693
rect 506 -401 552 -389
rect 506 -693 512 -401
rect 546 -693 552 -401
rect 506 -705 552 -693
rect 1564 -401 1610 -389
rect 1564 -693 1570 -401
rect 1604 -693 1610 -401
rect 1564 -705 1610 -693
rect 2622 -401 2668 -389
rect 2622 -693 2628 -401
rect 2662 -693 2668 -401
rect 2622 -705 2668 -693
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string FIXED_BBOX -2779 -1178 2779 1178
string parameters w 5 l 5 m 2 nf 5 diffcov 30 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 50 rlcov 50 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 30 viadrn 30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
