magic
tech sky130A
magscale 1 2
timestamp 1634908262
<< mvnmos >>
rect -229 2252 -29 2452
rect 29 2252 229 2452
rect -229 1958 -29 2158
rect 29 1958 229 2158
rect -229 1664 -29 1864
rect 29 1664 229 1864
rect -229 1370 -29 1570
rect 29 1370 229 1570
rect -229 1076 -29 1276
rect 29 1076 229 1276
rect -229 782 -29 982
rect 29 782 229 982
rect -229 488 -29 688
rect 29 488 229 688
rect -229 194 -29 394
rect 29 194 229 394
rect -229 -100 -29 100
rect 29 -100 229 100
rect -229 -394 -29 -194
rect 29 -394 229 -194
rect -229 -688 -29 -488
rect 29 -688 229 -488
rect -229 -982 -29 -782
rect 29 -982 229 -782
rect -229 -1276 -29 -1076
rect 29 -1276 229 -1076
rect -229 -1570 -29 -1370
rect 29 -1570 229 -1370
rect -229 -1864 -29 -1664
rect 29 -1864 229 -1664
rect -229 -2158 -29 -1958
rect 29 -2158 229 -1958
rect -229 -2452 -29 -2252
rect 29 -2452 229 -2252
<< mvndiff >>
rect -287 2378 -229 2452
rect -287 2326 -275 2378
rect -241 2326 -229 2378
rect -287 2252 -229 2326
rect -29 2378 29 2452
rect -29 2326 -17 2378
rect 17 2326 29 2378
rect -29 2252 29 2326
rect 229 2378 287 2452
rect 229 2326 241 2378
rect 275 2326 287 2378
rect 229 2252 287 2326
rect -287 2084 -229 2158
rect -287 2032 -275 2084
rect -241 2032 -229 2084
rect -287 1958 -229 2032
rect -29 2084 29 2158
rect -29 2032 -17 2084
rect 17 2032 29 2084
rect -29 1958 29 2032
rect 229 2084 287 2158
rect 229 2032 241 2084
rect 275 2032 287 2084
rect 229 1958 287 2032
rect -287 1790 -229 1864
rect -287 1738 -275 1790
rect -241 1738 -229 1790
rect -287 1664 -229 1738
rect -29 1790 29 1864
rect -29 1738 -17 1790
rect 17 1738 29 1790
rect -29 1664 29 1738
rect 229 1790 287 1864
rect 229 1738 241 1790
rect 275 1738 287 1790
rect 229 1664 287 1738
rect -287 1496 -229 1570
rect -287 1444 -275 1496
rect -241 1444 -229 1496
rect -287 1370 -229 1444
rect -29 1496 29 1570
rect -29 1444 -17 1496
rect 17 1444 29 1496
rect -29 1370 29 1444
rect 229 1496 287 1570
rect 229 1444 241 1496
rect 275 1444 287 1496
rect 229 1370 287 1444
rect -287 1202 -229 1276
rect -287 1150 -275 1202
rect -241 1150 -229 1202
rect -287 1076 -229 1150
rect -29 1202 29 1276
rect -29 1150 -17 1202
rect 17 1150 29 1202
rect -29 1076 29 1150
rect 229 1202 287 1276
rect 229 1150 241 1202
rect 275 1150 287 1202
rect 229 1076 287 1150
rect -287 908 -229 982
rect -287 856 -275 908
rect -241 856 -229 908
rect -287 782 -229 856
rect -29 908 29 982
rect -29 856 -17 908
rect 17 856 29 908
rect -29 782 29 856
rect 229 908 287 982
rect 229 856 241 908
rect 275 856 287 908
rect 229 782 287 856
rect -287 614 -229 688
rect -287 562 -275 614
rect -241 562 -229 614
rect -287 488 -229 562
rect -29 614 29 688
rect -29 562 -17 614
rect 17 562 29 614
rect -29 488 29 562
rect 229 614 287 688
rect 229 562 241 614
rect 275 562 287 614
rect 229 488 287 562
rect -287 320 -229 394
rect -287 268 -275 320
rect -241 268 -229 320
rect -287 194 -229 268
rect -29 320 29 394
rect -29 268 -17 320
rect 17 268 29 320
rect -29 194 29 268
rect 229 320 287 394
rect 229 268 241 320
rect 275 268 287 320
rect 229 194 287 268
rect -287 26 -229 100
rect -287 -26 -275 26
rect -241 -26 -229 26
rect -287 -100 -229 -26
rect -29 26 29 100
rect -29 -26 -17 26
rect 17 -26 29 26
rect -29 -100 29 -26
rect 229 26 287 100
rect 229 -26 241 26
rect 275 -26 287 26
rect 229 -100 287 -26
rect -287 -268 -229 -194
rect -287 -320 -275 -268
rect -241 -320 -229 -268
rect -287 -394 -229 -320
rect -29 -268 29 -194
rect -29 -320 -17 -268
rect 17 -320 29 -268
rect -29 -394 29 -320
rect 229 -268 287 -194
rect 229 -320 241 -268
rect 275 -320 287 -268
rect 229 -394 287 -320
rect -287 -562 -229 -488
rect -287 -614 -275 -562
rect -241 -614 -229 -562
rect -287 -688 -229 -614
rect -29 -562 29 -488
rect -29 -614 -17 -562
rect 17 -614 29 -562
rect -29 -688 29 -614
rect 229 -562 287 -488
rect 229 -614 241 -562
rect 275 -614 287 -562
rect 229 -688 287 -614
rect -287 -856 -229 -782
rect -287 -908 -275 -856
rect -241 -908 -229 -856
rect -287 -982 -229 -908
rect -29 -856 29 -782
rect -29 -908 -17 -856
rect 17 -908 29 -856
rect -29 -982 29 -908
rect 229 -856 287 -782
rect 229 -908 241 -856
rect 275 -908 287 -856
rect 229 -982 287 -908
rect -287 -1150 -229 -1076
rect -287 -1202 -275 -1150
rect -241 -1202 -229 -1150
rect -287 -1276 -229 -1202
rect -29 -1150 29 -1076
rect -29 -1202 -17 -1150
rect 17 -1202 29 -1150
rect -29 -1276 29 -1202
rect 229 -1150 287 -1076
rect 229 -1202 241 -1150
rect 275 -1202 287 -1150
rect 229 -1276 287 -1202
rect -287 -1444 -229 -1370
rect -287 -1496 -275 -1444
rect -241 -1496 -229 -1444
rect -287 -1570 -229 -1496
rect -29 -1444 29 -1370
rect -29 -1496 -17 -1444
rect 17 -1496 29 -1444
rect -29 -1570 29 -1496
rect 229 -1444 287 -1370
rect 229 -1496 241 -1444
rect 275 -1496 287 -1444
rect 229 -1570 287 -1496
rect -287 -1738 -229 -1664
rect -287 -1790 -275 -1738
rect -241 -1790 -229 -1738
rect -287 -1864 -229 -1790
rect -29 -1738 29 -1664
rect -29 -1790 -17 -1738
rect 17 -1790 29 -1738
rect -29 -1864 29 -1790
rect 229 -1738 287 -1664
rect 229 -1790 241 -1738
rect 275 -1790 287 -1738
rect 229 -1864 287 -1790
rect -287 -2032 -229 -1958
rect -287 -2084 -275 -2032
rect -241 -2084 -229 -2032
rect -287 -2158 -229 -2084
rect -29 -2032 29 -1958
rect -29 -2084 -17 -2032
rect 17 -2084 29 -2032
rect -29 -2158 29 -2084
rect 229 -2032 287 -1958
rect 229 -2084 241 -2032
rect 275 -2084 287 -2032
rect 229 -2158 287 -2084
rect -287 -2326 -229 -2252
rect -287 -2378 -275 -2326
rect -241 -2378 -229 -2326
rect -287 -2452 -229 -2378
rect -29 -2326 29 -2252
rect -29 -2378 -17 -2326
rect 17 -2378 29 -2326
rect -29 -2452 29 -2378
rect 229 -2326 287 -2252
rect 229 -2378 241 -2326
rect 275 -2378 287 -2326
rect 229 -2452 287 -2378
<< mvndiffc >>
rect -275 2326 -241 2378
rect -17 2326 17 2378
rect 241 2326 275 2378
rect -275 2032 -241 2084
rect -17 2032 17 2084
rect 241 2032 275 2084
rect -275 1738 -241 1790
rect -17 1738 17 1790
rect 241 1738 275 1790
rect -275 1444 -241 1496
rect -17 1444 17 1496
rect 241 1444 275 1496
rect -275 1150 -241 1202
rect -17 1150 17 1202
rect 241 1150 275 1202
rect -275 856 -241 908
rect -17 856 17 908
rect 241 856 275 908
rect -275 562 -241 614
rect -17 562 17 614
rect 241 562 275 614
rect -275 268 -241 320
rect -17 268 17 320
rect 241 268 275 320
rect -275 -26 -241 26
rect -17 -26 17 26
rect 241 -26 275 26
rect -275 -320 -241 -268
rect -17 -320 17 -268
rect 241 -320 275 -268
rect -275 -614 -241 -562
rect -17 -614 17 -562
rect 241 -614 275 -562
rect -275 -908 -241 -856
rect -17 -908 17 -856
rect 241 -908 275 -856
rect -275 -1202 -241 -1150
rect -17 -1202 17 -1150
rect 241 -1202 275 -1150
rect -275 -1496 -241 -1444
rect -17 -1496 17 -1444
rect 241 -1496 275 -1444
rect -275 -1790 -241 -1738
rect -17 -1790 17 -1738
rect 241 -1790 275 -1738
rect -275 -2084 -241 -2032
rect -17 -2084 17 -2032
rect 241 -2084 275 -2032
rect -275 -2378 -241 -2326
rect -17 -2378 17 -2326
rect 241 -2378 275 -2326
<< poly >>
rect -229 2452 -29 2478
rect 29 2452 229 2478
rect -229 2226 -29 2252
rect 29 2226 229 2252
rect -229 2158 -29 2184
rect 29 2158 229 2184
rect -229 1932 -29 1958
rect 29 1932 229 1958
rect -229 1864 -29 1890
rect 29 1864 229 1890
rect -229 1638 -29 1664
rect 29 1638 229 1664
rect -229 1570 -29 1596
rect 29 1570 229 1596
rect -229 1344 -29 1370
rect 29 1344 229 1370
rect -229 1276 -29 1302
rect 29 1276 229 1302
rect -229 1050 -29 1076
rect 29 1050 229 1076
rect -229 982 -29 1008
rect 29 982 229 1008
rect -229 756 -29 782
rect 29 756 229 782
rect -229 688 -29 714
rect 29 688 229 714
rect -229 462 -29 488
rect 29 462 229 488
rect -229 394 -29 420
rect 29 394 229 420
rect -229 168 -29 194
rect 29 168 229 194
rect -229 100 -29 126
rect 29 100 229 126
rect -229 -126 -29 -100
rect 29 -126 229 -100
rect -229 -194 -29 -168
rect 29 -194 229 -168
rect -229 -420 -29 -394
rect 29 -420 229 -394
rect -229 -488 -29 -462
rect 29 -488 229 -462
rect -229 -714 -29 -688
rect 29 -714 229 -688
rect -229 -782 -29 -756
rect 29 -782 229 -756
rect -229 -1008 -29 -982
rect 29 -1008 229 -982
rect -229 -1076 -29 -1050
rect 29 -1076 229 -1050
rect -229 -1302 -29 -1276
rect 29 -1302 229 -1276
rect -229 -1370 -29 -1344
rect 29 -1370 229 -1344
rect -229 -1596 -29 -1570
rect 29 -1596 229 -1570
rect -229 -1664 -29 -1638
rect 29 -1664 229 -1638
rect -229 -1890 -29 -1864
rect 29 -1890 229 -1864
rect -229 -1958 -29 -1932
rect 29 -1958 229 -1932
rect -229 -2184 -29 -2158
rect 29 -2184 229 -2158
rect -229 -2252 -29 -2226
rect 29 -2252 229 -2226
rect -229 -2478 -29 -2452
rect 29 -2478 229 -2452
<< locali >>
rect -275 2378 -241 2394
rect -275 2310 -241 2326
rect -17 2378 17 2394
rect -17 2310 17 2326
rect 241 2378 275 2394
rect 241 2310 275 2326
rect -275 2084 -241 2100
rect -275 2016 -241 2032
rect -17 2084 17 2100
rect -17 2016 17 2032
rect 241 2084 275 2100
rect 241 2016 275 2032
rect -275 1790 -241 1806
rect -275 1722 -241 1738
rect -17 1790 17 1806
rect -17 1722 17 1738
rect 241 1790 275 1806
rect 241 1722 275 1738
rect -275 1496 -241 1512
rect -275 1428 -241 1444
rect -17 1496 17 1512
rect -17 1428 17 1444
rect 241 1496 275 1512
rect 241 1428 275 1444
rect -275 1202 -241 1218
rect -275 1134 -241 1150
rect -17 1202 17 1218
rect -17 1134 17 1150
rect 241 1202 275 1218
rect 241 1134 275 1150
rect -275 908 -241 924
rect -275 840 -241 856
rect -17 908 17 924
rect -17 840 17 856
rect 241 908 275 924
rect 241 840 275 856
rect -275 614 -241 630
rect -275 546 -241 562
rect -17 614 17 630
rect -17 546 17 562
rect 241 614 275 630
rect 241 546 275 562
rect -275 320 -241 336
rect -275 252 -241 268
rect -17 320 17 336
rect -17 252 17 268
rect 241 320 275 336
rect 241 252 275 268
rect -275 26 -241 42
rect -275 -42 -241 -26
rect -17 26 17 42
rect -17 -42 17 -26
rect 241 26 275 42
rect 241 -42 275 -26
rect -275 -268 -241 -252
rect -275 -336 -241 -320
rect -17 -268 17 -252
rect -17 -336 17 -320
rect 241 -268 275 -252
rect 241 -336 275 -320
rect -275 -562 -241 -546
rect -275 -630 -241 -614
rect -17 -562 17 -546
rect -17 -630 17 -614
rect 241 -562 275 -546
rect 241 -630 275 -614
rect -275 -856 -241 -840
rect -275 -924 -241 -908
rect -17 -856 17 -840
rect -17 -924 17 -908
rect 241 -856 275 -840
rect 241 -924 275 -908
rect -275 -1150 -241 -1134
rect -275 -1218 -241 -1202
rect -17 -1150 17 -1134
rect -17 -1218 17 -1202
rect 241 -1150 275 -1134
rect 241 -1218 275 -1202
rect -275 -1444 -241 -1428
rect -275 -1512 -241 -1496
rect -17 -1444 17 -1428
rect -17 -1512 17 -1496
rect 241 -1444 275 -1428
rect 241 -1512 275 -1496
rect -275 -1738 -241 -1722
rect -275 -1806 -241 -1790
rect -17 -1738 17 -1722
rect -17 -1806 17 -1790
rect 241 -1738 275 -1722
rect 241 -1806 275 -1790
rect -275 -2032 -241 -2016
rect -275 -2100 -241 -2084
rect -17 -2032 17 -2016
rect -17 -2100 17 -2084
rect 241 -2032 275 -2016
rect 241 -2100 275 -2084
rect -275 -2326 -241 -2310
rect -275 -2394 -241 -2378
rect -17 -2326 17 -2310
rect -17 -2394 17 -2378
rect 241 -2326 275 -2310
rect 241 -2394 275 -2378
<< viali >>
rect -275 2326 -241 2378
rect -17 2326 17 2378
rect 241 2326 275 2378
rect -275 2032 -241 2084
rect -17 2032 17 2084
rect 241 2032 275 2084
rect -275 1738 -241 1790
rect -17 1738 17 1790
rect 241 1738 275 1790
rect -275 1444 -241 1496
rect -17 1444 17 1496
rect 241 1444 275 1496
rect -275 1150 -241 1202
rect -17 1150 17 1202
rect 241 1150 275 1202
rect -275 856 -241 908
rect -17 856 17 908
rect 241 856 275 908
rect -275 562 -241 614
rect -17 562 17 614
rect 241 562 275 614
rect -275 268 -241 320
rect -17 268 17 320
rect 241 268 275 320
rect -275 -26 -241 26
rect -17 -26 17 26
rect 241 -26 275 26
rect -275 -320 -241 -268
rect -17 -320 17 -268
rect 241 -320 275 -268
rect -275 -614 -241 -562
rect -17 -614 17 -562
rect 241 -614 275 -562
rect -275 -908 -241 -856
rect -17 -908 17 -856
rect 241 -908 275 -856
rect -275 -1202 -241 -1150
rect -17 -1202 17 -1150
rect 241 -1202 275 -1150
rect -275 -1496 -241 -1444
rect -17 -1496 17 -1444
rect 241 -1496 275 -1444
rect -275 -1790 -241 -1738
rect -17 -1790 17 -1738
rect 241 -1790 275 -1738
rect -275 -2084 -241 -2032
rect -17 -2084 17 -2032
rect 241 -2084 275 -2032
rect -275 -2378 -241 -2326
rect -17 -2378 17 -2326
rect 241 -2378 275 -2326
<< metal1 >>
rect -281 2378 -235 2390
rect -281 2326 -275 2378
rect -241 2326 -235 2378
rect -281 2314 -235 2326
rect -23 2378 23 2390
rect -23 2326 -17 2378
rect 17 2326 23 2378
rect -23 2314 23 2326
rect 235 2378 281 2390
rect 235 2326 241 2378
rect 275 2326 281 2378
rect 235 2314 281 2326
rect -281 2084 -235 2096
rect -281 2032 -275 2084
rect -241 2032 -235 2084
rect -281 2020 -235 2032
rect -23 2084 23 2096
rect -23 2032 -17 2084
rect 17 2032 23 2084
rect -23 2020 23 2032
rect 235 2084 281 2096
rect 235 2032 241 2084
rect 275 2032 281 2084
rect 235 2020 281 2032
rect -281 1790 -235 1802
rect -281 1738 -275 1790
rect -241 1738 -235 1790
rect -281 1726 -235 1738
rect -23 1790 23 1802
rect -23 1738 -17 1790
rect 17 1738 23 1790
rect -23 1726 23 1738
rect 235 1790 281 1802
rect 235 1738 241 1790
rect 275 1738 281 1790
rect 235 1726 281 1738
rect -281 1496 -235 1508
rect -281 1444 -275 1496
rect -241 1444 -235 1496
rect -281 1432 -235 1444
rect -23 1496 23 1508
rect -23 1444 -17 1496
rect 17 1444 23 1496
rect -23 1432 23 1444
rect 235 1496 281 1508
rect 235 1444 241 1496
rect 275 1444 281 1496
rect 235 1432 281 1444
rect -281 1202 -235 1214
rect -281 1150 -275 1202
rect -241 1150 -235 1202
rect -281 1138 -235 1150
rect -23 1202 23 1214
rect -23 1150 -17 1202
rect 17 1150 23 1202
rect -23 1138 23 1150
rect 235 1202 281 1214
rect 235 1150 241 1202
rect 275 1150 281 1202
rect 235 1138 281 1150
rect -281 908 -235 920
rect -281 856 -275 908
rect -241 856 -235 908
rect -281 844 -235 856
rect -23 908 23 920
rect -23 856 -17 908
rect 17 856 23 908
rect -23 844 23 856
rect 235 908 281 920
rect 235 856 241 908
rect 275 856 281 908
rect 235 844 281 856
rect -281 614 -235 626
rect -281 562 -275 614
rect -241 562 -235 614
rect -281 550 -235 562
rect -23 614 23 626
rect -23 562 -17 614
rect 17 562 23 614
rect -23 550 23 562
rect 235 614 281 626
rect 235 562 241 614
rect 275 562 281 614
rect 235 550 281 562
rect -281 320 -235 332
rect -281 268 -275 320
rect -241 268 -235 320
rect -281 256 -235 268
rect -23 320 23 332
rect -23 268 -17 320
rect 17 268 23 320
rect -23 256 23 268
rect 235 320 281 332
rect 235 268 241 320
rect 275 268 281 320
rect 235 256 281 268
rect -281 26 -235 38
rect -281 -26 -275 26
rect -241 -26 -235 26
rect -281 -38 -235 -26
rect -23 26 23 38
rect -23 -26 -17 26
rect 17 -26 23 26
rect -23 -38 23 -26
rect 235 26 281 38
rect 235 -26 241 26
rect 275 -26 281 26
rect 235 -38 281 -26
rect -281 -268 -235 -256
rect -281 -320 -275 -268
rect -241 -320 -235 -268
rect -281 -332 -235 -320
rect -23 -268 23 -256
rect -23 -320 -17 -268
rect 17 -320 23 -268
rect -23 -332 23 -320
rect 235 -268 281 -256
rect 235 -320 241 -268
rect 275 -320 281 -268
rect 235 -332 281 -320
rect -281 -562 -235 -550
rect -281 -614 -275 -562
rect -241 -614 -235 -562
rect -281 -626 -235 -614
rect -23 -562 23 -550
rect -23 -614 -17 -562
rect 17 -614 23 -562
rect -23 -626 23 -614
rect 235 -562 281 -550
rect 235 -614 241 -562
rect 275 -614 281 -562
rect 235 -626 281 -614
rect -281 -856 -235 -844
rect -281 -908 -275 -856
rect -241 -908 -235 -856
rect -281 -920 -235 -908
rect -23 -856 23 -844
rect -23 -908 -17 -856
rect 17 -908 23 -856
rect -23 -920 23 -908
rect 235 -856 281 -844
rect 235 -908 241 -856
rect 275 -908 281 -856
rect 235 -920 281 -908
rect -281 -1150 -235 -1138
rect -281 -1202 -275 -1150
rect -241 -1202 -235 -1150
rect -281 -1214 -235 -1202
rect -23 -1150 23 -1138
rect -23 -1202 -17 -1150
rect 17 -1202 23 -1150
rect -23 -1214 23 -1202
rect 235 -1150 281 -1138
rect 235 -1202 241 -1150
rect 275 -1202 281 -1150
rect 235 -1214 281 -1202
rect -281 -1444 -235 -1432
rect -281 -1496 -275 -1444
rect -241 -1496 -235 -1444
rect -281 -1508 -235 -1496
rect -23 -1444 23 -1432
rect -23 -1496 -17 -1444
rect 17 -1496 23 -1444
rect -23 -1508 23 -1496
rect 235 -1444 281 -1432
rect 235 -1496 241 -1444
rect 275 -1496 281 -1444
rect 235 -1508 281 -1496
rect -281 -1738 -235 -1726
rect -281 -1790 -275 -1738
rect -241 -1790 -235 -1738
rect -281 -1802 -235 -1790
rect -23 -1738 23 -1726
rect -23 -1790 -17 -1738
rect 17 -1790 23 -1738
rect -23 -1802 23 -1790
rect 235 -1738 281 -1726
rect 235 -1790 241 -1738
rect 275 -1790 281 -1738
rect 235 -1802 281 -1790
rect -281 -2032 -235 -2020
rect -281 -2084 -275 -2032
rect -241 -2084 -235 -2032
rect -281 -2096 -235 -2084
rect -23 -2032 23 -2020
rect -23 -2084 -17 -2032
rect 17 -2084 23 -2032
rect -23 -2096 23 -2084
rect 235 -2032 281 -2020
rect 235 -2084 241 -2032
rect 275 -2084 281 -2032
rect 235 -2096 281 -2084
rect -281 -2326 -235 -2314
rect -281 -2378 -275 -2326
rect -241 -2378 -235 -2326
rect -281 -2390 -235 -2378
rect -23 -2326 23 -2314
rect -23 -2378 -17 -2326
rect 17 -2378 23 -2326
rect -23 -2390 23 -2378
rect 235 -2326 281 -2314
rect 235 -2378 241 -2326
rect 275 -2378 281 -2326
rect 235 -2390 281 -2378
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string parameters w 1 l 1 m 17 nf 2 diffcov 30 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 30 viadrn 30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
