magic
tech sky130A
magscale 1 2
timestamp 1634225045
<< mvpsubdiff >>
rect -524 3768 -180 3870
rect -524 420 -446 3768
rect -218 420 -180 3768
rect -524 318 -180 420
<< mvpsubdiffcont >>
rect -446 420 -218 3768
<< poly >>
rect 362 4120 2488 4202
rect 216 3414 548 3484
rect 862 3412 1194 3482
rect 1574 3414 1906 3484
rect 2164 3414 2496 3484
rect 180 2718 512 2788
rect 886 2720 1218 2790
rect 1548 2720 1880 2790
rect 2126 2720 2458 2790
rect 184 2026 516 2096
rect 888 2028 1220 2098
rect 1526 2028 1858 2098
rect 2170 2028 2502 2098
rect 178 1332 510 1402
rect 858 1330 1190 1400
rect 1542 1330 1874 1400
rect 2176 1334 2508 1404
rect 172 638 504 708
rect 888 636 1220 706
rect 1518 638 1850 708
rect 2190 638 2522 708
<< locali >>
rect -70 4042 84 4186
rect 1318 4042 1380 4052
rect 2618 4042 2680 4072
rect -70 3988 2702 4042
rect -70 3948 84 3988
rect -524 3768 -180 3870
rect -14 3840 48 3948
rect -14 3794 52 3840
rect -524 420 -446 3768
rect -218 420 -180 3768
rect -524 318 -180 420
rect 2 312 48 3794
rect 662 328 708 3820
rect 1318 3818 1380 3988
rect 2618 3874 2680 3988
rect 1320 328 1366 3818
rect 1980 340 2026 3832
rect 2618 3802 2686 3874
rect 2640 344 2686 3802
rect 650 120 712 292
rect 1962 120 2024 284
rect 650 58 2034 120
rect 662 54 2034 58
rect 1038 -112 1112 54
rect 1962 50 2024 54
<< viali >>
rect -398 482 -250 3704
<< metal1 >>
rect -524 3704 -180 3870
rect -524 482 -398 3704
rect -250 482 -180 3704
rect -524 318 -180 482
use sky130_fd_pr__nfet_g5v0d10v5_GZ7LRN  sky130_fd_pr__nfet_g5v0d10v5_GZ7LRN_0
timestamp 1634224850
transform 1 0 1345 0 1 2061
box -1345 -2061 1345 2061
<< labels >>
flabel locali -34 4104 -34 4104 0 FreeSans 1600 0 0 0 d
flabel poly 1456 4172 1456 4172 0 FreeSans 1600 0 0 0 g
flabel locali 1074 -62 1074 -62 0 FreeSans 1600 0 0 0 s
flabel metal1 -428 3718 -428 3718 0 FreeSans 1600 0 0 0 sub
<< end >>
