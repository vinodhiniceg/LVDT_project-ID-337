magic
tech sky130A
magscale 1 2
timestamp 1634049374
<< pwell >>
rect -1010 -162 4674 10632
<< mvpsubdiff >>
rect -938 9182 -290 9430
rect -938 1494 -816 9182
rect -474 1494 -290 9182
rect -938 1184 -290 1494
<< mvpsubdiffcont >>
rect -816 1494 -474 9182
<< poly >>
rect 1054 10418 2830 10564
rect 734 8320 1560 8392
rect 2566 8314 3392 8386
rect 802 6222 1628 6294
rect 2644 6226 3470 6298
rect 534 4130 1360 4202
rect 2550 4126 3376 4198
rect 662 2040 1488 2112
rect 2658 2040 3484 2112
<< locali >>
rect -938 9182 -290 9430
rect -938 1494 -816 9182
rect -474 1494 -290 9182
rect -938 1184 -290 1494
rect -14 1390 52 9622
rect 2020 9546 2160 10122
rect -38 452 56 1390
rect 2050 1192 2116 9546
rect 4108 1342 4174 9720
rect 4102 452 4196 1342
rect -38 352 4196 452
rect -16 304 4196 352
<< viali >>
rect -784 1880 -522 8936
<< metal1 >>
rect -938 8936 -290 9430
rect -938 1880 -784 8936
rect -522 1880 -290 8936
rect -938 1184 -290 1880
use sky130_fd_pr__nfet_g5v0d10v5_C8B57Z  sky130_fd_pr__nfet_g5v0d10v5_C8B57Z_0 ~/layout test
timestamp 1634045799
transform 1 0 2087 0 1 5214
box -2087 -5214 2087 5214
<< end >>
