magic
tech sky130A
magscale 1 2
timestamp 1634121920
<< nwell >>
rect -464 -250 5454 2302
rect -430 -274 5454 -250
rect -202 -284 5454 -274
<< mvnsubdiff >>
rect -334 1852 -140 1894
rect -334 338 -310 1852
rect -168 338 -140 1852
rect -334 282 -140 338
<< mvnsubdiffcont >>
rect -310 338 -168 1852
<< poly >>
rect 468 2072 5264 2102
rect 184 1366 552 1436
rect 870 1362 1238 1432
rect 1482 1372 1850 1442
rect 2176 1372 2544 1442
rect 2844 1370 3212 1440
rect 3546 1364 3914 1434
rect 4200 1364 4568 1434
rect 4840 1360 5194 1442
rect 190 674 558 744
rect 866 674 1234 744
rect 1528 672 1896 742
rect 2174 678 2542 748
rect 2866 674 3234 744
rect 3532 676 3900 746
rect 4204 670 4572 740
rect 4828 672 5182 754
<< locali >>
rect 18 2016 102 2040
rect 18 2012 4714 2016
rect 5298 2012 5368 2016
rect 18 1948 5368 2012
rect -344 1852 -140 1914
rect -344 338 -310 1852
rect -168 338 -140 1852
rect 18 1746 102 1948
rect -344 282 -140 338
rect 30 246 94 1746
rect 694 404 746 1812
rect 1356 1728 1410 1948
rect 672 158 794 404
rect 1356 294 1408 1728
rect 2016 390 2068 1816
rect 2668 1740 2722 1948
rect 1994 158 2116 390
rect 2670 308 2722 1740
rect 3330 380 3382 1826
rect 3986 1730 4040 1948
rect 4672 1938 5368 1948
rect 3308 158 3430 380
rect 3988 332 4040 1730
rect 4644 370 4696 1874
rect 5298 1794 5368 1938
rect 4596 158 4718 370
rect 5304 368 5356 1794
rect 672 84 4718 158
rect 696 66 4718 84
rect 3308 60 3430 66
rect 4596 50 4718 66
<< viali >>
rect -286 396 -216 1800
<< metal1 >>
rect -344 1800 -140 1914
rect -344 396 -286 1800
rect -216 396 -140 1800
rect -344 282 -140 396
use sky130_fd_pr__pfet_g5v0d10v5_2CSA4Z  sky130_fd_pr__pfet_g5v0d10v5_2CSA4Z_0 ~/layout test
timestamp 1634118957
transform 1 0 2697 0 1 1056
box -2727 -1060 2727 1060
<< end >>
