magic
tech sky130A
magscale 1 2
timestamp 1634049309
<< pwell >>
rect -1164 -238 4674 8552
<< mvpsubdiff >>
rect -1042 7360 -556 7518
rect -1042 1414 -1002 7360
rect -608 1414 -556 7360
rect -1042 1238 -556 1414
<< mvpsubdiffcont >>
rect -1002 1414 -608 7360
<< poly >>
rect 1382 8330 3204 8372
rect 476 6226 1552 6300
rect 2540 6218 3616 6292
rect 526 4134 1602 4208
rect 2620 4132 3696 4206
rect 480 2036 1556 2110
rect 2550 2032 3626 2106
<< locali >>
rect 2052 7868 2112 8156
rect -1042 7360 -556 7518
rect -1042 1414 -1002 7360
rect -608 1414 -556 7360
rect -1042 1238 -556 1414
rect -2 1026 48 7522
rect 2028 7310 2132 7868
rect 2064 1040 2114 7310
rect 4112 1094 4162 7590
rect 4 510 60 924
rect 4120 510 4176 916
rect 2 412 4176 510
rect 4120 406 4176 412
<< viali >>
rect -962 1658 -650 7226
<< metal1 >>
rect -1042 7226 -556 7518
rect -1042 1658 -962 7226
rect -650 1658 -556 7226
rect -1042 1238 -556 1658
use sky130_fd_pr__nfet_g5v0d10v5_S5BDQR  sky130_fd_pr__nfet_g5v0d10v5_S5BDQR_0 ~/layout test
timestamp 1634046683
transform 1 0 2087 0 1 4167
box -2087 -4167 2087 4167
<< end >>
