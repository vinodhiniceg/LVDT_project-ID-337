magic
tech sky130A
magscale 1 2
timestamp 1634120139
<< nwell >>
rect -426 -360 5484 1588
<< mvnsubdiff >>
rect -326 1270 -56 1332
rect -326 204 -302 1270
rect -108 204 -56 1270
rect -326 96 -56 204
<< mvnsubdiffcont >>
rect -302 204 -108 1270
<< poly >>
rect 206 670 578 740
rect 888 668 1260 738
rect 1514 676 1886 746
rect 2212 674 2584 744
rect 2842 670 3214 740
rect 3506 672 3878 742
rect 4172 670 4544 740
rect 4784 670 5156 740
<< locali >>
rect -326 1270 -56 1332
rect 2678 1292 2748 1310
rect 36 1284 5364 1292
rect -326 204 -302 1270
rect -108 204 -56 1270
rect 28 1210 5364 1284
rect 28 1040 98 1210
rect 1360 1146 1430 1210
rect 2678 1158 2748 1210
rect 34 340 92 1040
rect 690 350 748 1146
rect 1354 1036 1430 1146
rect -326 96 -56 204
rect 680 152 776 350
rect 1354 344 1412 1036
rect 2006 370 2064 1154
rect 2674 1066 2748 1158
rect 1996 152 2092 370
rect 2674 356 2732 1066
rect 3324 362 3382 1142
rect 3982 1048 4052 1210
rect 3324 152 3420 362
rect 3994 340 4052 1048
rect 4644 366 4702 1126
rect 5288 1048 5358 1210
rect 4634 152 4730 366
rect 5300 324 5358 1048
rect 680 84 4730 152
rect 680 68 776 84
rect 3324 80 3420 84
<< viali >>
rect -256 266 -148 1224
<< metal1 >>
rect -326 1224 -56 1332
rect -326 266 -256 1224
rect -148 266 -56 1224
rect -326 96 -56 266
use sky130_fd_pr__pfet_g5v0d10v5_JRTA4Z  sky130_fd_pr__pfet_g5v0d10v5_JRTA4Z_0 ~/layout test
timestamp 1634119395
transform 1 0 2697 0 1 709
box -2727 -713 2727 713
<< end >>
